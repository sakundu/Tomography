VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram45_256x12
  FOREIGN fakeram45_256x12 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 57.570 BY 133.000 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.765 0.070 2.835 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.285 0.070 5.355 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.805 0.070 7.875 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.325 0.070 10.395 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.845 0.070 12.915 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.365 0.070 15.435 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.885 0.070 17.955 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.405 0.070 20.475 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.925 0.070 22.995 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.445 0.070 25.515 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.965 0.070 28.035 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.485 0.070 30.555 ;
    END
  END w_mask_in[11]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.725 0.070 32.795 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.245 0.070 35.315 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.765 0.070 37.835 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.285 0.070 40.355 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.805 0.070 42.875 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.325 0.070 45.395 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.845 0.070 47.915 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.365 0.070 50.435 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.885 0.070 52.955 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.405 0.070 55.475 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.925 0.070 57.995 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.445 0.070 60.515 ;
    END
  END rd_out[11]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 62.685 0.070 62.755 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 65.205 0.070 65.275 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 67.725 0.070 67.795 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.245 0.070 70.315 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.765 0.070 72.835 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.285 0.070 75.355 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.805 0.070 77.875 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.325 0.070 80.395 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.845 0.070 82.915 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.365 0.070 85.435 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 87.885 0.070 87.955 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 90.405 0.070 90.475 ;
    END
  END wd_in[11]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 92.645 0.070 92.715 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 95.165 0.070 95.235 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 97.685 0.070 97.755 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 100.205 0.070 100.275 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 102.725 0.070 102.795 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 105.245 0.070 105.315 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 107.765 0.070 107.835 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 110.285 0.070 110.355 ;
    END
  END addr_in[7]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 112.525 0.070 112.595 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 115.045 0.070 115.115 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 117.565 0.070 117.635 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 2.660 2.800 2.940 130.200 ;
      RECT 7.140 2.800 7.420 130.200 ;
      RECT 11.620 2.800 11.900 130.200 ;
      RECT 16.100 2.800 16.380 130.200 ;
      RECT 20.580 2.800 20.860 130.200 ;
      RECT 25.060 2.800 25.340 130.200 ;
      RECT 29.540 2.800 29.820 130.200 ;
      RECT 34.020 2.800 34.300 130.200 ;
      RECT 38.500 2.800 38.780 130.200 ;
      RECT 42.980 2.800 43.260 130.200 ;
      RECT 47.460 2.800 47.740 130.200 ;
      RECT 51.940 2.800 52.220 130.200 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 4.900 2.800 5.180 130.200 ;
      RECT 9.380 2.800 9.660 130.200 ;
      RECT 13.860 2.800 14.140 130.200 ;
      RECT 18.340 2.800 18.620 130.200 ;
      RECT 22.820 2.800 23.100 130.200 ;
      RECT 27.300 2.800 27.580 130.200 ;
      RECT 31.780 2.800 32.060 130.200 ;
      RECT 36.260 2.800 36.540 130.200 ;
      RECT 40.740 2.800 41.020 130.200 ;
      RECT 45.220 2.800 45.500 130.200 ;
      RECT 49.700 2.800 49.980 130.200 ;
      RECT 54.180 2.800 54.460 130.200 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 57.570 133.000 ;
    LAYER metal2 ;
    RECT 0 0 57.570 133.000 ;
    LAYER metal3 ;
    RECT 0.070 0 57.570 133.000 ;
    RECT 0 0.000 0.070 2.765 ;
    RECT 0 2.835 0.070 5.285 ;
    RECT 0 5.355 0.070 7.805 ;
    RECT 0 7.875 0.070 10.325 ;
    RECT 0 10.395 0.070 12.845 ;
    RECT 0 12.915 0.070 15.365 ;
    RECT 0 15.435 0.070 17.885 ;
    RECT 0 17.955 0.070 20.405 ;
    RECT 0 20.475 0.070 22.925 ;
    RECT 0 22.995 0.070 25.445 ;
    RECT 0 25.515 0.070 27.965 ;
    RECT 0 28.035 0.070 30.485 ;
    RECT 0 30.555 0.070 32.725 ;
    RECT 0 32.795 0.070 35.245 ;
    RECT 0 35.315 0.070 37.765 ;
    RECT 0 37.835 0.070 40.285 ;
    RECT 0 40.355 0.070 42.805 ;
    RECT 0 42.875 0.070 45.325 ;
    RECT 0 45.395 0.070 47.845 ;
    RECT 0 47.915 0.070 50.365 ;
    RECT 0 50.435 0.070 52.885 ;
    RECT 0 52.955 0.070 55.405 ;
    RECT 0 55.475 0.070 57.925 ;
    RECT 0 57.995 0.070 60.445 ;
    RECT 0 60.515 0.070 62.685 ;
    RECT 0 62.755 0.070 65.205 ;
    RECT 0 65.275 0.070 67.725 ;
    RECT 0 67.795 0.070 70.245 ;
    RECT 0 70.315 0.070 72.765 ;
    RECT 0 72.835 0.070 75.285 ;
    RECT 0 75.355 0.070 77.805 ;
    RECT 0 77.875 0.070 80.325 ;
    RECT 0 80.395 0.070 82.845 ;
    RECT 0 82.915 0.070 85.365 ;
    RECT 0 85.435 0.070 87.885 ;
    RECT 0 87.955 0.070 90.405 ;
    RECT 0 90.475 0.070 92.645 ;
    RECT 0 92.715 0.070 95.165 ;
    RECT 0 95.235 0.070 97.685 ;
    RECT 0 97.755 0.070 100.205 ;
    RECT 0 100.275 0.070 102.725 ;
    RECT 0 102.795 0.070 105.245 ;
    RECT 0 105.315 0.070 107.765 ;
    RECT 0 107.835 0.070 110.285 ;
    RECT 0 110.355 0.070 112.525 ;
    RECT 0 112.595 0.070 115.045 ;
    RECT 0 115.115 0.070 117.565 ;
    RECT 0 117.635 0.070 133.000 ;
    LAYER metal4 ;
    RECT 0 0 57.570 2.800 ;
    RECT 0 130.200 57.570 133.000 ;
    RECT 0.000 2.800 2.660 130.200 ;
    RECT 2.940 2.800 4.900 130.200 ;
    RECT 5.180 2.800 7.140 130.200 ;
    RECT 7.420 2.800 9.380 130.200 ;
    RECT 9.660 2.800 11.620 130.200 ;
    RECT 11.900 2.800 13.860 130.200 ;
    RECT 14.140 2.800 16.100 130.200 ;
    RECT 16.380 2.800 18.340 130.200 ;
    RECT 18.620 2.800 20.580 130.200 ;
    RECT 20.860 2.800 22.820 130.200 ;
    RECT 23.100 2.800 25.060 130.200 ;
    RECT 25.340 2.800 27.300 130.200 ;
    RECT 27.580 2.800 29.540 130.200 ;
    RECT 29.820 2.800 31.780 130.200 ;
    RECT 32.060 2.800 34.020 130.200 ;
    RECT 34.300 2.800 36.260 130.200 ;
    RECT 36.540 2.800 38.500 130.200 ;
    RECT 38.780 2.800 40.740 130.200 ;
    RECT 41.020 2.800 42.980 130.200 ;
    RECT 43.260 2.800 45.220 130.200 ;
    RECT 45.500 2.800 47.460 130.200 ;
    RECT 47.740 2.800 49.700 130.200 ;
    RECT 49.980 2.800 51.940 130.200 ;
    RECT 52.220 2.800 54.180 130.200 ;
    RECT 54.460 2.800 57.570 130.200 ;
    LAYER OVERLAP ;
    RECT 0 0 57.570 133.000 ;
  END
END fakeram45_256x12

END LIBRARY
