module mesh(clk, in, out);
input clk, in;
output out;
AOI211_X1 g_4_4 (.ZN (n_4_4) );
AOI211_X1 g_5_2 (.ZN (n_5_2) );
AOI211_X1 g_7_1 (.ZN (n_7_1), .A (n_4_4) );
AOI211_X1 g_9_2 (.ZN (n_9_2), .A (n_5_2) );
AOI211_X1 g_11_1 (.ZN (n_11_1), .A (n_7_1) );
AOI211_X1 g_13_2 (.ZN (n_13_2), .A (n_9_2), .B (n_4_4) );
AOI211_X1 g_15_1 (.ZN (n_15_1), .A (n_11_1), .B (n_5_2) );
AOI211_X1 g_17_2 (.ZN (n_17_2), .A (n_13_2), .B (n_7_1), .C1 (n_4_4) );
AOI211_X1 g_19_1 (.ZN (n_19_1), .A (n_15_1), .B (n_9_2), .C1 (n_5_2) );
AOI211_X1 g_21_2 (.ZN (n_21_2), .A (n_17_2), .B (n_11_1), .C1 (n_7_1) );
AOI211_X1 g_23_1 (.ZN (n_23_1), .A (n_19_1), .B (n_13_2), .C1 (n_9_2), .C2 (n_4_4) );
AOI211_X1 g_25_2 (.ZN (n_25_2), .A (n_21_2), .B (n_15_1), .C1 (n_11_1), .C2 (n_5_2) );
AOI211_X1 g_27_1 (.ZN (n_27_1), .A (n_23_1), .B (n_17_2), .C1 (n_13_2), .C2 (n_7_1) );
AOI211_X1 g_29_2 (.ZN (n_29_2), .A (n_25_2), .B (n_19_1), .C1 (n_15_1), .C2 (n_9_2) );
AOI211_X1 g_31_1 (.ZN (n_31_1), .A (n_27_1), .B (n_21_2), .C1 (n_17_2), .C2 (n_11_1) );
AOI211_X1 g_33_2 (.ZN (n_33_2), .A (n_29_2), .B (n_23_1), .C1 (n_19_1), .C2 (n_13_2) );
AOI211_X1 g_35_1 (.ZN (n_35_1), .A (n_31_1), .B (n_25_2), .C1 (n_21_2), .C2 (n_15_1) );
AOI211_X1 g_37_2 (.ZN (n_37_2), .A (n_33_2), .B (n_27_1), .C1 (n_23_1), .C2 (n_17_2) );
AOI211_X1 g_39_1 (.ZN (n_39_1), .A (n_35_1), .B (n_29_2), .C1 (n_25_2), .C2 (n_19_1) );
AOI211_X1 g_41_2 (.ZN (n_41_2), .A (n_37_2), .B (n_31_1), .C1 (n_27_1), .C2 (n_21_2) );
AOI211_X1 g_43_1 (.ZN (n_43_1), .A (n_39_1), .B (n_33_2), .C1 (n_29_2), .C2 (n_23_1) );
AOI211_X1 g_45_2 (.ZN (n_45_2), .A (n_41_2), .B (n_35_1), .C1 (n_31_1), .C2 (n_25_2) );
AOI211_X1 g_47_1 (.ZN (n_47_1), .A (n_43_1), .B (n_37_2), .C1 (n_33_2), .C2 (n_27_1) );
AOI211_X1 g_49_2 (.ZN (n_49_2), .A (n_45_2), .B (n_39_1), .C1 (n_35_1), .C2 (n_29_2) );
AOI211_X1 g_51_1 (.ZN (n_51_1), .A (n_47_1), .B (n_41_2), .C1 (n_37_2), .C2 (n_31_1) );
AOI211_X1 g_53_2 (.ZN (n_53_2), .A (n_49_2), .B (n_43_1), .C1 (n_39_1), .C2 (n_33_2) );
AOI211_X1 g_55_1 (.ZN (n_55_1), .A (n_51_1), .B (n_45_2), .C1 (n_41_2), .C2 (n_35_1) );
AOI211_X1 g_57_2 (.ZN (n_57_2), .A (n_53_2), .B (n_47_1), .C1 (n_43_1), .C2 (n_37_2) );
AOI211_X1 g_59_1 (.ZN (n_59_1), .A (n_55_1), .B (n_49_2), .C1 (n_45_2), .C2 (n_39_1) );
AOI211_X1 g_61_2 (.ZN (n_61_2), .A (n_57_2), .B (n_51_1), .C1 (n_47_1), .C2 (n_41_2) );
AOI211_X1 g_63_1 (.ZN (n_63_1), .A (n_59_1), .B (n_53_2), .C1 (n_49_2), .C2 (n_43_1) );
AOI211_X1 g_65_2 (.ZN (n_65_2), .A (n_61_2), .B (n_55_1), .C1 (n_51_1), .C2 (n_45_2) );
AOI211_X1 g_67_1 (.ZN (n_67_1), .A (n_63_1), .B (n_57_2), .C1 (n_53_2), .C2 (n_47_1) );
AOI211_X1 g_69_2 (.ZN (n_69_2), .A (n_65_2), .B (n_59_1), .C1 (n_55_1), .C2 (n_49_2) );
AOI211_X1 g_71_1 (.ZN (n_71_1), .A (n_67_1), .B (n_61_2), .C1 (n_57_2), .C2 (n_51_1) );
AOI211_X1 g_73_2 (.ZN (n_73_2), .A (n_69_2), .B (n_63_1), .C1 (n_59_1), .C2 (n_53_2) );
AOI211_X1 g_75_1 (.ZN (n_75_1), .A (n_71_1), .B (n_65_2), .C1 (n_61_2), .C2 (n_55_1) );
AOI211_X1 g_77_2 (.ZN (n_77_2), .A (n_73_2), .B (n_67_1), .C1 (n_63_1), .C2 (n_57_2) );
AOI211_X1 g_79_1 (.ZN (n_79_1), .A (n_75_1), .B (n_69_2), .C1 (n_65_2), .C2 (n_59_1) );
AOI211_X1 g_81_2 (.ZN (n_81_2), .A (n_77_2), .B (n_71_1), .C1 (n_67_1), .C2 (n_61_2) );
AOI211_X1 g_83_1 (.ZN (n_83_1), .A (n_79_1), .B (n_73_2), .C1 (n_69_2), .C2 (n_63_1) );
AOI211_X1 g_85_2 (.ZN (n_85_2), .A (n_81_2), .B (n_75_1), .C1 (n_71_1), .C2 (n_65_2) );
AOI211_X1 g_87_1 (.ZN (n_87_1), .A (n_83_1), .B (n_77_2), .C1 (n_73_2), .C2 (n_67_1) );
AOI211_X1 g_89_2 (.ZN (n_89_2), .A (n_85_2), .B (n_79_1), .C1 (n_75_1), .C2 (n_69_2) );
AOI211_X1 g_91_1 (.ZN (n_91_1), .A (n_87_1), .B (n_81_2), .C1 (n_77_2), .C2 (n_71_1) );
AOI211_X1 g_93_2 (.ZN (n_93_2), .A (n_89_2), .B (n_83_1), .C1 (n_79_1), .C2 (n_73_2) );
AOI211_X1 g_95_1 (.ZN (n_95_1), .A (n_91_1), .B (n_85_2), .C1 (n_81_2), .C2 (n_75_1) );
AOI211_X1 g_97_2 (.ZN (n_97_2), .A (n_93_2), .B (n_87_1), .C1 (n_83_1), .C2 (n_77_2) );
AOI211_X1 g_99_1 (.ZN (n_99_1), .A (n_95_1), .B (n_89_2), .C1 (n_85_2), .C2 (n_79_1) );
AOI211_X1 g_101_2 (.ZN (n_101_2), .A (n_97_2), .B (n_91_1), .C1 (n_87_1), .C2 (n_81_2) );
AOI211_X1 g_103_1 (.ZN (n_103_1), .A (n_99_1), .B (n_93_2), .C1 (n_89_2), .C2 (n_83_1) );
AOI211_X1 g_105_2 (.ZN (n_105_2), .A (n_101_2), .B (n_95_1), .C1 (n_91_1), .C2 (n_85_2) );
AOI211_X1 g_107_1 (.ZN (n_107_1), .A (n_103_1), .B (n_97_2), .C1 (n_93_2), .C2 (n_87_1) );
AOI211_X1 g_109_2 (.ZN (n_109_2), .A (n_105_2), .B (n_99_1), .C1 (n_95_1), .C2 (n_89_2) );
AOI211_X1 g_111_1 (.ZN (n_111_1), .A (n_107_1), .B (n_101_2), .C1 (n_97_2), .C2 (n_91_1) );
AOI211_X1 g_113_2 (.ZN (n_113_2), .A (n_109_2), .B (n_103_1), .C1 (n_99_1), .C2 (n_93_2) );
AOI211_X1 g_115_1 (.ZN (n_115_1), .A (n_111_1), .B (n_105_2), .C1 (n_101_2), .C2 (n_95_1) );
AOI211_X1 g_117_2 (.ZN (n_117_2), .A (n_113_2), .B (n_107_1), .C1 (n_103_1), .C2 (n_97_2) );
AOI211_X1 g_119_1 (.ZN (n_119_1), .A (n_115_1), .B (n_109_2), .C1 (n_105_2), .C2 (n_99_1) );
AOI211_X1 g_121_2 (.ZN (n_121_2), .A (n_117_2), .B (n_111_1), .C1 (n_107_1), .C2 (n_101_2) );
AOI211_X1 g_123_1 (.ZN (n_123_1), .A (n_119_1), .B (n_113_2), .C1 (n_109_2), .C2 (n_103_1) );
AOI211_X1 g_125_2 (.ZN (n_125_2), .A (n_121_2), .B (n_115_1), .C1 (n_111_1), .C2 (n_105_2) );
AOI211_X1 g_127_1 (.ZN (n_127_1), .A (n_123_1), .B (n_117_2), .C1 (n_113_2), .C2 (n_107_1) );
AOI211_X1 g_129_2 (.ZN (n_129_2), .A (n_125_2), .B (n_119_1), .C1 (n_115_1), .C2 (n_109_2) );
AOI211_X1 g_131_1 (.ZN (n_131_1), .A (n_127_1), .B (n_121_2), .C1 (n_117_2), .C2 (n_111_1) );
AOI211_X1 g_133_2 (.ZN (n_133_2), .A (n_129_2), .B (n_123_1), .C1 (n_119_1), .C2 (n_113_2) );
AOI211_X1 g_135_1 (.ZN (n_135_1), .A (n_131_1), .B (n_125_2), .C1 (n_121_2), .C2 (n_115_1) );
AOI211_X1 g_137_2 (.ZN (n_137_2), .A (n_133_2), .B (n_127_1), .C1 (n_123_1), .C2 (n_117_2) );
AOI211_X1 g_139_1 (.ZN (n_139_1), .A (n_135_1), .B (n_129_2), .C1 (n_125_2), .C2 (n_119_1) );
AOI211_X1 g_141_2 (.ZN (n_141_2), .A (n_137_2), .B (n_131_1), .C1 (n_127_1), .C2 (n_121_2) );
AOI211_X1 g_143_1 (.ZN (n_143_1), .A (n_139_1), .B (n_133_2), .C1 (n_129_2), .C2 (n_123_1) );
AOI211_X1 g_145_2 (.ZN (n_145_2), .A (n_141_2), .B (n_135_1), .C1 (n_131_1), .C2 (n_125_2) );
AOI211_X1 g_147_1 (.ZN (n_147_1), .A (n_143_1), .B (n_137_2), .C1 (n_133_2), .C2 (n_127_1) );
AOI211_X1 g_149_2 (.ZN (n_149_2), .A (n_145_2), .B (n_139_1), .C1 (n_135_1), .C2 (n_129_2) );
AOI211_X1 g_150_4 (.ZN (n_150_4), .A (n_147_1), .B (n_141_2), .C1 (n_137_2), .C2 (n_131_1) );
AOI211_X1 g_149_6 (.ZN (n_149_6), .A (n_149_2), .B (n_143_1), .C1 (n_139_1), .C2 (n_133_2) );
AOI211_X1 g_150_8 (.ZN (n_150_8), .A (n_150_4), .B (n_145_2), .C1 (n_141_2), .C2 (n_135_1) );
AOI211_X1 g_149_10 (.ZN (n_149_10), .A (n_149_6), .B (n_147_1), .C1 (n_143_1), .C2 (n_137_2) );
AOI211_X1 g_150_12 (.ZN (n_150_12), .A (n_150_8), .B (n_149_2), .C1 (n_145_2), .C2 (n_139_1) );
AOI211_X1 g_149_14 (.ZN (n_149_14), .A (n_149_10), .B (n_150_4), .C1 (n_147_1), .C2 (n_141_2) );
AOI211_X1 g_150_16 (.ZN (n_150_16), .A (n_150_12), .B (n_149_6), .C1 (n_149_2), .C2 (n_143_1) );
AOI211_X1 g_149_18 (.ZN (n_149_18), .A (n_149_14), .B (n_150_8), .C1 (n_150_4), .C2 (n_145_2) );
AOI211_X1 g_150_20 (.ZN (n_150_20), .A (n_150_16), .B (n_149_10), .C1 (n_149_6), .C2 (n_147_1) );
AOI211_X1 g_149_22 (.ZN (n_149_22), .A (n_149_18), .B (n_150_12), .C1 (n_150_8), .C2 (n_149_2) );
AOI211_X1 g_150_24 (.ZN (n_150_24), .A (n_150_20), .B (n_149_14), .C1 (n_149_10), .C2 (n_150_4) );
AOI211_X1 g_149_26 (.ZN (n_149_26), .A (n_149_22), .B (n_150_16), .C1 (n_150_12), .C2 (n_149_6) );
AOI211_X1 g_150_28 (.ZN (n_150_28), .A (n_150_24), .B (n_149_18), .C1 (n_149_14), .C2 (n_150_8) );
AOI211_X1 g_149_30 (.ZN (n_149_30), .A (n_149_26), .B (n_150_20), .C1 (n_150_16), .C2 (n_149_10) );
AOI211_X1 g_150_32 (.ZN (n_150_32), .A (n_150_28), .B (n_149_22), .C1 (n_149_18), .C2 (n_150_12) );
AOI211_X1 g_149_34 (.ZN (n_149_34), .A (n_149_30), .B (n_150_24), .C1 (n_150_20), .C2 (n_149_14) );
AOI211_X1 g_150_36 (.ZN (n_150_36), .A (n_150_32), .B (n_149_26), .C1 (n_149_22), .C2 (n_150_16) );
AOI211_X1 g_149_38 (.ZN (n_149_38), .A (n_149_34), .B (n_150_28), .C1 (n_150_24), .C2 (n_149_18) );
AOI211_X1 g_150_40 (.ZN (n_150_40), .A (n_150_36), .B (n_149_30), .C1 (n_149_26), .C2 (n_150_20) );
AOI211_X1 g_149_42 (.ZN (n_149_42), .A (n_149_38), .B (n_150_32), .C1 (n_150_28), .C2 (n_149_22) );
AOI211_X1 g_150_44 (.ZN (n_150_44), .A (n_150_40), .B (n_149_34), .C1 (n_149_30), .C2 (n_150_24) );
AOI211_X1 g_149_46 (.ZN (n_149_46), .A (n_149_42), .B (n_150_36), .C1 (n_150_32), .C2 (n_149_26) );
AOI211_X1 g_150_48 (.ZN (n_150_48), .A (n_150_44), .B (n_149_38), .C1 (n_149_34), .C2 (n_150_28) );
AOI211_X1 g_149_50 (.ZN (n_149_50), .A (n_149_46), .B (n_150_40), .C1 (n_150_36), .C2 (n_149_30) );
AOI211_X1 g_150_52 (.ZN (n_150_52), .A (n_150_48), .B (n_149_42), .C1 (n_149_38), .C2 (n_150_32) );
AOI211_X1 g_149_54 (.ZN (n_149_54), .A (n_149_50), .B (n_150_44), .C1 (n_150_40), .C2 (n_149_34) );
AOI211_X1 g_150_56 (.ZN (n_150_56), .A (n_150_52), .B (n_149_46), .C1 (n_149_42), .C2 (n_150_36) );
AOI211_X1 g_149_58 (.ZN (n_149_58), .A (n_149_54), .B (n_150_48), .C1 (n_150_44), .C2 (n_149_38) );
AOI211_X1 g_150_60 (.ZN (n_150_60), .A (n_150_56), .B (n_149_50), .C1 (n_149_46), .C2 (n_150_40) );
AOI211_X1 g_149_62 (.ZN (n_149_62), .A (n_149_58), .B (n_150_52), .C1 (n_150_48), .C2 (n_149_42) );
AOI211_X1 g_150_64 (.ZN (n_150_64), .A (n_150_60), .B (n_149_54), .C1 (n_149_50), .C2 (n_150_44) );
AOI211_X1 g_149_66 (.ZN (n_149_66), .A (n_149_62), .B (n_150_56), .C1 (n_150_52), .C2 (n_149_46) );
AOI211_X1 g_150_68 (.ZN (n_150_68), .A (n_150_64), .B (n_149_58), .C1 (n_149_54), .C2 (n_150_48) );
AOI211_X1 g_149_70 (.ZN (n_149_70), .A (n_149_66), .B (n_150_60), .C1 (n_150_56), .C2 (n_149_50) );
AOI211_X1 g_150_72 (.ZN (n_150_72), .A (n_150_68), .B (n_149_62), .C1 (n_149_58), .C2 (n_150_52) );
AOI211_X1 g_149_74 (.ZN (n_149_74), .A (n_149_70), .B (n_150_64), .C1 (n_150_60), .C2 (n_149_54) );
AOI211_X1 g_150_76 (.ZN (n_150_76), .A (n_150_72), .B (n_149_66), .C1 (n_149_62), .C2 (n_150_56) );
AOI211_X1 g_149_78 (.ZN (n_149_78), .A (n_149_74), .B (n_150_68), .C1 (n_150_64), .C2 (n_149_58) );
AOI211_X1 g_150_80 (.ZN (n_150_80), .A (n_150_76), .B (n_149_70), .C1 (n_149_66), .C2 (n_150_60) );
AOI211_X1 g_149_82 (.ZN (n_149_82), .A (n_149_78), .B (n_150_72), .C1 (n_150_68), .C2 (n_149_62) );
AOI211_X1 g_150_84 (.ZN (n_150_84), .A (n_150_80), .B (n_149_74), .C1 (n_149_70), .C2 (n_150_64) );
AOI211_X1 g_149_86 (.ZN (n_149_86), .A (n_149_82), .B (n_150_76), .C1 (n_150_72), .C2 (n_149_66) );
AOI211_X1 g_150_88 (.ZN (n_150_88), .A (n_150_84), .B (n_149_78), .C1 (n_149_74), .C2 (n_150_68) );
AOI211_X1 g_149_90 (.ZN (n_149_90), .A (n_149_86), .B (n_150_80), .C1 (n_150_76), .C2 (n_149_70) );
AOI211_X1 g_150_92 (.ZN (n_150_92), .A (n_150_88), .B (n_149_82), .C1 (n_149_78), .C2 (n_150_72) );
AOI211_X1 g_149_94 (.ZN (n_149_94), .A (n_149_90), .B (n_150_84), .C1 (n_150_80), .C2 (n_149_74) );
AOI211_X1 g_150_96 (.ZN (n_150_96), .A (n_150_92), .B (n_149_86), .C1 (n_149_82), .C2 (n_150_76) );
AOI211_X1 g_149_98 (.ZN (n_149_98), .A (n_149_94), .B (n_150_88), .C1 (n_150_84), .C2 (n_149_78) );
AOI211_X1 g_150_100 (.ZN (n_150_100), .A (n_150_96), .B (n_149_90), .C1 (n_149_86), .C2 (n_150_80) );
AOI211_X1 g_149_102 (.ZN (n_149_102), .A (n_149_98), .B (n_150_92), .C1 (n_150_88), .C2 (n_149_82) );
AOI211_X1 g_150_104 (.ZN (n_150_104), .A (n_150_100), .B (n_149_94), .C1 (n_149_90), .C2 (n_150_84) );
AOI211_X1 g_149_106 (.ZN (n_149_106), .A (n_149_102), .B (n_150_96), .C1 (n_150_92), .C2 (n_149_86) );
AOI211_X1 g_150_108 (.ZN (n_150_108), .A (n_150_104), .B (n_149_98), .C1 (n_149_94), .C2 (n_150_88) );
AOI211_X1 g_149_110 (.ZN (n_149_110), .A (n_149_106), .B (n_150_100), .C1 (n_150_96), .C2 (n_149_90) );
AOI211_X1 g_150_112 (.ZN (n_150_112), .A (n_150_108), .B (n_149_102), .C1 (n_149_98), .C2 (n_150_92) );
AOI211_X1 g_149_114 (.ZN (n_149_114), .A (n_149_110), .B (n_150_104), .C1 (n_150_100), .C2 (n_149_94) );
AOI211_X1 g_150_116 (.ZN (n_150_116), .A (n_150_112), .B (n_149_106), .C1 (n_149_102), .C2 (n_150_96) );
AOI211_X1 g_149_118 (.ZN (n_149_118), .A (n_149_114), .B (n_150_108), .C1 (n_150_104), .C2 (n_149_98) );
AOI211_X1 g_150_120 (.ZN (n_150_120), .A (n_150_116), .B (n_149_110), .C1 (n_149_106), .C2 (n_150_100) );
AOI211_X1 g_149_122 (.ZN (n_149_122), .A (n_149_118), .B (n_150_112), .C1 (n_150_108), .C2 (n_149_102) );
AOI211_X1 g_150_124 (.ZN (n_150_124), .A (n_150_120), .B (n_149_114), .C1 (n_149_110), .C2 (n_150_104) );
AOI211_X1 g_149_126 (.ZN (n_149_126), .A (n_149_122), .B (n_150_116), .C1 (n_150_112), .C2 (n_149_106) );
AOI211_X1 g_150_128 (.ZN (n_150_128), .A (n_150_124), .B (n_149_118), .C1 (n_149_114), .C2 (n_150_108) );
AOI211_X1 g_149_130 (.ZN (n_149_130), .A (n_149_126), .B (n_150_120), .C1 (n_150_116), .C2 (n_149_110) );
AOI211_X1 g_150_132 (.ZN (n_150_132), .A (n_150_128), .B (n_149_122), .C1 (n_149_118), .C2 (n_150_112) );
AOI211_X1 g_149_134 (.ZN (n_149_134), .A (n_149_130), .B (n_150_124), .C1 (n_150_120), .C2 (n_149_114) );
AOI211_X1 g_150_136 (.ZN (n_150_136), .A (n_150_132), .B (n_149_126), .C1 (n_149_122), .C2 (n_150_116) );
AOI211_X1 g_149_138 (.ZN (n_149_138), .A (n_149_134), .B (n_150_128), .C1 (n_150_124), .C2 (n_149_118) );
AOI211_X1 g_150_140 (.ZN (n_150_140), .A (n_150_136), .B (n_149_130), .C1 (n_149_126), .C2 (n_150_120) );
AOI211_X1 g_149_142 (.ZN (n_149_142), .A (n_149_138), .B (n_150_132), .C1 (n_150_128), .C2 (n_149_122) );
AOI211_X1 g_150_144 (.ZN (n_150_144), .A (n_150_140), .B (n_149_134), .C1 (n_149_130), .C2 (n_150_124) );
AOI211_X1 g_149_146 (.ZN (n_149_146), .A (n_149_142), .B (n_150_136), .C1 (n_150_132), .C2 (n_149_126) );
AOI211_X1 g_150_148 (.ZN (n_150_148), .A (n_150_144), .B (n_149_138), .C1 (n_149_134), .C2 (n_150_128) );
AOI211_X1 g_149_150 (.ZN (n_149_150), .A (n_149_146), .B (n_150_140), .C1 (n_150_136), .C2 (n_149_130) );
AOI211_X1 g_147_149 (.ZN (n_147_149), .A (n_150_148), .B (n_149_142), .C1 (n_149_138), .C2 (n_150_132) );
AOI211_X1 g_145_150 (.ZN (n_145_150), .A (n_149_150), .B (n_150_144), .C1 (n_150_140), .C2 (n_149_134) );
AOI211_X1 g_143_149 (.ZN (n_143_149), .A (n_147_149), .B (n_149_146), .C1 (n_149_142), .C2 (n_150_136) );
AOI211_X1 g_141_150 (.ZN (n_141_150), .A (n_145_150), .B (n_150_148), .C1 (n_150_144), .C2 (n_149_138) );
AOI211_X1 g_139_149 (.ZN (n_139_149), .A (n_143_149), .B (n_149_150), .C1 (n_149_146), .C2 (n_150_140) );
AOI211_X1 g_137_150 (.ZN (n_137_150), .A (n_141_150), .B (n_147_149), .C1 (n_150_148), .C2 (n_149_142) );
AOI211_X1 g_135_149 (.ZN (n_135_149), .A (n_139_149), .B (n_145_150), .C1 (n_149_150), .C2 (n_150_144) );
AOI211_X1 g_133_150 (.ZN (n_133_150), .A (n_137_150), .B (n_143_149), .C1 (n_147_149), .C2 (n_149_146) );
AOI211_X1 g_131_149 (.ZN (n_131_149), .A (n_135_149), .B (n_141_150), .C1 (n_145_150), .C2 (n_150_148) );
AOI211_X1 g_129_150 (.ZN (n_129_150), .A (n_133_150), .B (n_139_149), .C1 (n_143_149), .C2 (n_149_150) );
AOI211_X1 g_127_149 (.ZN (n_127_149), .A (n_131_149), .B (n_137_150), .C1 (n_141_150), .C2 (n_147_149) );
AOI211_X1 g_125_150 (.ZN (n_125_150), .A (n_129_150), .B (n_135_149), .C1 (n_139_149), .C2 (n_145_150) );
AOI211_X1 g_123_149 (.ZN (n_123_149), .A (n_127_149), .B (n_133_150), .C1 (n_137_150), .C2 (n_143_149) );
AOI211_X1 g_121_150 (.ZN (n_121_150), .A (n_125_150), .B (n_131_149), .C1 (n_135_149), .C2 (n_141_150) );
AOI211_X1 g_119_149 (.ZN (n_119_149), .A (n_123_149), .B (n_129_150), .C1 (n_133_150), .C2 (n_139_149) );
AOI211_X1 g_117_150 (.ZN (n_117_150), .A (n_121_150), .B (n_127_149), .C1 (n_131_149), .C2 (n_137_150) );
AOI211_X1 g_115_149 (.ZN (n_115_149), .A (n_119_149), .B (n_125_150), .C1 (n_129_150), .C2 (n_135_149) );
AOI211_X1 g_113_150 (.ZN (n_113_150), .A (n_117_150), .B (n_123_149), .C1 (n_127_149), .C2 (n_133_150) );
AOI211_X1 g_111_149 (.ZN (n_111_149), .A (n_115_149), .B (n_121_150), .C1 (n_125_150), .C2 (n_131_149) );
AOI211_X1 g_109_150 (.ZN (n_109_150), .A (n_113_150), .B (n_119_149), .C1 (n_123_149), .C2 (n_129_150) );
AOI211_X1 g_107_149 (.ZN (n_107_149), .A (n_111_149), .B (n_117_150), .C1 (n_121_150), .C2 (n_127_149) );
AOI211_X1 g_105_150 (.ZN (n_105_150), .A (n_109_150), .B (n_115_149), .C1 (n_119_149), .C2 (n_125_150) );
AOI211_X1 g_103_149 (.ZN (n_103_149), .A (n_107_149), .B (n_113_150), .C1 (n_117_150), .C2 (n_123_149) );
AOI211_X1 g_101_150 (.ZN (n_101_150), .A (n_105_150), .B (n_111_149), .C1 (n_115_149), .C2 (n_121_150) );
AOI211_X1 g_99_149 (.ZN (n_99_149), .A (n_103_149), .B (n_109_150), .C1 (n_113_150), .C2 (n_119_149) );
AOI211_X1 g_97_150 (.ZN (n_97_150), .A (n_101_150), .B (n_107_149), .C1 (n_111_149), .C2 (n_117_150) );
AOI211_X1 g_95_149 (.ZN (n_95_149), .A (n_99_149), .B (n_105_150), .C1 (n_109_150), .C2 (n_115_149) );
AOI211_X1 g_93_150 (.ZN (n_93_150), .A (n_97_150), .B (n_103_149), .C1 (n_107_149), .C2 (n_113_150) );
AOI211_X1 g_91_149 (.ZN (n_91_149), .A (n_95_149), .B (n_101_150), .C1 (n_105_150), .C2 (n_111_149) );
AOI211_X1 g_89_150 (.ZN (n_89_150), .A (n_93_150), .B (n_99_149), .C1 (n_103_149), .C2 (n_109_150) );
AOI211_X1 g_87_149 (.ZN (n_87_149), .A (n_91_149), .B (n_97_150), .C1 (n_101_150), .C2 (n_107_149) );
AOI211_X1 g_85_150 (.ZN (n_85_150), .A (n_89_150), .B (n_95_149), .C1 (n_99_149), .C2 (n_105_150) );
AOI211_X1 g_83_149 (.ZN (n_83_149), .A (n_87_149), .B (n_93_150), .C1 (n_97_150), .C2 (n_103_149) );
AOI211_X1 g_81_150 (.ZN (n_81_150), .A (n_85_150), .B (n_91_149), .C1 (n_95_149), .C2 (n_101_150) );
AOI211_X1 g_79_149 (.ZN (n_79_149), .A (n_83_149), .B (n_89_150), .C1 (n_93_150), .C2 (n_99_149) );
AOI211_X1 g_77_150 (.ZN (n_77_150), .A (n_81_150), .B (n_87_149), .C1 (n_91_149), .C2 (n_97_150) );
AOI211_X1 g_75_149 (.ZN (n_75_149), .A (n_79_149), .B (n_85_150), .C1 (n_89_150), .C2 (n_95_149) );
AOI211_X1 g_73_150 (.ZN (n_73_150), .A (n_77_150), .B (n_83_149), .C1 (n_87_149), .C2 (n_93_150) );
AOI211_X1 g_71_149 (.ZN (n_71_149), .A (n_75_149), .B (n_81_150), .C1 (n_85_150), .C2 (n_91_149) );
AOI211_X1 g_69_150 (.ZN (n_69_150), .A (n_73_150), .B (n_79_149), .C1 (n_83_149), .C2 (n_89_150) );
AOI211_X1 g_67_149 (.ZN (n_67_149), .A (n_71_149), .B (n_77_150), .C1 (n_81_150), .C2 (n_87_149) );
AOI211_X1 g_65_150 (.ZN (n_65_150), .A (n_69_150), .B (n_75_149), .C1 (n_79_149), .C2 (n_85_150) );
AOI211_X1 g_63_149 (.ZN (n_63_149), .A (n_67_149), .B (n_73_150), .C1 (n_77_150), .C2 (n_83_149) );
AOI211_X1 g_61_150 (.ZN (n_61_150), .A (n_65_150), .B (n_71_149), .C1 (n_75_149), .C2 (n_81_150) );
AOI211_X1 g_59_149 (.ZN (n_59_149), .A (n_63_149), .B (n_69_150), .C1 (n_73_150), .C2 (n_79_149) );
AOI211_X1 g_57_150 (.ZN (n_57_150), .A (n_61_150), .B (n_67_149), .C1 (n_71_149), .C2 (n_77_150) );
AOI211_X1 g_55_149 (.ZN (n_55_149), .A (n_59_149), .B (n_65_150), .C1 (n_69_150), .C2 (n_75_149) );
AOI211_X1 g_53_150 (.ZN (n_53_150), .A (n_57_150), .B (n_63_149), .C1 (n_67_149), .C2 (n_73_150) );
AOI211_X1 g_51_149 (.ZN (n_51_149), .A (n_55_149), .B (n_61_150), .C1 (n_65_150), .C2 (n_71_149) );
AOI211_X1 g_49_150 (.ZN (n_49_150), .A (n_53_150), .B (n_59_149), .C1 (n_63_149), .C2 (n_69_150) );
AOI211_X1 g_47_149 (.ZN (n_47_149), .A (n_51_149), .B (n_57_150), .C1 (n_61_150), .C2 (n_67_149) );
AOI211_X1 g_45_150 (.ZN (n_45_150), .A (n_49_150), .B (n_55_149), .C1 (n_59_149), .C2 (n_65_150) );
AOI211_X1 g_43_149 (.ZN (n_43_149), .A (n_47_149), .B (n_53_150), .C1 (n_57_150), .C2 (n_63_149) );
AOI211_X1 g_41_150 (.ZN (n_41_150), .A (n_45_150), .B (n_51_149), .C1 (n_55_149), .C2 (n_61_150) );
AOI211_X1 g_39_149 (.ZN (n_39_149), .A (n_43_149), .B (n_49_150), .C1 (n_53_150), .C2 (n_59_149) );
AOI211_X1 g_37_150 (.ZN (n_37_150), .A (n_41_150), .B (n_47_149), .C1 (n_51_149), .C2 (n_57_150) );
AOI211_X1 g_35_149 (.ZN (n_35_149), .A (n_39_149), .B (n_45_150), .C1 (n_49_150), .C2 (n_55_149) );
AOI211_X1 g_33_150 (.ZN (n_33_150), .A (n_37_150), .B (n_43_149), .C1 (n_47_149), .C2 (n_53_150) );
AOI211_X1 g_31_149 (.ZN (n_31_149), .A (n_35_149), .B (n_41_150), .C1 (n_45_150), .C2 (n_51_149) );
AOI211_X1 g_29_150 (.ZN (n_29_150), .A (n_33_150), .B (n_39_149), .C1 (n_43_149), .C2 (n_49_150) );
AOI211_X1 g_27_149 (.ZN (n_27_149), .A (n_31_149), .B (n_37_150), .C1 (n_41_150), .C2 (n_47_149) );
AOI211_X1 g_25_150 (.ZN (n_25_150), .A (n_29_150), .B (n_35_149), .C1 (n_39_149), .C2 (n_45_150) );
AOI211_X1 g_23_149 (.ZN (n_23_149), .A (n_27_149), .B (n_33_150), .C1 (n_37_150), .C2 (n_43_149) );
AOI211_X1 g_21_150 (.ZN (n_21_150), .A (n_25_150), .B (n_31_149), .C1 (n_35_149), .C2 (n_41_150) );
AOI211_X1 g_19_149 (.ZN (n_19_149), .A (n_23_149), .B (n_29_150), .C1 (n_33_150), .C2 (n_39_149) );
AOI211_X1 g_17_150 (.ZN (n_17_150), .A (n_21_150), .B (n_27_149), .C1 (n_31_149), .C2 (n_37_150) );
AOI211_X1 g_15_149 (.ZN (n_15_149), .A (n_19_149), .B (n_25_150), .C1 (n_29_150), .C2 (n_35_149) );
AOI211_X1 g_13_150 (.ZN (n_13_150), .A (n_17_150), .B (n_23_149), .C1 (n_27_149), .C2 (n_33_150) );
AOI211_X1 g_11_149 (.ZN (n_11_149), .A (n_15_149), .B (n_21_150), .C1 (n_25_150), .C2 (n_31_149) );
AOI211_X1 g_9_150 (.ZN (n_9_150), .A (n_13_150), .B (n_19_149), .C1 (n_23_149), .C2 (n_29_150) );
AOI211_X1 g_7_149 (.ZN (n_7_149), .A (n_11_149), .B (n_17_150), .C1 (n_21_150), .C2 (n_27_149) );
AOI211_X1 g_5_150 (.ZN (n_5_150), .A (n_9_150), .B (n_15_149), .C1 (n_19_149), .C2 (n_25_150) );
AOI211_X1 g_3_149 (.ZN (n_3_149), .A (n_7_149), .B (n_13_150), .C1 (n_17_150), .C2 (n_23_149) );
AOI211_X1 g_1_150 (.ZN (n_1_150), .A (n_5_150), .B (n_11_149), .C1 (n_15_149), .C2 (n_21_150) );
AOI211_X1 g_2_148 (.ZN (n_2_148), .A (n_3_149), .B (n_9_150), .C1 (n_13_150), .C2 (n_19_149) );
AOI211_X1 g_1_146 (.ZN (n_1_146), .A (n_1_150), .B (n_7_149), .C1 (n_11_149), .C2 (n_17_150) );
AOI211_X1 g_2_144 (.ZN (n_2_144), .A (n_2_148), .B (n_5_150), .C1 (n_9_150), .C2 (n_15_149) );
AOI211_X1 g_1_142 (.ZN (n_1_142), .A (n_1_146), .B (n_3_149), .C1 (n_7_149), .C2 (n_13_150) );
AOI211_X1 g_2_140 (.ZN (n_2_140), .A (n_2_144), .B (n_1_150), .C1 (n_5_150), .C2 (n_11_149) );
AOI211_X1 g_1_138 (.ZN (n_1_138), .A (n_1_142), .B (n_2_148), .C1 (n_3_149), .C2 (n_9_150) );
AOI211_X1 g_2_136 (.ZN (n_2_136), .A (n_2_140), .B (n_1_146), .C1 (n_1_150), .C2 (n_7_149) );
AOI211_X1 g_1_134 (.ZN (n_1_134), .A (n_1_138), .B (n_2_144), .C1 (n_2_148), .C2 (n_5_150) );
AOI211_X1 g_2_132 (.ZN (n_2_132), .A (n_2_136), .B (n_1_142), .C1 (n_1_146), .C2 (n_3_149) );
AOI211_X1 g_1_130 (.ZN (n_1_130), .A (n_1_134), .B (n_2_140), .C1 (n_2_144), .C2 (n_1_150) );
AOI211_X1 g_2_128 (.ZN (n_2_128), .A (n_2_132), .B (n_1_138), .C1 (n_1_142), .C2 (n_2_148) );
AOI211_X1 g_1_126 (.ZN (n_1_126), .A (n_1_130), .B (n_2_136), .C1 (n_2_140), .C2 (n_1_146) );
AOI211_X1 g_2_124 (.ZN (n_2_124), .A (n_2_128), .B (n_1_134), .C1 (n_1_138), .C2 (n_2_144) );
AOI211_X1 g_1_122 (.ZN (n_1_122), .A (n_1_126), .B (n_2_132), .C1 (n_2_136), .C2 (n_1_142) );
AOI211_X1 g_2_120 (.ZN (n_2_120), .A (n_2_124), .B (n_1_130), .C1 (n_1_134), .C2 (n_2_140) );
AOI211_X1 g_1_118 (.ZN (n_1_118), .A (n_1_122), .B (n_2_128), .C1 (n_2_132), .C2 (n_1_138) );
AOI211_X1 g_2_116 (.ZN (n_2_116), .A (n_2_120), .B (n_1_126), .C1 (n_1_130), .C2 (n_2_136) );
AOI211_X1 g_1_114 (.ZN (n_1_114), .A (n_1_118), .B (n_2_124), .C1 (n_2_128), .C2 (n_1_134) );
AOI211_X1 g_2_112 (.ZN (n_2_112), .A (n_2_116), .B (n_1_122), .C1 (n_1_126), .C2 (n_2_132) );
AOI211_X1 g_1_110 (.ZN (n_1_110), .A (n_1_114), .B (n_2_120), .C1 (n_2_124), .C2 (n_1_130) );
AOI211_X1 g_2_108 (.ZN (n_2_108), .A (n_2_112), .B (n_1_118), .C1 (n_1_122), .C2 (n_2_128) );
AOI211_X1 g_1_106 (.ZN (n_1_106), .A (n_1_110), .B (n_2_116), .C1 (n_2_120), .C2 (n_1_126) );
AOI211_X1 g_2_104 (.ZN (n_2_104), .A (n_2_108), .B (n_1_114), .C1 (n_1_118), .C2 (n_2_124) );
AOI211_X1 g_1_102 (.ZN (n_1_102), .A (n_1_106), .B (n_2_112), .C1 (n_2_116), .C2 (n_1_122) );
AOI211_X1 g_2_100 (.ZN (n_2_100), .A (n_2_104), .B (n_1_110), .C1 (n_1_114), .C2 (n_2_120) );
AOI211_X1 g_1_98 (.ZN (n_1_98), .A (n_1_102), .B (n_2_108), .C1 (n_2_112), .C2 (n_1_118) );
AOI211_X1 g_2_96 (.ZN (n_2_96), .A (n_2_100), .B (n_1_106), .C1 (n_1_110), .C2 (n_2_116) );
AOI211_X1 g_1_94 (.ZN (n_1_94), .A (n_1_98), .B (n_2_104), .C1 (n_2_108), .C2 (n_1_114) );
AOI211_X1 g_2_92 (.ZN (n_2_92), .A (n_2_96), .B (n_1_102), .C1 (n_1_106), .C2 (n_2_112) );
AOI211_X1 g_1_90 (.ZN (n_1_90), .A (n_1_94), .B (n_2_100), .C1 (n_2_104), .C2 (n_1_110) );
AOI211_X1 g_2_88 (.ZN (n_2_88), .A (n_2_92), .B (n_1_98), .C1 (n_1_102), .C2 (n_2_108) );
AOI211_X1 g_1_86 (.ZN (n_1_86), .A (n_1_90), .B (n_2_96), .C1 (n_2_100), .C2 (n_1_106) );
AOI211_X1 g_2_84 (.ZN (n_2_84), .A (n_2_88), .B (n_1_94), .C1 (n_1_98), .C2 (n_2_104) );
AOI211_X1 g_1_82 (.ZN (n_1_82), .A (n_1_86), .B (n_2_92), .C1 (n_2_96), .C2 (n_1_102) );
AOI211_X1 g_2_80 (.ZN (n_2_80), .A (n_2_84), .B (n_1_90), .C1 (n_1_94), .C2 (n_2_100) );
AOI211_X1 g_1_78 (.ZN (n_1_78), .A (n_1_82), .B (n_2_88), .C1 (n_2_92), .C2 (n_1_98) );
AOI211_X1 g_2_76 (.ZN (n_2_76), .A (n_2_80), .B (n_1_86), .C1 (n_1_90), .C2 (n_2_96) );
AOI211_X1 g_1_74 (.ZN (n_1_74), .A (n_1_78), .B (n_2_84), .C1 (n_2_88), .C2 (n_1_94) );
AOI211_X1 g_2_72 (.ZN (n_2_72), .A (n_2_76), .B (n_1_82), .C1 (n_1_86), .C2 (n_2_92) );
AOI211_X1 g_1_70 (.ZN (n_1_70), .A (n_1_74), .B (n_2_80), .C1 (n_2_84), .C2 (n_1_90) );
AOI211_X1 g_2_68 (.ZN (n_2_68), .A (n_2_72), .B (n_1_78), .C1 (n_1_82), .C2 (n_2_88) );
AOI211_X1 g_1_66 (.ZN (n_1_66), .A (n_1_70), .B (n_2_76), .C1 (n_2_80), .C2 (n_1_86) );
AOI211_X1 g_2_64 (.ZN (n_2_64), .A (n_2_68), .B (n_1_74), .C1 (n_1_78), .C2 (n_2_84) );
AOI211_X1 g_1_62 (.ZN (n_1_62), .A (n_1_66), .B (n_2_72), .C1 (n_2_76), .C2 (n_1_82) );
AOI211_X1 g_2_60 (.ZN (n_2_60), .A (n_2_64), .B (n_1_70), .C1 (n_1_74), .C2 (n_2_80) );
AOI211_X1 g_1_58 (.ZN (n_1_58), .A (n_1_62), .B (n_2_68), .C1 (n_2_72), .C2 (n_1_78) );
AOI211_X1 g_2_56 (.ZN (n_2_56), .A (n_2_60), .B (n_1_66), .C1 (n_1_70), .C2 (n_2_76) );
AOI211_X1 g_1_54 (.ZN (n_1_54), .A (n_1_58), .B (n_2_64), .C1 (n_2_68), .C2 (n_1_74) );
AOI211_X1 g_2_52 (.ZN (n_2_52), .A (n_2_56), .B (n_1_62), .C1 (n_1_66), .C2 (n_2_72) );
AOI211_X1 g_1_50 (.ZN (n_1_50), .A (n_1_54), .B (n_2_60), .C1 (n_2_64), .C2 (n_1_70) );
AOI211_X1 g_2_48 (.ZN (n_2_48), .A (n_2_52), .B (n_1_58), .C1 (n_1_62), .C2 (n_2_68) );
AOI211_X1 g_1_46 (.ZN (n_1_46), .A (n_1_50), .B (n_2_56), .C1 (n_2_60), .C2 (n_1_66) );
AOI211_X1 g_2_44 (.ZN (n_2_44), .A (n_2_48), .B (n_1_54), .C1 (n_1_58), .C2 (n_2_64) );
AOI211_X1 g_1_42 (.ZN (n_1_42), .A (n_1_46), .B (n_2_52), .C1 (n_2_56), .C2 (n_1_62) );
AOI211_X1 g_2_40 (.ZN (n_2_40), .A (n_2_44), .B (n_1_50), .C1 (n_1_54), .C2 (n_2_60) );
AOI211_X1 g_1_38 (.ZN (n_1_38), .A (n_1_42), .B (n_2_48), .C1 (n_2_52), .C2 (n_1_58) );
AOI211_X1 g_2_36 (.ZN (n_2_36), .A (n_2_40), .B (n_1_46), .C1 (n_1_50), .C2 (n_2_56) );
AOI211_X1 g_1_34 (.ZN (n_1_34), .A (n_1_38), .B (n_2_44), .C1 (n_2_48), .C2 (n_1_54) );
AOI211_X1 g_2_32 (.ZN (n_2_32), .A (n_2_36), .B (n_1_42), .C1 (n_1_46), .C2 (n_2_52) );
AOI211_X1 g_1_30 (.ZN (n_1_30), .A (n_1_34), .B (n_2_40), .C1 (n_2_44), .C2 (n_1_50) );
AOI211_X1 g_2_28 (.ZN (n_2_28), .A (n_2_32), .B (n_1_38), .C1 (n_1_42), .C2 (n_2_48) );
AOI211_X1 g_1_26 (.ZN (n_1_26), .A (n_1_30), .B (n_2_36), .C1 (n_2_40), .C2 (n_1_46) );
AOI211_X1 g_2_24 (.ZN (n_2_24), .A (n_2_28), .B (n_1_34), .C1 (n_1_38), .C2 (n_2_44) );
AOI211_X1 g_1_22 (.ZN (n_1_22), .A (n_1_26), .B (n_2_32), .C1 (n_2_36), .C2 (n_1_42) );
AOI211_X1 g_2_20 (.ZN (n_2_20), .A (n_2_24), .B (n_1_30), .C1 (n_1_34), .C2 (n_2_40) );
AOI211_X1 g_1_18 (.ZN (n_1_18), .A (n_1_22), .B (n_2_28), .C1 (n_2_32), .C2 (n_1_38) );
AOI211_X1 g_2_16 (.ZN (n_2_16), .A (n_2_20), .B (n_1_26), .C1 (n_1_30), .C2 (n_2_36) );
AOI211_X1 g_1_14 (.ZN (n_1_14), .A (n_1_18), .B (n_2_24), .C1 (n_2_28), .C2 (n_1_34) );
AOI211_X1 g_2_12 (.ZN (n_2_12), .A (n_2_16), .B (n_1_22), .C1 (n_1_26), .C2 (n_2_32) );
AOI211_X1 g_1_10 (.ZN (n_1_10), .A (n_1_14), .B (n_2_20), .C1 (n_2_24), .C2 (n_1_30) );
AOI211_X1 g_2_8 (.ZN (n_2_8), .A (n_2_12), .B (n_1_18), .C1 (n_1_22), .C2 (n_2_28) );
AOI211_X1 g_1_6 (.ZN (n_1_6), .A (n_1_10), .B (n_2_16), .C1 (n_2_20), .C2 (n_1_26) );
AOI211_X1 g_2_4 (.ZN (n_2_4), .A (n_2_8), .B (n_1_14), .C1 (n_1_18), .C2 (n_2_24) );
AOI211_X1 g_1_2 (.ZN (n_1_2), .A (n_1_6), .B (n_2_12), .C1 (n_2_16), .C2 (n_1_22) );
AOI211_X1 g_3_1 (.ZN (n_3_1), .A (n_2_4), .B (n_1_10), .C1 (n_1_14), .C2 (n_2_20) );
AOI211_X1 g_2_3 (.ZN (n_2_3), .A (n_1_2), .B (n_2_8), .C1 (n_2_12), .C2 (n_1_18) );
AOI211_X1 g_1_1 (.ZN (n_1_1), .A (n_3_1), .B (n_1_6), .C1 (n_1_10), .C2 (n_2_16) );
AOI211_X1 g_3_2 (.ZN (n_3_2), .A (n_2_3), .B (n_2_4), .C1 (n_2_8), .C2 (n_1_14) );
AOI211_X1 g_5_1 (.ZN (n_5_1), .A (n_1_1), .B (n_1_2), .C1 (n_1_6), .C2 (n_2_12) );
AOI211_X1 g_4_3 (.ZN (n_4_3), .A (n_3_2), .B (n_3_1), .C1 (n_2_4), .C2 (n_1_10) );
AOI211_X1 g_2_2 (.ZN (n_2_2), .A (n_5_1), .B (n_2_3), .C1 (n_1_2), .C2 (n_2_8) );
AOI211_X1 g_4_1 (.ZN (n_4_1), .A (n_4_3), .B (n_1_1), .C1 (n_3_1), .C2 (n_1_6) );
AOI211_X1 g_6_2 (.ZN (n_6_2), .A (n_2_2), .B (n_3_2), .C1 (n_2_3), .C2 (n_2_4) );
AOI211_X1 g_8_1 (.ZN (n_8_1), .A (n_4_1), .B (n_5_1), .C1 (n_1_1), .C2 (n_1_2) );
AOI211_X1 g_7_3 (.ZN (n_7_3), .A (n_6_2), .B (n_4_3), .C1 (n_3_2), .C2 (n_3_1) );
AOI211_X1 g_6_1 (.ZN (n_6_1), .A (n_8_1), .B (n_2_2), .C1 (n_5_1), .C2 (n_2_3) );
AOI211_X1 g_4_2 (.ZN (n_4_2), .A (n_7_3), .B (n_4_1), .C1 (n_4_3), .C2 (n_1_1) );
AOI211_X1 g_2_1 (.ZN (n_2_1), .A (n_6_1), .B (n_6_2), .C1 (n_2_2), .C2 (n_3_2) );
AOI211_X1 g_1_3 (.ZN (n_1_3), .A (n_4_2), .B (n_8_1), .C1 (n_4_1), .C2 (n_5_1) );
AOI211_X1 g_2_5 (.ZN (n_2_5), .A (n_2_1), .B (n_7_3), .C1 (n_6_2), .C2 (n_4_3) );
AOI211_X1 g_3_3 (.ZN (n_3_3), .A (n_1_3), .B (n_6_1), .C1 (n_8_1), .C2 (n_2_2) );
AOI211_X1 g_1_4 (.ZN (n_1_4), .A (n_2_5), .B (n_4_2), .C1 (n_7_3), .C2 (n_4_1) );
AOI211_X1 g_3_5 (.ZN (n_3_5), .A (n_3_3), .B (n_2_1), .C1 (n_6_1), .C2 (n_6_2) );
AOI211_X1 g_5_4 (.ZN (n_5_4), .A (n_1_4), .B (n_1_3), .C1 (n_4_2), .C2 (n_8_1) );
AOI211_X1 g_4_6 (.ZN (n_4_6), .A (n_3_5), .B (n_2_5), .C1 (n_2_1), .C2 (n_7_3) );
AOI211_X1 g_3_4 (.ZN (n_3_4), .A (n_5_4), .B (n_3_3), .C1 (n_1_3), .C2 (n_6_1) );
AOI211_X1 g_1_5 (.ZN (n_1_5), .A (n_4_6), .B (n_1_4), .C1 (n_2_5), .C2 (n_4_2) );
AOI211_X1 g_2_7 (.ZN (n_2_7), .A (n_3_4), .B (n_3_5), .C1 (n_3_3), .C2 (n_2_1) );
AOI211_X1 g_1_9 (.ZN (n_1_9), .A (n_1_5), .B (n_5_4), .C1 (n_1_4), .C2 (n_1_3) );
AOI211_X1 g_2_11 (.ZN (n_2_11), .A (n_2_7), .B (n_4_6), .C1 (n_3_5), .C2 (n_2_5) );
AOI211_X1 g_1_13 (.ZN (n_1_13), .A (n_1_9), .B (n_3_4), .C1 (n_5_4), .C2 (n_3_3) );
AOI211_X1 g_2_15 (.ZN (n_2_15), .A (n_2_11), .B (n_1_5), .C1 (n_4_6), .C2 (n_1_4) );
AOI211_X1 g_1_17 (.ZN (n_1_17), .A (n_1_13), .B (n_2_7), .C1 (n_3_4), .C2 (n_3_5) );
AOI211_X1 g_2_19 (.ZN (n_2_19), .A (n_2_15), .B (n_1_9), .C1 (n_1_5), .C2 (n_5_4) );
AOI211_X1 g_1_21 (.ZN (n_1_21), .A (n_1_17), .B (n_2_11), .C1 (n_2_7), .C2 (n_4_6) );
AOI211_X1 g_2_23 (.ZN (n_2_23), .A (n_2_19), .B (n_1_13), .C1 (n_1_9), .C2 (n_3_4) );
AOI211_X1 g_1_25 (.ZN (n_1_25), .A (n_1_21), .B (n_2_15), .C1 (n_2_11), .C2 (n_1_5) );
AOI211_X1 g_2_27 (.ZN (n_2_27), .A (n_2_23), .B (n_1_17), .C1 (n_1_13), .C2 (n_2_7) );
AOI211_X1 g_1_29 (.ZN (n_1_29), .A (n_1_25), .B (n_2_19), .C1 (n_2_15), .C2 (n_1_9) );
AOI211_X1 g_2_31 (.ZN (n_2_31), .A (n_2_27), .B (n_1_21), .C1 (n_1_17), .C2 (n_2_11) );
AOI211_X1 g_1_33 (.ZN (n_1_33), .A (n_1_29), .B (n_2_23), .C1 (n_2_19), .C2 (n_1_13) );
AOI211_X1 g_2_35 (.ZN (n_2_35), .A (n_2_31), .B (n_1_25), .C1 (n_1_21), .C2 (n_2_15) );
AOI211_X1 g_1_37 (.ZN (n_1_37), .A (n_1_33), .B (n_2_27), .C1 (n_2_23), .C2 (n_1_17) );
AOI211_X1 g_2_39 (.ZN (n_2_39), .A (n_2_35), .B (n_1_29), .C1 (n_1_25), .C2 (n_2_19) );
AOI211_X1 g_1_41 (.ZN (n_1_41), .A (n_1_37), .B (n_2_31), .C1 (n_2_27), .C2 (n_1_21) );
AOI211_X1 g_2_43 (.ZN (n_2_43), .A (n_2_39), .B (n_1_33), .C1 (n_1_29), .C2 (n_2_23) );
AOI211_X1 g_1_45 (.ZN (n_1_45), .A (n_1_41), .B (n_2_35), .C1 (n_2_31), .C2 (n_1_25) );
AOI211_X1 g_2_47 (.ZN (n_2_47), .A (n_2_43), .B (n_1_37), .C1 (n_1_33), .C2 (n_2_27) );
AOI211_X1 g_1_49 (.ZN (n_1_49), .A (n_1_45), .B (n_2_39), .C1 (n_2_35), .C2 (n_1_29) );
AOI211_X1 g_2_51 (.ZN (n_2_51), .A (n_2_47), .B (n_1_41), .C1 (n_1_37), .C2 (n_2_31) );
AOI211_X1 g_1_53 (.ZN (n_1_53), .A (n_1_49), .B (n_2_43), .C1 (n_2_39), .C2 (n_1_33) );
AOI211_X1 g_2_55 (.ZN (n_2_55), .A (n_2_51), .B (n_1_45), .C1 (n_1_41), .C2 (n_2_35) );
AOI211_X1 g_1_57 (.ZN (n_1_57), .A (n_1_53), .B (n_2_47), .C1 (n_2_43), .C2 (n_1_37) );
AOI211_X1 g_2_59 (.ZN (n_2_59), .A (n_2_55), .B (n_1_49), .C1 (n_1_45), .C2 (n_2_39) );
AOI211_X1 g_1_61 (.ZN (n_1_61), .A (n_1_57), .B (n_2_51), .C1 (n_2_47), .C2 (n_1_41) );
AOI211_X1 g_2_63 (.ZN (n_2_63), .A (n_2_59), .B (n_1_53), .C1 (n_1_49), .C2 (n_2_43) );
AOI211_X1 g_1_65 (.ZN (n_1_65), .A (n_1_61), .B (n_2_55), .C1 (n_2_51), .C2 (n_1_45) );
AOI211_X1 g_2_67 (.ZN (n_2_67), .A (n_2_63), .B (n_1_57), .C1 (n_1_53), .C2 (n_2_47) );
AOI211_X1 g_1_69 (.ZN (n_1_69), .A (n_1_65), .B (n_2_59), .C1 (n_2_55), .C2 (n_1_49) );
AOI211_X1 g_2_71 (.ZN (n_2_71), .A (n_2_67), .B (n_1_61), .C1 (n_1_57), .C2 (n_2_51) );
AOI211_X1 g_1_73 (.ZN (n_1_73), .A (n_1_69), .B (n_2_63), .C1 (n_2_59), .C2 (n_1_53) );
AOI211_X1 g_2_75 (.ZN (n_2_75), .A (n_2_71), .B (n_1_65), .C1 (n_1_61), .C2 (n_2_55) );
AOI211_X1 g_1_77 (.ZN (n_1_77), .A (n_1_73), .B (n_2_67), .C1 (n_2_63), .C2 (n_1_57) );
AOI211_X1 g_2_79 (.ZN (n_2_79), .A (n_2_75), .B (n_1_69), .C1 (n_1_65), .C2 (n_2_59) );
AOI211_X1 g_1_81 (.ZN (n_1_81), .A (n_1_77), .B (n_2_71), .C1 (n_2_67), .C2 (n_1_61) );
AOI211_X1 g_2_83 (.ZN (n_2_83), .A (n_2_79), .B (n_1_73), .C1 (n_1_69), .C2 (n_2_63) );
AOI211_X1 g_1_85 (.ZN (n_1_85), .A (n_1_81), .B (n_2_75), .C1 (n_2_71), .C2 (n_1_65) );
AOI211_X1 g_2_87 (.ZN (n_2_87), .A (n_2_83), .B (n_1_77), .C1 (n_1_73), .C2 (n_2_67) );
AOI211_X1 g_1_89 (.ZN (n_1_89), .A (n_1_85), .B (n_2_79), .C1 (n_2_75), .C2 (n_1_69) );
AOI211_X1 g_2_91 (.ZN (n_2_91), .A (n_2_87), .B (n_1_81), .C1 (n_1_77), .C2 (n_2_71) );
AOI211_X1 g_1_93 (.ZN (n_1_93), .A (n_1_89), .B (n_2_83), .C1 (n_2_79), .C2 (n_1_73) );
AOI211_X1 g_2_95 (.ZN (n_2_95), .A (n_2_91), .B (n_1_85), .C1 (n_1_81), .C2 (n_2_75) );
AOI211_X1 g_1_97 (.ZN (n_1_97), .A (n_1_93), .B (n_2_87), .C1 (n_2_83), .C2 (n_1_77) );
AOI211_X1 g_2_99 (.ZN (n_2_99), .A (n_2_95), .B (n_1_89), .C1 (n_1_85), .C2 (n_2_79) );
AOI211_X1 g_1_101 (.ZN (n_1_101), .A (n_1_97), .B (n_2_91), .C1 (n_2_87), .C2 (n_1_81) );
AOI211_X1 g_2_103 (.ZN (n_2_103), .A (n_2_99), .B (n_1_93), .C1 (n_1_89), .C2 (n_2_83) );
AOI211_X1 g_1_105 (.ZN (n_1_105), .A (n_1_101), .B (n_2_95), .C1 (n_2_91), .C2 (n_1_85) );
AOI211_X1 g_2_107 (.ZN (n_2_107), .A (n_2_103), .B (n_1_97), .C1 (n_1_93), .C2 (n_2_87) );
AOI211_X1 g_1_109 (.ZN (n_1_109), .A (n_1_105), .B (n_2_99), .C1 (n_2_95), .C2 (n_1_89) );
AOI211_X1 g_2_111 (.ZN (n_2_111), .A (n_2_107), .B (n_1_101), .C1 (n_1_97), .C2 (n_2_91) );
AOI211_X1 g_1_113 (.ZN (n_1_113), .A (n_1_109), .B (n_2_103), .C1 (n_2_99), .C2 (n_1_93) );
AOI211_X1 g_2_115 (.ZN (n_2_115), .A (n_2_111), .B (n_1_105), .C1 (n_1_101), .C2 (n_2_95) );
AOI211_X1 g_1_117 (.ZN (n_1_117), .A (n_1_113), .B (n_2_107), .C1 (n_2_103), .C2 (n_1_97) );
AOI211_X1 g_2_119 (.ZN (n_2_119), .A (n_2_115), .B (n_1_109), .C1 (n_1_105), .C2 (n_2_99) );
AOI211_X1 g_1_121 (.ZN (n_1_121), .A (n_1_117), .B (n_2_111), .C1 (n_2_107), .C2 (n_1_101) );
AOI211_X1 g_2_123 (.ZN (n_2_123), .A (n_2_119), .B (n_1_113), .C1 (n_1_109), .C2 (n_2_103) );
AOI211_X1 g_1_125 (.ZN (n_1_125), .A (n_1_121), .B (n_2_115), .C1 (n_2_111), .C2 (n_1_105) );
AOI211_X1 g_2_127 (.ZN (n_2_127), .A (n_2_123), .B (n_1_117), .C1 (n_1_113), .C2 (n_2_107) );
AOI211_X1 g_1_129 (.ZN (n_1_129), .A (n_1_125), .B (n_2_119), .C1 (n_2_115), .C2 (n_1_109) );
AOI211_X1 g_2_131 (.ZN (n_2_131), .A (n_2_127), .B (n_1_121), .C1 (n_1_117), .C2 (n_2_111) );
AOI211_X1 g_1_133 (.ZN (n_1_133), .A (n_1_129), .B (n_2_123), .C1 (n_2_119), .C2 (n_1_113) );
AOI211_X1 g_2_135 (.ZN (n_2_135), .A (n_2_131), .B (n_1_125), .C1 (n_1_121), .C2 (n_2_115) );
AOI211_X1 g_1_137 (.ZN (n_1_137), .A (n_1_133), .B (n_2_127), .C1 (n_2_123), .C2 (n_1_117) );
AOI211_X1 g_2_139 (.ZN (n_2_139), .A (n_2_135), .B (n_1_129), .C1 (n_1_125), .C2 (n_2_119) );
AOI211_X1 g_1_141 (.ZN (n_1_141), .A (n_1_137), .B (n_2_131), .C1 (n_2_127), .C2 (n_1_121) );
AOI211_X1 g_2_143 (.ZN (n_2_143), .A (n_2_139), .B (n_1_133), .C1 (n_1_129), .C2 (n_2_123) );
AOI211_X1 g_1_145 (.ZN (n_1_145), .A (n_1_141), .B (n_2_135), .C1 (n_2_131), .C2 (n_1_125) );
AOI211_X1 g_2_147 (.ZN (n_2_147), .A (n_2_143), .B (n_1_137), .C1 (n_1_133), .C2 (n_2_127) );
AOI211_X1 g_1_149 (.ZN (n_1_149), .A (n_1_145), .B (n_2_139), .C1 (n_2_135), .C2 (n_1_129) );
AOI211_X1 g_3_150 (.ZN (n_3_150), .A (n_2_147), .B (n_1_141), .C1 (n_1_137), .C2 (n_2_131) );
AOI211_X1 g_5_149 (.ZN (n_5_149), .A (n_1_149), .B (n_2_143), .C1 (n_2_139), .C2 (n_1_133) );
AOI211_X1 g_7_150 (.ZN (n_7_150), .A (n_3_150), .B (n_1_145), .C1 (n_1_141), .C2 (n_2_135) );
AOI211_X1 g_9_149 (.ZN (n_9_149), .A (n_5_149), .B (n_2_147), .C1 (n_2_143), .C2 (n_1_137) );
AOI211_X1 g_11_150 (.ZN (n_11_150), .A (n_7_150), .B (n_1_149), .C1 (n_1_145), .C2 (n_2_139) );
AOI211_X1 g_13_149 (.ZN (n_13_149), .A (n_9_149), .B (n_3_150), .C1 (n_2_147), .C2 (n_1_141) );
AOI211_X1 g_15_150 (.ZN (n_15_150), .A (n_11_150), .B (n_5_149), .C1 (n_1_149), .C2 (n_2_143) );
AOI211_X1 g_17_149 (.ZN (n_17_149), .A (n_13_149), .B (n_7_150), .C1 (n_3_150), .C2 (n_1_145) );
AOI211_X1 g_19_150 (.ZN (n_19_150), .A (n_15_150), .B (n_9_149), .C1 (n_5_149), .C2 (n_2_147) );
AOI211_X1 g_21_149 (.ZN (n_21_149), .A (n_17_149), .B (n_11_150), .C1 (n_7_150), .C2 (n_1_149) );
AOI211_X1 g_23_150 (.ZN (n_23_150), .A (n_19_150), .B (n_13_149), .C1 (n_9_149), .C2 (n_3_150) );
AOI211_X1 g_25_149 (.ZN (n_25_149), .A (n_21_149), .B (n_15_150), .C1 (n_11_150), .C2 (n_5_149) );
AOI211_X1 g_27_150 (.ZN (n_27_150), .A (n_23_150), .B (n_17_149), .C1 (n_13_149), .C2 (n_7_150) );
AOI211_X1 g_29_149 (.ZN (n_29_149), .A (n_25_149), .B (n_19_150), .C1 (n_15_150), .C2 (n_9_149) );
AOI211_X1 g_31_150 (.ZN (n_31_150), .A (n_27_150), .B (n_21_149), .C1 (n_17_149), .C2 (n_11_150) );
AOI211_X1 g_33_149 (.ZN (n_33_149), .A (n_29_149), .B (n_23_150), .C1 (n_19_150), .C2 (n_13_149) );
AOI211_X1 g_35_150 (.ZN (n_35_150), .A (n_31_150), .B (n_25_149), .C1 (n_21_149), .C2 (n_15_150) );
AOI211_X1 g_37_149 (.ZN (n_37_149), .A (n_33_149), .B (n_27_150), .C1 (n_23_150), .C2 (n_17_149) );
AOI211_X1 g_39_150 (.ZN (n_39_150), .A (n_35_150), .B (n_29_149), .C1 (n_25_149), .C2 (n_19_150) );
AOI211_X1 g_41_149 (.ZN (n_41_149), .A (n_37_149), .B (n_31_150), .C1 (n_27_150), .C2 (n_21_149) );
AOI211_X1 g_43_150 (.ZN (n_43_150), .A (n_39_150), .B (n_33_149), .C1 (n_29_149), .C2 (n_23_150) );
AOI211_X1 g_45_149 (.ZN (n_45_149), .A (n_41_149), .B (n_35_150), .C1 (n_31_150), .C2 (n_25_149) );
AOI211_X1 g_47_150 (.ZN (n_47_150), .A (n_43_150), .B (n_37_149), .C1 (n_33_149), .C2 (n_27_150) );
AOI211_X1 g_49_149 (.ZN (n_49_149), .A (n_45_149), .B (n_39_150), .C1 (n_35_150), .C2 (n_29_149) );
AOI211_X1 g_51_150 (.ZN (n_51_150), .A (n_47_150), .B (n_41_149), .C1 (n_37_149), .C2 (n_31_150) );
AOI211_X1 g_53_149 (.ZN (n_53_149), .A (n_49_149), .B (n_43_150), .C1 (n_39_150), .C2 (n_33_149) );
AOI211_X1 g_55_150 (.ZN (n_55_150), .A (n_51_150), .B (n_45_149), .C1 (n_41_149), .C2 (n_35_150) );
AOI211_X1 g_57_149 (.ZN (n_57_149), .A (n_53_149), .B (n_47_150), .C1 (n_43_150), .C2 (n_37_149) );
AOI211_X1 g_59_150 (.ZN (n_59_150), .A (n_55_150), .B (n_49_149), .C1 (n_45_149), .C2 (n_39_150) );
AOI211_X1 g_61_149 (.ZN (n_61_149), .A (n_57_149), .B (n_51_150), .C1 (n_47_150), .C2 (n_41_149) );
AOI211_X1 g_63_150 (.ZN (n_63_150), .A (n_59_150), .B (n_53_149), .C1 (n_49_149), .C2 (n_43_150) );
AOI211_X1 g_65_149 (.ZN (n_65_149), .A (n_61_149), .B (n_55_150), .C1 (n_51_150), .C2 (n_45_149) );
AOI211_X1 g_67_150 (.ZN (n_67_150), .A (n_63_150), .B (n_57_149), .C1 (n_53_149), .C2 (n_47_150) );
AOI211_X1 g_69_149 (.ZN (n_69_149), .A (n_65_149), .B (n_59_150), .C1 (n_55_150), .C2 (n_49_149) );
AOI211_X1 g_71_150 (.ZN (n_71_150), .A (n_67_150), .B (n_61_149), .C1 (n_57_149), .C2 (n_51_150) );
AOI211_X1 g_73_149 (.ZN (n_73_149), .A (n_69_149), .B (n_63_150), .C1 (n_59_150), .C2 (n_53_149) );
AOI211_X1 g_75_150 (.ZN (n_75_150), .A (n_71_150), .B (n_65_149), .C1 (n_61_149), .C2 (n_55_150) );
AOI211_X1 g_77_149 (.ZN (n_77_149), .A (n_73_149), .B (n_67_150), .C1 (n_63_150), .C2 (n_57_149) );
AOI211_X1 g_79_150 (.ZN (n_79_150), .A (n_75_150), .B (n_69_149), .C1 (n_65_149), .C2 (n_59_150) );
AOI211_X1 g_81_149 (.ZN (n_81_149), .A (n_77_149), .B (n_71_150), .C1 (n_67_150), .C2 (n_61_149) );
AOI211_X1 g_83_150 (.ZN (n_83_150), .A (n_79_150), .B (n_73_149), .C1 (n_69_149), .C2 (n_63_150) );
AOI211_X1 g_85_149 (.ZN (n_85_149), .A (n_81_149), .B (n_75_150), .C1 (n_71_150), .C2 (n_65_149) );
AOI211_X1 g_87_150 (.ZN (n_87_150), .A (n_83_150), .B (n_77_149), .C1 (n_73_149), .C2 (n_67_150) );
AOI211_X1 g_89_149 (.ZN (n_89_149), .A (n_85_149), .B (n_79_150), .C1 (n_75_150), .C2 (n_69_149) );
AOI211_X1 g_91_150 (.ZN (n_91_150), .A (n_87_150), .B (n_81_149), .C1 (n_77_149), .C2 (n_71_150) );
AOI211_X1 g_93_149 (.ZN (n_93_149), .A (n_89_149), .B (n_83_150), .C1 (n_79_150), .C2 (n_73_149) );
AOI211_X1 g_95_150 (.ZN (n_95_150), .A (n_91_150), .B (n_85_149), .C1 (n_81_149), .C2 (n_75_150) );
AOI211_X1 g_97_149 (.ZN (n_97_149), .A (n_93_149), .B (n_87_150), .C1 (n_83_150), .C2 (n_77_149) );
AOI211_X1 g_99_150 (.ZN (n_99_150), .A (n_95_150), .B (n_89_149), .C1 (n_85_149), .C2 (n_79_150) );
AOI211_X1 g_101_149 (.ZN (n_101_149), .A (n_97_149), .B (n_91_150), .C1 (n_87_150), .C2 (n_81_149) );
AOI211_X1 g_103_150 (.ZN (n_103_150), .A (n_99_150), .B (n_93_149), .C1 (n_89_149), .C2 (n_83_150) );
AOI211_X1 g_105_149 (.ZN (n_105_149), .A (n_101_149), .B (n_95_150), .C1 (n_91_150), .C2 (n_85_149) );
AOI211_X1 g_107_150 (.ZN (n_107_150), .A (n_103_150), .B (n_97_149), .C1 (n_93_149), .C2 (n_87_150) );
AOI211_X1 g_109_149 (.ZN (n_109_149), .A (n_105_149), .B (n_99_150), .C1 (n_95_150), .C2 (n_89_149) );
AOI211_X1 g_111_150 (.ZN (n_111_150), .A (n_107_150), .B (n_101_149), .C1 (n_97_149), .C2 (n_91_150) );
AOI211_X1 g_113_149 (.ZN (n_113_149), .A (n_109_149), .B (n_103_150), .C1 (n_99_150), .C2 (n_93_149) );
AOI211_X1 g_115_150 (.ZN (n_115_150), .A (n_111_150), .B (n_105_149), .C1 (n_101_149), .C2 (n_95_150) );
AOI211_X1 g_117_149 (.ZN (n_117_149), .A (n_113_149), .B (n_107_150), .C1 (n_103_150), .C2 (n_97_149) );
AOI211_X1 g_119_150 (.ZN (n_119_150), .A (n_115_150), .B (n_109_149), .C1 (n_105_149), .C2 (n_99_150) );
AOI211_X1 g_121_149 (.ZN (n_121_149), .A (n_117_149), .B (n_111_150), .C1 (n_107_150), .C2 (n_101_149) );
AOI211_X1 g_123_150 (.ZN (n_123_150), .A (n_119_150), .B (n_113_149), .C1 (n_109_149), .C2 (n_103_150) );
AOI211_X1 g_125_149 (.ZN (n_125_149), .A (n_121_149), .B (n_115_150), .C1 (n_111_150), .C2 (n_105_149) );
AOI211_X1 g_127_150 (.ZN (n_127_150), .A (n_123_150), .B (n_117_149), .C1 (n_113_149), .C2 (n_107_150) );
AOI211_X1 g_129_149 (.ZN (n_129_149), .A (n_125_149), .B (n_119_150), .C1 (n_115_150), .C2 (n_109_149) );
AOI211_X1 g_131_150 (.ZN (n_131_150), .A (n_127_150), .B (n_121_149), .C1 (n_117_149), .C2 (n_111_150) );
AOI211_X1 g_133_149 (.ZN (n_133_149), .A (n_129_149), .B (n_123_150), .C1 (n_119_150), .C2 (n_113_149) );
AOI211_X1 g_135_150 (.ZN (n_135_150), .A (n_131_150), .B (n_125_149), .C1 (n_121_149), .C2 (n_115_150) );
AOI211_X1 g_137_149 (.ZN (n_137_149), .A (n_133_149), .B (n_127_150), .C1 (n_123_150), .C2 (n_117_149) );
AOI211_X1 g_139_150 (.ZN (n_139_150), .A (n_135_150), .B (n_129_149), .C1 (n_125_149), .C2 (n_119_150) );
AOI211_X1 g_141_149 (.ZN (n_141_149), .A (n_137_149), .B (n_131_150), .C1 (n_127_150), .C2 (n_121_149) );
AOI211_X1 g_143_150 (.ZN (n_143_150), .A (n_139_150), .B (n_133_149), .C1 (n_129_149), .C2 (n_123_150) );
AOI211_X1 g_145_149 (.ZN (n_145_149), .A (n_141_149), .B (n_135_150), .C1 (n_131_150), .C2 (n_125_149) );
AOI211_X1 g_147_150 (.ZN (n_147_150), .A (n_143_150), .B (n_137_149), .C1 (n_133_149), .C2 (n_127_150) );
AOI211_X1 g_149_149 (.ZN (n_149_149), .A (n_145_149), .B (n_139_150), .C1 (n_135_150), .C2 (n_129_149) );
AOI211_X1 g_150_147 (.ZN (n_150_147), .A (n_147_150), .B (n_141_149), .C1 (n_137_149), .C2 (n_131_150) );
AOI211_X1 g_148_148 (.ZN (n_148_148), .A (n_149_149), .B (n_143_150), .C1 (n_139_150), .C2 (n_133_149) );
AOI211_X1 g_150_149 (.ZN (n_150_149), .A (n_150_147), .B (n_145_149), .C1 (n_141_149), .C2 (n_135_150) );
AOI211_X1 g_148_150 (.ZN (n_148_150), .A (n_148_148), .B (n_147_150), .C1 (n_143_150), .C2 (n_137_149) );
AOI211_X1 g_149_148 (.ZN (n_149_148), .A (n_150_149), .B (n_149_149), .C1 (n_145_149), .C2 (n_139_150) );
AOI211_X1 g_150_150 (.ZN (n_150_150), .A (n_148_150), .B (n_150_147), .C1 (n_147_150), .C2 (n_141_149) );
AOI211_X1 g_148_149 (.ZN (n_148_149), .A (n_149_148), .B (n_148_148), .C1 (n_149_149), .C2 (n_143_150) );
AOI211_X1 g_146_150 (.ZN (n_146_150), .A (n_150_150), .B (n_150_149), .C1 (n_150_147), .C2 (n_145_149) );
AOI211_X1 g_147_148 (.ZN (n_147_148), .A (n_148_149), .B (n_148_150), .C1 (n_148_148), .C2 (n_147_150) );
AOI211_X1 g_149_147 (.ZN (n_149_147), .A (n_146_150), .B (n_149_148), .C1 (n_150_149), .C2 (n_149_149) );
AOI211_X1 g_150_145 (.ZN (n_150_145), .A (n_147_148), .B (n_150_150), .C1 (n_148_150), .C2 (n_150_147) );
AOI211_X1 g_148_146 (.ZN (n_148_146), .A (n_149_147), .B (n_148_149), .C1 (n_149_148), .C2 (n_148_148) );
AOI211_X1 g_146_147 (.ZN (n_146_147), .A (n_150_145), .B (n_146_150), .C1 (n_150_150), .C2 (n_150_149) );
AOI211_X1 g_144_148 (.ZN (n_144_148), .A (n_148_146), .B (n_147_148), .C1 (n_148_149), .C2 (n_148_150) );
AOI211_X1 g_146_149 (.ZN (n_146_149), .A (n_146_147), .B (n_149_147), .C1 (n_146_150), .C2 (n_149_148) );
AOI211_X1 g_144_150 (.ZN (n_144_150), .A (n_144_148), .B (n_150_145), .C1 (n_147_148), .C2 (n_150_150) );
AOI211_X1 g_145_148 (.ZN (n_145_148), .A (n_146_149), .B (n_148_146), .C1 (n_149_147), .C2 (n_148_149) );
AOI211_X1 g_147_147 (.ZN (n_147_147), .A (n_144_150), .B (n_146_147), .C1 (n_150_145), .C2 (n_146_150) );
AOI211_X1 g_148_145 (.ZN (n_148_145), .A (n_145_148), .B (n_144_148), .C1 (n_148_146), .C2 (n_147_148) );
AOI211_X1 g_150_146 (.ZN (n_150_146), .A (n_147_147), .B (n_146_149), .C1 (n_146_147), .C2 (n_149_147) );
AOI211_X1 g_149_144 (.ZN (n_149_144), .A (n_148_145), .B (n_144_150), .C1 (n_144_148), .C2 (n_150_145) );
AOI211_X1 g_150_142 (.ZN (n_150_142), .A (n_150_146), .B (n_145_148), .C1 (n_146_149), .C2 (n_148_146) );
AOI211_X1 g_149_140 (.ZN (n_149_140), .A (n_149_144), .B (n_147_147), .C1 (n_144_150), .C2 (n_146_147) );
AOI211_X1 g_150_138 (.ZN (n_150_138), .A (n_150_142), .B (n_148_145), .C1 (n_145_148), .C2 (n_144_148) );
AOI211_X1 g_149_136 (.ZN (n_149_136), .A (n_149_140), .B (n_150_146), .C1 (n_147_147), .C2 (n_146_149) );
AOI211_X1 g_150_134 (.ZN (n_150_134), .A (n_150_138), .B (n_149_144), .C1 (n_148_145), .C2 (n_144_150) );
AOI211_X1 g_149_132 (.ZN (n_149_132), .A (n_149_136), .B (n_150_142), .C1 (n_150_146), .C2 (n_145_148) );
AOI211_X1 g_150_130 (.ZN (n_150_130), .A (n_150_134), .B (n_149_140), .C1 (n_149_144), .C2 (n_147_147) );
AOI211_X1 g_149_128 (.ZN (n_149_128), .A (n_149_132), .B (n_150_138), .C1 (n_150_142), .C2 (n_148_145) );
AOI211_X1 g_150_126 (.ZN (n_150_126), .A (n_150_130), .B (n_149_136), .C1 (n_149_140), .C2 (n_150_146) );
AOI211_X1 g_149_124 (.ZN (n_149_124), .A (n_149_128), .B (n_150_134), .C1 (n_150_138), .C2 (n_149_144) );
AOI211_X1 g_150_122 (.ZN (n_150_122), .A (n_150_126), .B (n_149_132), .C1 (n_149_136), .C2 (n_150_142) );
AOI211_X1 g_149_120 (.ZN (n_149_120), .A (n_149_124), .B (n_150_130), .C1 (n_150_134), .C2 (n_149_140) );
AOI211_X1 g_150_118 (.ZN (n_150_118), .A (n_150_122), .B (n_149_128), .C1 (n_149_132), .C2 (n_150_138) );
AOI211_X1 g_149_116 (.ZN (n_149_116), .A (n_149_120), .B (n_150_126), .C1 (n_150_130), .C2 (n_149_136) );
AOI211_X1 g_150_114 (.ZN (n_150_114), .A (n_150_118), .B (n_149_124), .C1 (n_149_128), .C2 (n_150_134) );
AOI211_X1 g_149_112 (.ZN (n_149_112), .A (n_149_116), .B (n_150_122), .C1 (n_150_126), .C2 (n_149_132) );
AOI211_X1 g_150_110 (.ZN (n_150_110), .A (n_150_114), .B (n_149_120), .C1 (n_149_124), .C2 (n_150_130) );
AOI211_X1 g_149_108 (.ZN (n_149_108), .A (n_149_112), .B (n_150_118), .C1 (n_150_122), .C2 (n_149_128) );
AOI211_X1 g_150_106 (.ZN (n_150_106), .A (n_150_110), .B (n_149_116), .C1 (n_149_120), .C2 (n_150_126) );
AOI211_X1 g_149_104 (.ZN (n_149_104), .A (n_149_108), .B (n_150_114), .C1 (n_150_118), .C2 (n_149_124) );
AOI211_X1 g_150_102 (.ZN (n_150_102), .A (n_150_106), .B (n_149_112), .C1 (n_149_116), .C2 (n_150_122) );
AOI211_X1 g_149_100 (.ZN (n_149_100), .A (n_149_104), .B (n_150_110), .C1 (n_150_114), .C2 (n_149_120) );
AOI211_X1 g_150_98 (.ZN (n_150_98), .A (n_150_102), .B (n_149_108), .C1 (n_149_112), .C2 (n_150_118) );
AOI211_X1 g_149_96 (.ZN (n_149_96), .A (n_149_100), .B (n_150_106), .C1 (n_150_110), .C2 (n_149_116) );
AOI211_X1 g_150_94 (.ZN (n_150_94), .A (n_150_98), .B (n_149_104), .C1 (n_149_108), .C2 (n_150_114) );
AOI211_X1 g_149_92 (.ZN (n_149_92), .A (n_149_96), .B (n_150_102), .C1 (n_150_106), .C2 (n_149_112) );
AOI211_X1 g_150_90 (.ZN (n_150_90), .A (n_150_94), .B (n_149_100), .C1 (n_149_104), .C2 (n_150_110) );
AOI211_X1 g_149_88 (.ZN (n_149_88), .A (n_149_92), .B (n_150_98), .C1 (n_150_102), .C2 (n_149_108) );
AOI211_X1 g_150_86 (.ZN (n_150_86), .A (n_150_90), .B (n_149_96), .C1 (n_149_100), .C2 (n_150_106) );
AOI211_X1 g_149_84 (.ZN (n_149_84), .A (n_149_88), .B (n_150_94), .C1 (n_150_98), .C2 (n_149_104) );
AOI211_X1 g_150_82 (.ZN (n_150_82), .A (n_150_86), .B (n_149_92), .C1 (n_149_96), .C2 (n_150_102) );
AOI211_X1 g_149_80 (.ZN (n_149_80), .A (n_149_84), .B (n_150_90), .C1 (n_150_94), .C2 (n_149_100) );
AOI211_X1 g_150_78 (.ZN (n_150_78), .A (n_150_82), .B (n_149_88), .C1 (n_149_92), .C2 (n_150_98) );
AOI211_X1 g_149_76 (.ZN (n_149_76), .A (n_149_80), .B (n_150_86), .C1 (n_150_90), .C2 (n_149_96) );
AOI211_X1 g_150_74 (.ZN (n_150_74), .A (n_150_78), .B (n_149_84), .C1 (n_149_88), .C2 (n_150_94) );
AOI211_X1 g_149_72 (.ZN (n_149_72), .A (n_149_76), .B (n_150_82), .C1 (n_150_86), .C2 (n_149_92) );
AOI211_X1 g_150_70 (.ZN (n_150_70), .A (n_150_74), .B (n_149_80), .C1 (n_149_84), .C2 (n_150_90) );
AOI211_X1 g_149_68 (.ZN (n_149_68), .A (n_149_72), .B (n_150_78), .C1 (n_150_82), .C2 (n_149_88) );
AOI211_X1 g_150_66 (.ZN (n_150_66), .A (n_150_70), .B (n_149_76), .C1 (n_149_80), .C2 (n_150_86) );
AOI211_X1 g_149_64 (.ZN (n_149_64), .A (n_149_68), .B (n_150_74), .C1 (n_150_78), .C2 (n_149_84) );
AOI211_X1 g_150_62 (.ZN (n_150_62), .A (n_150_66), .B (n_149_72), .C1 (n_149_76), .C2 (n_150_82) );
AOI211_X1 g_149_60 (.ZN (n_149_60), .A (n_149_64), .B (n_150_70), .C1 (n_150_74), .C2 (n_149_80) );
AOI211_X1 g_150_58 (.ZN (n_150_58), .A (n_150_62), .B (n_149_68), .C1 (n_149_72), .C2 (n_150_78) );
AOI211_X1 g_149_56 (.ZN (n_149_56), .A (n_149_60), .B (n_150_66), .C1 (n_150_70), .C2 (n_149_76) );
AOI211_X1 g_150_54 (.ZN (n_150_54), .A (n_150_58), .B (n_149_64), .C1 (n_149_68), .C2 (n_150_74) );
AOI211_X1 g_149_52 (.ZN (n_149_52), .A (n_149_56), .B (n_150_62), .C1 (n_150_66), .C2 (n_149_72) );
AOI211_X1 g_150_50 (.ZN (n_150_50), .A (n_150_54), .B (n_149_60), .C1 (n_149_64), .C2 (n_150_70) );
AOI211_X1 g_149_48 (.ZN (n_149_48), .A (n_149_52), .B (n_150_58), .C1 (n_150_62), .C2 (n_149_68) );
AOI211_X1 g_150_46 (.ZN (n_150_46), .A (n_150_50), .B (n_149_56), .C1 (n_149_60), .C2 (n_150_66) );
AOI211_X1 g_149_44 (.ZN (n_149_44), .A (n_149_48), .B (n_150_54), .C1 (n_150_58), .C2 (n_149_64) );
AOI211_X1 g_150_42 (.ZN (n_150_42), .A (n_150_46), .B (n_149_52), .C1 (n_149_56), .C2 (n_150_62) );
AOI211_X1 g_149_40 (.ZN (n_149_40), .A (n_149_44), .B (n_150_50), .C1 (n_150_54), .C2 (n_149_60) );
AOI211_X1 g_150_38 (.ZN (n_150_38), .A (n_150_42), .B (n_149_48), .C1 (n_149_52), .C2 (n_150_58) );
AOI211_X1 g_149_36 (.ZN (n_149_36), .A (n_149_40), .B (n_150_46), .C1 (n_150_50), .C2 (n_149_56) );
AOI211_X1 g_150_34 (.ZN (n_150_34), .A (n_150_38), .B (n_149_44), .C1 (n_149_48), .C2 (n_150_54) );
AOI211_X1 g_149_32 (.ZN (n_149_32), .A (n_149_36), .B (n_150_42), .C1 (n_150_46), .C2 (n_149_52) );
AOI211_X1 g_150_30 (.ZN (n_150_30), .A (n_150_34), .B (n_149_40), .C1 (n_149_44), .C2 (n_150_50) );
AOI211_X1 g_149_28 (.ZN (n_149_28), .A (n_149_32), .B (n_150_38), .C1 (n_150_42), .C2 (n_149_48) );
AOI211_X1 g_150_26 (.ZN (n_150_26), .A (n_150_30), .B (n_149_36), .C1 (n_149_40), .C2 (n_150_46) );
AOI211_X1 g_149_24 (.ZN (n_149_24), .A (n_149_28), .B (n_150_34), .C1 (n_150_38), .C2 (n_149_44) );
AOI211_X1 g_150_22 (.ZN (n_150_22), .A (n_150_26), .B (n_149_32), .C1 (n_149_36), .C2 (n_150_42) );
AOI211_X1 g_149_20 (.ZN (n_149_20), .A (n_149_24), .B (n_150_30), .C1 (n_150_34), .C2 (n_149_40) );
AOI211_X1 g_150_18 (.ZN (n_150_18), .A (n_150_22), .B (n_149_28), .C1 (n_149_32), .C2 (n_150_38) );
AOI211_X1 g_149_16 (.ZN (n_149_16), .A (n_149_20), .B (n_150_26), .C1 (n_150_30), .C2 (n_149_36) );
AOI211_X1 g_150_14 (.ZN (n_150_14), .A (n_150_18), .B (n_149_24), .C1 (n_149_28), .C2 (n_150_34) );
AOI211_X1 g_149_12 (.ZN (n_149_12), .A (n_149_16), .B (n_150_22), .C1 (n_150_26), .C2 (n_149_32) );
AOI211_X1 g_150_10 (.ZN (n_150_10), .A (n_150_14), .B (n_149_20), .C1 (n_149_24), .C2 (n_150_30) );
AOI211_X1 g_149_8 (.ZN (n_149_8), .A (n_149_12), .B (n_150_18), .C1 (n_150_22), .C2 (n_149_28) );
AOI211_X1 g_150_6 (.ZN (n_150_6), .A (n_150_10), .B (n_149_16), .C1 (n_149_20), .C2 (n_150_26) );
AOI211_X1 g_149_4 (.ZN (n_149_4), .A (n_149_8), .B (n_150_14), .C1 (n_150_18), .C2 (n_149_24) );
AOI211_X1 g_150_2 (.ZN (n_150_2), .A (n_150_6), .B (n_149_12), .C1 (n_149_16), .C2 (n_150_22) );
AOI211_X1 g_148_1 (.ZN (n_148_1), .A (n_149_4), .B (n_150_10), .C1 (n_150_14), .C2 (n_149_20) );
AOI211_X1 g_147_3 (.ZN (n_147_3), .A (n_150_2), .B (n_149_8), .C1 (n_149_12), .C2 (n_150_18) );
AOI211_X1 g_146_1 (.ZN (n_146_1), .A (n_148_1), .B (n_150_6), .C1 (n_150_10), .C2 (n_149_16) );
AOI211_X1 g_148_2 (.ZN (n_148_2), .A (n_147_3), .B (n_149_4), .C1 (n_149_8), .C2 (n_150_14) );
AOI211_X1 g_150_1 (.ZN (n_150_1), .A (n_146_1), .B (n_150_2), .C1 (n_150_6), .C2 (n_149_12) );
AOI211_X1 g_149_3 (.ZN (n_149_3), .A (n_148_2), .B (n_148_1), .C1 (n_149_4), .C2 (n_150_10) );
AOI211_X1 g_150_5 (.ZN (n_150_5), .A (n_150_1), .B (n_147_3), .C1 (n_150_2), .C2 (n_149_8) );
AOI211_X1 g_148_4 (.ZN (n_148_4), .A (n_149_3), .B (n_146_1), .C1 (n_148_1), .C2 (n_150_6) );
AOI211_X1 g_150_3 (.ZN (n_150_3), .A (n_150_5), .B (n_148_2), .C1 (n_147_3), .C2 (n_149_4) );
AOI211_X1 g_149_1 (.ZN (n_149_1), .A (n_148_4), .B (n_150_1), .C1 (n_146_1), .C2 (n_150_2) );
AOI211_X1 g_147_2 (.ZN (n_147_2), .A (n_150_3), .B (n_149_3), .C1 (n_148_2), .C2 (n_148_1) );
AOI211_X1 g_145_1 (.ZN (n_145_1), .A (n_149_1), .B (n_150_5), .C1 (n_150_1), .C2 (n_147_3) );
AOI211_X1 g_146_3 (.ZN (n_146_3), .A (n_147_2), .B (n_148_4), .C1 (n_149_3), .C2 (n_146_1) );
AOI211_X1 g_144_2 (.ZN (n_144_2), .A (n_145_1), .B (n_150_3), .C1 (n_150_5), .C2 (n_148_2) );
AOI211_X1 g_142_1 (.ZN (n_142_1), .A (n_146_3), .B (n_149_1), .C1 (n_148_4), .C2 (n_150_1) );
AOI211_X1 g_140_2 (.ZN (n_140_2), .A (n_144_2), .B (n_147_2), .C1 (n_150_3), .C2 (n_149_3) );
AOI211_X1 g_138_1 (.ZN (n_138_1), .A (n_142_1), .B (n_145_1), .C1 (n_149_1), .C2 (n_150_5) );
AOI211_X1 g_136_2 (.ZN (n_136_2), .A (n_140_2), .B (n_146_3), .C1 (n_147_2), .C2 (n_148_4) );
AOI211_X1 g_134_1 (.ZN (n_134_1), .A (n_138_1), .B (n_144_2), .C1 (n_145_1), .C2 (n_150_3) );
AOI211_X1 g_132_2 (.ZN (n_132_2), .A (n_136_2), .B (n_142_1), .C1 (n_146_3), .C2 (n_149_1) );
AOI211_X1 g_130_1 (.ZN (n_130_1), .A (n_134_1), .B (n_140_2), .C1 (n_144_2), .C2 (n_147_2) );
AOI211_X1 g_128_2 (.ZN (n_128_2), .A (n_132_2), .B (n_138_1), .C1 (n_142_1), .C2 (n_145_1) );
AOI211_X1 g_126_1 (.ZN (n_126_1), .A (n_130_1), .B (n_136_2), .C1 (n_140_2), .C2 (n_146_3) );
AOI211_X1 g_124_2 (.ZN (n_124_2), .A (n_128_2), .B (n_134_1), .C1 (n_138_1), .C2 (n_144_2) );
AOI211_X1 g_122_1 (.ZN (n_122_1), .A (n_126_1), .B (n_132_2), .C1 (n_136_2), .C2 (n_142_1) );
AOI211_X1 g_120_2 (.ZN (n_120_2), .A (n_124_2), .B (n_130_1), .C1 (n_134_1), .C2 (n_140_2) );
AOI211_X1 g_118_1 (.ZN (n_118_1), .A (n_122_1), .B (n_128_2), .C1 (n_132_2), .C2 (n_138_1) );
AOI211_X1 g_116_2 (.ZN (n_116_2), .A (n_120_2), .B (n_126_1), .C1 (n_130_1), .C2 (n_136_2) );
AOI211_X1 g_114_1 (.ZN (n_114_1), .A (n_118_1), .B (n_124_2), .C1 (n_128_2), .C2 (n_134_1) );
AOI211_X1 g_112_2 (.ZN (n_112_2), .A (n_116_2), .B (n_122_1), .C1 (n_126_1), .C2 (n_132_2) );
AOI211_X1 g_110_1 (.ZN (n_110_1), .A (n_114_1), .B (n_120_2), .C1 (n_124_2), .C2 (n_130_1) );
AOI211_X1 g_108_2 (.ZN (n_108_2), .A (n_112_2), .B (n_118_1), .C1 (n_122_1), .C2 (n_128_2) );
AOI211_X1 g_106_1 (.ZN (n_106_1), .A (n_110_1), .B (n_116_2), .C1 (n_120_2), .C2 (n_126_1) );
AOI211_X1 g_104_2 (.ZN (n_104_2), .A (n_108_2), .B (n_114_1), .C1 (n_118_1), .C2 (n_124_2) );
AOI211_X1 g_102_1 (.ZN (n_102_1), .A (n_106_1), .B (n_112_2), .C1 (n_116_2), .C2 (n_122_1) );
AOI211_X1 g_100_2 (.ZN (n_100_2), .A (n_104_2), .B (n_110_1), .C1 (n_114_1), .C2 (n_120_2) );
AOI211_X1 g_98_1 (.ZN (n_98_1), .A (n_102_1), .B (n_108_2), .C1 (n_112_2), .C2 (n_118_1) );
AOI211_X1 g_96_2 (.ZN (n_96_2), .A (n_100_2), .B (n_106_1), .C1 (n_110_1), .C2 (n_116_2) );
AOI211_X1 g_94_1 (.ZN (n_94_1), .A (n_98_1), .B (n_104_2), .C1 (n_108_2), .C2 (n_114_1) );
AOI211_X1 g_92_2 (.ZN (n_92_2), .A (n_96_2), .B (n_102_1), .C1 (n_106_1), .C2 (n_112_2) );
AOI211_X1 g_90_1 (.ZN (n_90_1), .A (n_94_1), .B (n_100_2), .C1 (n_104_2), .C2 (n_110_1) );
AOI211_X1 g_88_2 (.ZN (n_88_2), .A (n_92_2), .B (n_98_1), .C1 (n_102_1), .C2 (n_108_2) );
AOI211_X1 g_86_1 (.ZN (n_86_1), .A (n_90_1), .B (n_96_2), .C1 (n_100_2), .C2 (n_106_1) );
AOI211_X1 g_84_2 (.ZN (n_84_2), .A (n_88_2), .B (n_94_1), .C1 (n_98_1), .C2 (n_104_2) );
AOI211_X1 g_82_1 (.ZN (n_82_1), .A (n_86_1), .B (n_92_2), .C1 (n_96_2), .C2 (n_102_1) );
AOI211_X1 g_80_2 (.ZN (n_80_2), .A (n_84_2), .B (n_90_1), .C1 (n_94_1), .C2 (n_100_2) );
AOI211_X1 g_78_1 (.ZN (n_78_1), .A (n_82_1), .B (n_88_2), .C1 (n_92_2), .C2 (n_98_1) );
AOI211_X1 g_76_2 (.ZN (n_76_2), .A (n_80_2), .B (n_86_1), .C1 (n_90_1), .C2 (n_96_2) );
AOI211_X1 g_74_1 (.ZN (n_74_1), .A (n_78_1), .B (n_84_2), .C1 (n_88_2), .C2 (n_94_1) );
AOI211_X1 g_72_2 (.ZN (n_72_2), .A (n_76_2), .B (n_82_1), .C1 (n_86_1), .C2 (n_92_2) );
AOI211_X1 g_70_1 (.ZN (n_70_1), .A (n_74_1), .B (n_80_2), .C1 (n_84_2), .C2 (n_90_1) );
AOI211_X1 g_68_2 (.ZN (n_68_2), .A (n_72_2), .B (n_78_1), .C1 (n_82_1), .C2 (n_88_2) );
AOI211_X1 g_66_1 (.ZN (n_66_1), .A (n_70_1), .B (n_76_2), .C1 (n_80_2), .C2 (n_86_1) );
AOI211_X1 g_64_2 (.ZN (n_64_2), .A (n_68_2), .B (n_74_1), .C1 (n_78_1), .C2 (n_84_2) );
AOI211_X1 g_62_1 (.ZN (n_62_1), .A (n_66_1), .B (n_72_2), .C1 (n_76_2), .C2 (n_82_1) );
AOI211_X1 g_60_2 (.ZN (n_60_2), .A (n_64_2), .B (n_70_1), .C1 (n_74_1), .C2 (n_80_2) );
AOI211_X1 g_58_1 (.ZN (n_58_1), .A (n_62_1), .B (n_68_2), .C1 (n_72_2), .C2 (n_78_1) );
AOI211_X1 g_56_2 (.ZN (n_56_2), .A (n_60_2), .B (n_66_1), .C1 (n_70_1), .C2 (n_76_2) );
AOI211_X1 g_54_1 (.ZN (n_54_1), .A (n_58_1), .B (n_64_2), .C1 (n_68_2), .C2 (n_74_1) );
AOI211_X1 g_52_2 (.ZN (n_52_2), .A (n_56_2), .B (n_62_1), .C1 (n_66_1), .C2 (n_72_2) );
AOI211_X1 g_50_1 (.ZN (n_50_1), .A (n_54_1), .B (n_60_2), .C1 (n_64_2), .C2 (n_70_1) );
AOI211_X1 g_48_2 (.ZN (n_48_2), .A (n_52_2), .B (n_58_1), .C1 (n_62_1), .C2 (n_68_2) );
AOI211_X1 g_46_1 (.ZN (n_46_1), .A (n_50_1), .B (n_56_2), .C1 (n_60_2), .C2 (n_66_1) );
AOI211_X1 g_44_2 (.ZN (n_44_2), .A (n_48_2), .B (n_54_1), .C1 (n_58_1), .C2 (n_64_2) );
AOI211_X1 g_42_1 (.ZN (n_42_1), .A (n_46_1), .B (n_52_2), .C1 (n_56_2), .C2 (n_62_1) );
AOI211_X1 g_40_2 (.ZN (n_40_2), .A (n_44_2), .B (n_50_1), .C1 (n_54_1), .C2 (n_60_2) );
AOI211_X1 g_38_1 (.ZN (n_38_1), .A (n_42_1), .B (n_48_2), .C1 (n_52_2), .C2 (n_58_1) );
AOI211_X1 g_36_2 (.ZN (n_36_2), .A (n_40_2), .B (n_46_1), .C1 (n_50_1), .C2 (n_56_2) );
AOI211_X1 g_34_1 (.ZN (n_34_1), .A (n_38_1), .B (n_44_2), .C1 (n_48_2), .C2 (n_54_1) );
AOI211_X1 g_32_2 (.ZN (n_32_2), .A (n_36_2), .B (n_42_1), .C1 (n_46_1), .C2 (n_52_2) );
AOI211_X1 g_30_1 (.ZN (n_30_1), .A (n_34_1), .B (n_40_2), .C1 (n_44_2), .C2 (n_50_1) );
AOI211_X1 g_28_2 (.ZN (n_28_2), .A (n_32_2), .B (n_38_1), .C1 (n_42_1), .C2 (n_48_2) );
AOI211_X1 g_26_1 (.ZN (n_26_1), .A (n_30_1), .B (n_36_2), .C1 (n_40_2), .C2 (n_46_1) );
AOI211_X1 g_24_2 (.ZN (n_24_2), .A (n_28_2), .B (n_34_1), .C1 (n_38_1), .C2 (n_44_2) );
AOI211_X1 g_22_1 (.ZN (n_22_1), .A (n_26_1), .B (n_32_2), .C1 (n_36_2), .C2 (n_42_1) );
AOI211_X1 g_20_2 (.ZN (n_20_2), .A (n_24_2), .B (n_30_1), .C1 (n_34_1), .C2 (n_40_2) );
AOI211_X1 g_18_1 (.ZN (n_18_1), .A (n_22_1), .B (n_28_2), .C1 (n_32_2), .C2 (n_38_1) );
AOI211_X1 g_16_2 (.ZN (n_16_2), .A (n_20_2), .B (n_26_1), .C1 (n_30_1), .C2 (n_36_2) );
AOI211_X1 g_14_1 (.ZN (n_14_1), .A (n_18_1), .B (n_24_2), .C1 (n_28_2), .C2 (n_34_1) );
AOI211_X1 g_12_2 (.ZN (n_12_2), .A (n_16_2), .B (n_22_1), .C1 (n_26_1), .C2 (n_32_2) );
AOI211_X1 g_10_1 (.ZN (n_10_1), .A (n_14_1), .B (n_20_2), .C1 (n_24_2), .C2 (n_30_1) );
AOI211_X1 g_8_2 (.ZN (n_8_2), .A (n_12_2), .B (n_18_1), .C1 (n_22_1), .C2 (n_28_2) );
AOI211_X1 g_6_3 (.ZN (n_6_3), .A (n_10_1), .B (n_16_2), .C1 (n_20_2), .C2 (n_26_1) );
AOI211_X1 g_5_5 (.ZN (n_5_5), .A (n_8_2), .B (n_14_1), .C1 (n_18_1), .C2 (n_24_2) );
AOI211_X1 g_3_6 (.ZN (n_3_6), .A (n_6_3), .B (n_12_2), .C1 (n_16_2), .C2 (n_22_1) );
AOI211_X1 g_1_7 (.ZN (n_1_7), .A (n_5_5), .B (n_10_1), .C1 (n_14_1), .C2 (n_20_2) );
AOI211_X1 g_2_9 (.ZN (n_2_9), .A (n_3_6), .B (n_8_2), .C1 (n_12_2), .C2 (n_18_1) );
AOI211_X1 g_1_11 (.ZN (n_1_11), .A (n_1_7), .B (n_6_3), .C1 (n_10_1), .C2 (n_16_2) );
AOI211_X1 g_3_10 (.ZN (n_3_10), .A (n_2_9), .B (n_5_5), .C1 (n_8_2), .C2 (n_14_1) );
AOI211_X1 g_4_8 (.ZN (n_4_8), .A (n_1_11), .B (n_3_6), .C1 (n_6_3), .C2 (n_12_2) );
AOI211_X1 g_6_7 (.ZN (n_6_7), .A (n_3_10), .B (n_1_7), .C1 (n_5_5), .C2 (n_10_1) );
AOI211_X1 g_7_5 (.ZN (n_7_5), .A (n_4_8), .B (n_2_9), .C1 (n_3_6), .C2 (n_8_2) );
AOI211_X1 g_5_6 (.ZN (n_5_6), .A (n_6_7), .B (n_1_11), .C1 (n_1_7), .C2 (n_6_3) );
AOI211_X1 g_3_7 (.ZN (n_3_7), .A (n_7_5), .B (n_3_10), .C1 (n_2_9), .C2 (n_5_5) );
AOI211_X1 g_1_8 (.ZN (n_1_8), .A (n_5_6), .B (n_4_8), .C1 (n_1_11), .C2 (n_3_6) );
AOI211_X1 g_2_6 (.ZN (n_2_6), .A (n_3_7), .B (n_6_7), .C1 (n_3_10), .C2 (n_1_7) );
AOI211_X1 g_4_5 (.ZN (n_4_5), .A (n_1_8), .B (n_7_5), .C1 (n_4_8), .C2 (n_2_9) );
AOI211_X1 g_5_3 (.ZN (n_5_3), .A (n_2_6), .B (n_5_6), .C1 (n_6_7), .C2 (n_1_11) );
AOI211_X1 g_7_2 (.ZN (n_7_2), .A (n_4_5), .B (n_3_7), .C1 (n_7_5), .C2 (n_3_10) );
AOI211_X1 g_9_1 (.ZN (n_9_1), .A (n_5_3), .B (n_1_8), .C1 (n_5_6), .C2 (n_4_8) );
AOI211_X1 g_8_3 (.ZN (n_8_3), .A (n_7_2), .B (n_2_6), .C1 (n_3_7), .C2 (n_6_7) );
AOI211_X1 g_6_4 (.ZN (n_6_4), .A (n_9_1), .B (n_4_5), .C1 (n_1_8), .C2 (n_7_5) );
AOI211_X1 g_7_6 (.ZN (n_7_6), .A (n_8_3), .B (n_5_3), .C1 (n_2_6), .C2 (n_5_6) );
AOI211_X1 g_8_4 (.ZN (n_8_4), .A (n_6_4), .B (n_7_2), .C1 (n_4_5), .C2 (n_3_7) );
AOI211_X1 g_10_3 (.ZN (n_10_3), .A (n_7_6), .B (n_9_1), .C1 (n_5_3), .C2 (n_1_8) );
AOI211_X1 g_9_5 (.ZN (n_9_5), .A (n_8_4), .B (n_8_3), .C1 (n_7_2), .C2 (n_2_6) );
AOI211_X1 g_7_4 (.ZN (n_7_4), .A (n_10_3), .B (n_6_4), .C1 (n_9_1), .C2 (n_4_5) );
AOI211_X1 g_9_3 (.ZN (n_9_3), .A (n_9_5), .B (n_7_6), .C1 (n_8_3), .C2 (n_5_3) );
AOI211_X1 g_11_2 (.ZN (n_11_2), .A (n_7_4), .B (n_8_4), .C1 (n_6_4), .C2 (n_7_2) );
AOI211_X1 g_13_1 (.ZN (n_13_1), .A (n_9_3), .B (n_10_3), .C1 (n_7_6), .C2 (n_9_1) );
AOI211_X1 g_14_3 (.ZN (n_14_3), .A (n_11_2), .B (n_9_5), .C1 (n_8_4), .C2 (n_8_3) );
AOI211_X1 g_12_4 (.ZN (n_12_4), .A (n_13_1), .B (n_7_4), .C1 (n_10_3), .C2 (n_6_4) );
AOI211_X1 g_10_5 (.ZN (n_10_5), .A (n_14_3), .B (n_9_3), .C1 (n_9_5), .C2 (n_7_6) );
AOI211_X1 g_11_3 (.ZN (n_11_3), .A (n_12_4), .B (n_11_2), .C1 (n_7_4), .C2 (n_8_4) );
AOI211_X1 g_12_1 (.ZN (n_12_1), .A (n_10_5), .B (n_13_1), .C1 (n_9_3), .C2 (n_10_3) );
AOI211_X1 g_10_2 (.ZN (n_10_2), .A (n_11_3), .B (n_14_3), .C1 (n_11_2), .C2 (n_9_5) );
AOI211_X1 g_9_4 (.ZN (n_9_4), .A (n_12_1), .B (n_12_4), .C1 (n_13_1), .C2 (n_7_4) );
AOI211_X1 g_8_6 (.ZN (n_8_6), .A (n_10_2), .B (n_10_5), .C1 (n_14_3), .C2 (n_9_3) );
AOI211_X1 g_6_5 (.ZN (n_6_5), .A (n_9_4), .B (n_11_3), .C1 (n_12_4), .C2 (n_11_2) );
AOI211_X1 g_5_7 (.ZN (n_5_7), .A (n_8_6), .B (n_12_1), .C1 (n_10_5), .C2 (n_13_1) );
AOI211_X1 g_3_8 (.ZN (n_3_8), .A (n_6_5), .B (n_10_2), .C1 (n_11_3), .C2 (n_14_3) );
AOI211_X1 g_2_10 (.ZN (n_2_10), .A (n_5_7), .B (n_9_4), .C1 (n_12_1), .C2 (n_12_4) );
AOI211_X1 g_1_12 (.ZN (n_1_12), .A (n_3_8), .B (n_8_6), .C1 (n_10_2), .C2 (n_10_5) );
AOI211_X1 g_3_13 (.ZN (n_3_13), .A (n_2_10), .B (n_6_5), .C1 (n_9_4), .C2 (n_11_3) );
AOI211_X1 g_4_11 (.ZN (n_4_11), .A (n_1_12), .B (n_5_7), .C1 (n_8_6), .C2 (n_12_1) );
AOI211_X1 g_3_9 (.ZN (n_3_9), .A (n_3_13), .B (n_3_8), .C1 (n_6_5), .C2 (n_10_2) );
AOI211_X1 g_4_7 (.ZN (n_4_7), .A (n_4_11), .B (n_2_10), .C1 (n_5_7), .C2 (n_9_4) );
AOI211_X1 g_5_9 (.ZN (n_5_9), .A (n_3_9), .B (n_1_12), .C1 (n_3_8), .C2 (n_8_6) );
AOI211_X1 g_7_8 (.ZN (n_7_8), .A (n_4_7), .B (n_3_13), .C1 (n_2_10), .C2 (n_6_5) );
AOI211_X1 g_6_6 (.ZN (n_6_6), .A (n_5_9), .B (n_4_11), .C1 (n_1_12), .C2 (n_5_7) );
AOI211_X1 g_8_5 (.ZN (n_8_5), .A (n_7_8), .B (n_3_9), .C1 (n_3_13), .C2 (n_3_8) );
AOI211_X1 g_10_4 (.ZN (n_10_4), .A (n_6_6), .B (n_4_7), .C1 (n_4_11), .C2 (n_2_10) );
AOI211_X1 g_12_3 (.ZN (n_12_3), .A (n_8_5), .B (n_5_9), .C1 (n_3_9), .C2 (n_1_12) );
AOI211_X1 g_14_2 (.ZN (n_14_2), .A (n_10_4), .B (n_7_8), .C1 (n_4_7), .C2 (n_3_13) );
AOI211_X1 g_16_1 (.ZN (n_16_1), .A (n_12_3), .B (n_6_6), .C1 (n_5_9), .C2 (n_4_11) );
AOI211_X1 g_15_3 (.ZN (n_15_3), .A (n_14_2), .B (n_8_5), .C1 (n_7_8), .C2 (n_3_9) );
AOI211_X1 g_13_4 (.ZN (n_13_4), .A (n_16_1), .B (n_10_4), .C1 (n_6_6), .C2 (n_4_7) );
AOI211_X1 g_11_5 (.ZN (n_11_5), .A (n_15_3), .B (n_12_3), .C1 (n_8_5), .C2 (n_5_9) );
AOI211_X1 g_9_6 (.ZN (n_9_6), .A (n_13_4), .B (n_14_2), .C1 (n_10_4), .C2 (n_7_8) );
AOI211_X1 g_7_7 (.ZN (n_7_7), .A (n_11_5), .B (n_16_1), .C1 (n_12_3), .C2 (n_6_6) );
AOI211_X1 g_5_8 (.ZN (n_5_8), .A (n_9_6), .B (n_15_3), .C1 (n_14_2), .C2 (n_8_5) );
AOI211_X1 g_4_10 (.ZN (n_4_10), .A (n_7_7), .B (n_13_4), .C1 (n_16_1), .C2 (n_10_4) );
AOI211_X1 g_6_9 (.ZN (n_6_9), .A (n_5_8), .B (n_11_5), .C1 (n_15_3), .C2 (n_12_3) );
AOI211_X1 g_8_8 (.ZN (n_8_8), .A (n_4_10), .B (n_9_6), .C1 (n_13_4), .C2 (n_14_2) );
AOI211_X1 g_10_7 (.ZN (n_10_7), .A (n_6_9), .B (n_7_7), .C1 (n_11_5), .C2 (n_16_1) );
AOI211_X1 g_12_6 (.ZN (n_12_6), .A (n_8_8), .B (n_5_8), .C1 (n_9_6), .C2 (n_15_3) );
AOI211_X1 g_11_4 (.ZN (n_11_4), .A (n_10_7), .B (n_4_10), .C1 (n_7_7), .C2 (n_13_4) );
AOI211_X1 g_13_3 (.ZN (n_13_3), .A (n_12_6), .B (n_6_9), .C1 (n_5_8), .C2 (n_11_5) );
AOI211_X1 g_15_2 (.ZN (n_15_2), .A (n_11_4), .B (n_8_8), .C1 (n_4_10), .C2 (n_9_6) );
AOI211_X1 g_17_1 (.ZN (n_17_1), .A (n_13_3), .B (n_10_7), .C1 (n_6_9), .C2 (n_7_7) );
AOI211_X1 g_18_3 (.ZN (n_18_3), .A (n_15_2), .B (n_12_6), .C1 (n_8_8), .C2 (n_5_8) );
AOI211_X1 g_16_4 (.ZN (n_16_4), .A (n_17_1), .B (n_11_4), .C1 (n_10_7), .C2 (n_4_10) );
AOI211_X1 g_14_5 (.ZN (n_14_5), .A (n_18_3), .B (n_13_3), .C1 (n_12_6), .C2 (n_6_9) );
AOI211_X1 g_13_7 (.ZN (n_13_7), .A (n_16_4), .B (n_15_2), .C1 (n_11_4), .C2 (n_8_8) );
AOI211_X1 g_12_5 (.ZN (n_12_5), .A (n_14_5), .B (n_17_1), .C1 (n_13_3), .C2 (n_10_7) );
AOI211_X1 g_14_4 (.ZN (n_14_4), .A (n_13_7), .B (n_18_3), .C1 (n_15_2), .C2 (n_12_6) );
AOI211_X1 g_16_3 (.ZN (n_16_3), .A (n_12_5), .B (n_16_4), .C1 (n_17_1), .C2 (n_11_4) );
AOI211_X1 g_18_2 (.ZN (n_18_2), .A (n_14_4), .B (n_14_5), .C1 (n_18_3), .C2 (n_13_3) );
AOI211_X1 g_20_1 (.ZN (n_20_1), .A (n_16_3), .B (n_13_7), .C1 (n_16_4), .C2 (n_15_2) );
AOI211_X1 g_19_3 (.ZN (n_19_3), .A (n_18_2), .B (n_12_5), .C1 (n_14_5), .C2 (n_17_1) );
AOI211_X1 g_17_4 (.ZN (n_17_4), .A (n_20_1), .B (n_14_4), .C1 (n_13_7), .C2 (n_18_3) );
AOI211_X1 g_15_5 (.ZN (n_15_5), .A (n_19_3), .B (n_16_3), .C1 (n_12_5), .C2 (n_16_4) );
AOI211_X1 g_13_6 (.ZN (n_13_6), .A (n_17_4), .B (n_18_2), .C1 (n_14_4), .C2 (n_14_5) );
AOI211_X1 g_11_7 (.ZN (n_11_7), .A (n_15_5), .B (n_20_1), .C1 (n_16_3), .C2 (n_13_7) );
AOI211_X1 g_9_8 (.ZN (n_9_8), .A (n_13_6), .B (n_19_3), .C1 (n_18_2), .C2 (n_12_5) );
AOI211_X1 g_10_6 (.ZN (n_10_6), .A (n_11_7), .B (n_17_4), .C1 (n_20_1), .C2 (n_14_4) );
AOI211_X1 g_8_7 (.ZN (n_8_7), .A (n_9_8), .B (n_15_5), .C1 (n_19_3), .C2 (n_16_3) );
AOI211_X1 g_6_8 (.ZN (n_6_8), .A (n_10_6), .B (n_13_6), .C1 (n_17_4), .C2 (n_18_2) );
AOI211_X1 g_4_9 (.ZN (n_4_9), .A (n_8_7), .B (n_11_7), .C1 (n_15_5), .C2 (n_20_1) );
AOI211_X1 g_3_11 (.ZN (n_3_11), .A (n_6_8), .B (n_9_8), .C1 (n_13_6), .C2 (n_19_3) );
AOI211_X1 g_5_10 (.ZN (n_5_10), .A (n_4_9), .B (n_10_6), .C1 (n_11_7), .C2 (n_17_4) );
AOI211_X1 g_7_9 (.ZN (n_7_9), .A (n_3_11), .B (n_8_7), .C1 (n_9_8), .C2 (n_15_5) );
AOI211_X1 g_6_11 (.ZN (n_6_11), .A (n_5_10), .B (n_6_8), .C1 (n_10_6), .C2 (n_13_6) );
AOI211_X1 g_8_10 (.ZN (n_8_10), .A (n_7_9), .B (n_4_9), .C1 (n_8_7), .C2 (n_11_7) );
AOI211_X1 g_10_9 (.ZN (n_10_9), .A (n_6_11), .B (n_3_11), .C1 (n_6_8), .C2 (n_9_8) );
AOI211_X1 g_9_7 (.ZN (n_9_7), .A (n_8_10), .B (n_5_10), .C1 (n_4_9), .C2 (n_10_6) );
AOI211_X1 g_11_6 (.ZN (n_11_6), .A (n_10_9), .B (n_7_9), .C1 (n_3_11), .C2 (n_8_7) );
AOI211_X1 g_13_5 (.ZN (n_13_5), .A (n_9_7), .B (n_6_11), .C1 (n_5_10), .C2 (n_6_8) );
AOI211_X1 g_15_4 (.ZN (n_15_4), .A (n_11_6), .B (n_8_10), .C1 (n_7_9), .C2 (n_4_9) );
AOI211_X1 g_17_3 (.ZN (n_17_3), .A (n_13_5), .B (n_10_9), .C1 (n_6_11), .C2 (n_3_11) );
AOI211_X1 g_19_2 (.ZN (n_19_2), .A (n_15_4), .B (n_9_7), .C1 (n_8_10), .C2 (n_5_10) );
AOI211_X1 g_21_1 (.ZN (n_21_1), .A (n_17_3), .B (n_11_6), .C1 (n_10_9), .C2 (n_7_9) );
AOI211_X1 g_22_3 (.ZN (n_22_3), .A (n_19_2), .B (n_13_5), .C1 (n_9_7), .C2 (n_6_11) );
AOI211_X1 g_20_4 (.ZN (n_20_4), .A (n_21_1), .B (n_15_4), .C1 (n_11_6), .C2 (n_8_10) );
AOI211_X1 g_18_5 (.ZN (n_18_5), .A (n_22_3), .B (n_17_3), .C1 (n_13_5), .C2 (n_10_9) );
AOI211_X1 g_16_6 (.ZN (n_16_6), .A (n_20_4), .B (n_19_2), .C1 (n_15_4), .C2 (n_9_7) );
AOI211_X1 g_14_7 (.ZN (n_14_7), .A (n_18_5), .B (n_21_1), .C1 (n_17_3), .C2 (n_11_6) );
AOI211_X1 g_12_8 (.ZN (n_12_8), .A (n_16_6), .B (n_22_3), .C1 (n_19_2), .C2 (n_13_5) );
AOI211_X1 g_14_9 (.ZN (n_14_9), .A (n_14_7), .B (n_20_4), .C1 (n_21_1), .C2 (n_15_4) );
AOI211_X1 g_15_7 (.ZN (n_15_7), .A (n_12_8), .B (n_18_5), .C1 (n_22_3), .C2 (n_17_3) );
AOI211_X1 g_16_5 (.ZN (n_16_5), .A (n_14_9), .B (n_16_6), .C1 (n_20_4), .C2 (n_19_2) );
AOI211_X1 g_18_4 (.ZN (n_18_4), .A (n_15_7), .B (n_14_7), .C1 (n_18_5), .C2 (n_21_1) );
AOI211_X1 g_20_3 (.ZN (n_20_3), .A (n_16_5), .B (n_12_8), .C1 (n_16_6), .C2 (n_22_3) );
AOI211_X1 g_22_2 (.ZN (n_22_2), .A (n_18_4), .B (n_14_9), .C1 (n_14_7), .C2 (n_20_4) );
AOI211_X1 g_24_1 (.ZN (n_24_1), .A (n_20_3), .B (n_15_7), .C1 (n_12_8), .C2 (n_18_5) );
AOI211_X1 g_23_3 (.ZN (n_23_3), .A (n_22_2), .B (n_16_5), .C1 (n_14_9), .C2 (n_16_6) );
AOI211_X1 g_21_4 (.ZN (n_21_4), .A (n_24_1), .B (n_18_4), .C1 (n_15_7), .C2 (n_14_7) );
AOI211_X1 g_19_5 (.ZN (n_19_5), .A (n_23_3), .B (n_20_3), .C1 (n_16_5), .C2 (n_12_8) );
AOI211_X1 g_17_6 (.ZN (n_17_6), .A (n_21_4), .B (n_22_2), .C1 (n_18_4), .C2 (n_14_9) );
AOI211_X1 g_16_8 (.ZN (n_16_8), .A (n_19_5), .B (n_24_1), .C1 (n_20_3), .C2 (n_15_7) );
AOI211_X1 g_15_6 (.ZN (n_15_6), .A (n_17_6), .B (n_23_3), .C1 (n_22_2), .C2 (n_16_5) );
AOI211_X1 g_17_5 (.ZN (n_17_5), .A (n_16_8), .B (n_21_4), .C1 (n_24_1), .C2 (n_18_4) );
AOI211_X1 g_19_4 (.ZN (n_19_4), .A (n_15_6), .B (n_19_5), .C1 (n_23_3), .C2 (n_20_3) );
AOI211_X1 g_21_3 (.ZN (n_21_3), .A (n_17_5), .B (n_17_6), .C1 (n_21_4), .C2 (n_22_2) );
AOI211_X1 g_23_2 (.ZN (n_23_2), .A (n_19_4), .B (n_16_8), .C1 (n_19_5), .C2 (n_24_1) );
AOI211_X1 g_25_1 (.ZN (n_25_1), .A (n_21_3), .B (n_15_6), .C1 (n_17_6), .C2 (n_23_3) );
AOI211_X1 g_26_3 (.ZN (n_26_3), .A (n_23_2), .B (n_17_5), .C1 (n_16_8), .C2 (n_21_4) );
AOI211_X1 g_24_4 (.ZN (n_24_4), .A (n_25_1), .B (n_19_4), .C1 (n_15_6), .C2 (n_19_5) );
AOI211_X1 g_22_5 (.ZN (n_22_5), .A (n_26_3), .B (n_21_3), .C1 (n_17_5), .C2 (n_17_6) );
AOI211_X1 g_20_6 (.ZN (n_20_6), .A (n_24_4), .B (n_23_2), .C1 (n_19_4), .C2 (n_16_8) );
AOI211_X1 g_18_7 (.ZN (n_18_7), .A (n_22_5), .B (n_25_1), .C1 (n_21_3), .C2 (n_15_6) );
AOI211_X1 g_17_9 (.ZN (n_17_9), .A (n_20_6), .B (n_26_3), .C1 (n_23_2), .C2 (n_17_5) );
AOI211_X1 g_16_7 (.ZN (n_16_7), .A (n_18_7), .B (n_24_4), .C1 (n_25_1), .C2 (n_19_4) );
AOI211_X1 g_14_6 (.ZN (n_14_6), .A (n_17_9), .B (n_22_5), .C1 (n_26_3), .C2 (n_21_3) );
AOI211_X1 g_12_7 (.ZN (n_12_7), .A (n_16_7), .B (n_20_6), .C1 (n_24_4), .C2 (n_23_2) );
AOI211_X1 g_10_8 (.ZN (n_10_8), .A (n_14_6), .B (n_18_7), .C1 (n_22_5), .C2 (n_25_1) );
AOI211_X1 g_8_9 (.ZN (n_8_9), .A (n_12_7), .B (n_17_9), .C1 (n_20_6), .C2 (n_26_3) );
AOI211_X1 g_6_10 (.ZN (n_6_10), .A (n_10_8), .B (n_16_7), .C1 (n_18_7), .C2 (n_24_4) );
AOI211_X1 g_5_12 (.ZN (n_5_12), .A (n_8_9), .B (n_14_6), .C1 (n_17_9), .C2 (n_22_5) );
AOI211_X1 g_7_11 (.ZN (n_7_11), .A (n_6_10), .B (n_12_7), .C1 (n_16_7), .C2 (n_20_6) );
AOI211_X1 g_9_10 (.ZN (n_9_10), .A (n_5_12), .B (n_10_8), .C1 (n_14_6), .C2 (n_18_7) );
AOI211_X1 g_11_9 (.ZN (n_11_9), .A (n_7_11), .B (n_8_9), .C1 (n_12_7), .C2 (n_17_9) );
AOI211_X1 g_13_8 (.ZN (n_13_8), .A (n_9_10), .B (n_6_10), .C1 (n_10_8), .C2 (n_16_7) );
AOI211_X1 g_12_10 (.ZN (n_12_10), .A (n_11_9), .B (n_5_12), .C1 (n_8_9), .C2 (n_14_6) );
AOI211_X1 g_11_8 (.ZN (n_11_8), .A (n_13_8), .B (n_7_11), .C1 (n_6_10), .C2 (n_12_7) );
AOI211_X1 g_9_9 (.ZN (n_9_9), .A (n_12_10), .B (n_9_10), .C1 (n_5_12), .C2 (n_10_8) );
AOI211_X1 g_7_10 (.ZN (n_7_10), .A (n_11_8), .B (n_11_9), .C1 (n_7_11), .C2 (n_8_9) );
AOI211_X1 g_5_11 (.ZN (n_5_11), .A (n_9_9), .B (n_13_8), .C1 (n_9_10), .C2 (n_6_10) );
AOI211_X1 g_3_12 (.ZN (n_3_12), .A (n_7_10), .B (n_12_10), .C1 (n_11_9), .C2 (n_5_12) );
AOI211_X1 g_2_14 (.ZN (n_2_14), .A (n_5_11), .B (n_11_8), .C1 (n_13_8), .C2 (n_7_11) );
AOI211_X1 g_1_16 (.ZN (n_1_16), .A (n_3_12), .B (n_9_9), .C1 (n_12_10), .C2 (n_9_10) );
AOI211_X1 g_3_17 (.ZN (n_3_17), .A (n_2_14), .B (n_7_10), .C1 (n_11_8), .C2 (n_11_9) );
AOI211_X1 g_4_15 (.ZN (n_4_15), .A (n_1_16), .B (n_5_11), .C1 (n_9_9), .C2 (n_13_8) );
AOI211_X1 g_5_13 (.ZN (n_5_13), .A (n_3_17), .B (n_3_12), .C1 (n_7_10), .C2 (n_12_10) );
AOI211_X1 g_7_12 (.ZN (n_7_12), .A (n_4_15), .B (n_2_14), .C1 (n_5_11), .C2 (n_11_8) );
AOI211_X1 g_9_11 (.ZN (n_9_11), .A (n_5_13), .B (n_1_16), .C1 (n_3_12), .C2 (n_9_9) );
AOI211_X1 g_11_10 (.ZN (n_11_10), .A (n_7_12), .B (n_3_17), .C1 (n_2_14), .C2 (n_7_10) );
AOI211_X1 g_13_9 (.ZN (n_13_9), .A (n_9_11), .B (n_4_15), .C1 (n_1_16), .C2 (n_5_11) );
AOI211_X1 g_15_8 (.ZN (n_15_8), .A (n_11_10), .B (n_5_13), .C1 (n_3_17), .C2 (n_3_12) );
AOI211_X1 g_17_7 (.ZN (n_17_7), .A (n_13_9), .B (n_7_12), .C1 (n_4_15), .C2 (n_2_14) );
AOI211_X1 g_19_6 (.ZN (n_19_6), .A (n_15_8), .B (n_9_11), .C1 (n_5_13), .C2 (n_1_16) );
AOI211_X1 g_21_5 (.ZN (n_21_5), .A (n_17_7), .B (n_11_10), .C1 (n_7_12), .C2 (n_3_17) );
AOI211_X1 g_23_4 (.ZN (n_23_4), .A (n_19_6), .B (n_13_9), .C1 (n_9_11), .C2 (n_4_15) );
AOI211_X1 g_25_3 (.ZN (n_25_3), .A (n_21_5), .B (n_15_8), .C1 (n_11_10), .C2 (n_5_13) );
AOI211_X1 g_27_2 (.ZN (n_27_2), .A (n_23_4), .B (n_17_7), .C1 (n_13_9), .C2 (n_7_12) );
AOI211_X1 g_29_1 (.ZN (n_29_1), .A (n_25_3), .B (n_19_6), .C1 (n_15_8), .C2 (n_9_11) );
AOI211_X1 g_30_3 (.ZN (n_30_3), .A (n_27_2), .B (n_21_5), .C1 (n_17_7), .C2 (n_11_10) );
AOI211_X1 g_28_4 (.ZN (n_28_4), .A (n_29_1), .B (n_23_4), .C1 (n_19_6), .C2 (n_13_9) );
AOI211_X1 g_26_5 (.ZN (n_26_5), .A (n_30_3), .B (n_25_3), .C1 (n_21_5), .C2 (n_15_8) );
AOI211_X1 g_27_3 (.ZN (n_27_3), .A (n_28_4), .B (n_27_2), .C1 (n_23_4), .C2 (n_17_7) );
AOI211_X1 g_28_1 (.ZN (n_28_1), .A (n_26_5), .B (n_29_1), .C1 (n_25_3), .C2 (n_19_6) );
AOI211_X1 g_26_2 (.ZN (n_26_2), .A (n_27_3), .B (n_30_3), .C1 (n_27_2), .C2 (n_21_5) );
AOI211_X1 g_24_3 (.ZN (n_24_3), .A (n_28_1), .B (n_28_4), .C1 (n_29_1), .C2 (n_23_4) );
AOI211_X1 g_22_4 (.ZN (n_22_4), .A (n_26_2), .B (n_26_5), .C1 (n_30_3), .C2 (n_25_3) );
AOI211_X1 g_20_5 (.ZN (n_20_5), .A (n_24_3), .B (n_27_3), .C1 (n_28_4), .C2 (n_27_2) );
AOI211_X1 g_18_6 (.ZN (n_18_6), .A (n_22_4), .B (n_28_1), .C1 (n_26_5), .C2 (n_29_1) );
AOI211_X1 g_19_8 (.ZN (n_19_8), .A (n_20_5), .B (n_26_2), .C1 (n_27_3), .C2 (n_30_3) );
AOI211_X1 g_21_7 (.ZN (n_21_7), .A (n_18_6), .B (n_24_3), .C1 (n_28_1), .C2 (n_28_4) );
AOI211_X1 g_23_6 (.ZN (n_23_6), .A (n_19_8), .B (n_22_4), .C1 (n_26_2), .C2 (n_26_5) );
AOI211_X1 g_25_5 (.ZN (n_25_5), .A (n_21_7), .B (n_20_5), .C1 (n_24_3), .C2 (n_27_3) );
AOI211_X1 g_27_4 (.ZN (n_27_4), .A (n_23_6), .B (n_18_6), .C1 (n_22_4), .C2 (n_28_1) );
AOI211_X1 g_29_3 (.ZN (n_29_3), .A (n_25_5), .B (n_19_8), .C1 (n_20_5), .C2 (n_26_2) );
AOI211_X1 g_31_2 (.ZN (n_31_2), .A (n_27_4), .B (n_21_7), .C1 (n_18_6), .C2 (n_24_3) );
AOI211_X1 g_33_1 (.ZN (n_33_1), .A (n_29_3), .B (n_23_6), .C1 (n_19_8), .C2 (n_22_4) );
AOI211_X1 g_34_3 (.ZN (n_34_3), .A (n_31_2), .B (n_25_5), .C1 (n_21_7), .C2 (n_20_5) );
AOI211_X1 g_32_4 (.ZN (n_32_4), .A (n_33_1), .B (n_27_4), .C1 (n_23_6), .C2 (n_18_6) );
AOI211_X1 g_30_5 (.ZN (n_30_5), .A (n_34_3), .B (n_29_3), .C1 (n_25_5), .C2 (n_19_8) );
AOI211_X1 g_31_3 (.ZN (n_31_3), .A (n_32_4), .B (n_31_2), .C1 (n_27_4), .C2 (n_21_7) );
AOI211_X1 g_32_1 (.ZN (n_32_1), .A (n_30_5), .B (n_33_1), .C1 (n_29_3), .C2 (n_23_6) );
AOI211_X1 g_30_2 (.ZN (n_30_2), .A (n_31_3), .B (n_34_3), .C1 (n_31_2), .C2 (n_25_5) );
AOI211_X1 g_28_3 (.ZN (n_28_3), .A (n_32_1), .B (n_32_4), .C1 (n_33_1), .C2 (n_27_4) );
AOI211_X1 g_26_4 (.ZN (n_26_4), .A (n_30_2), .B (n_30_5), .C1 (n_34_3), .C2 (n_29_3) );
AOI211_X1 g_24_5 (.ZN (n_24_5), .A (n_28_3), .B (n_31_3), .C1 (n_32_4), .C2 (n_31_2) );
AOI211_X1 g_22_6 (.ZN (n_22_6), .A (n_26_4), .B (n_32_1), .C1 (n_30_5), .C2 (n_33_1) );
AOI211_X1 g_20_7 (.ZN (n_20_7), .A (n_24_5), .B (n_30_2), .C1 (n_31_3), .C2 (n_34_3) );
AOI211_X1 g_18_8 (.ZN (n_18_8), .A (n_22_6), .B (n_28_3), .C1 (n_32_1), .C2 (n_32_4) );
AOI211_X1 g_16_9 (.ZN (n_16_9), .A (n_20_7), .B (n_26_4), .C1 (n_30_2), .C2 (n_30_5) );
AOI211_X1 g_14_8 (.ZN (n_14_8), .A (n_18_8), .B (n_24_5), .C1 (n_28_3), .C2 (n_31_3) );
AOI211_X1 g_12_9 (.ZN (n_12_9), .A (n_16_9), .B (n_22_6), .C1 (n_26_4), .C2 (n_32_1) );
AOI211_X1 g_10_10 (.ZN (n_10_10), .A (n_14_8), .B (n_20_7), .C1 (n_24_5), .C2 (n_30_2) );
AOI211_X1 g_8_11 (.ZN (n_8_11), .A (n_12_9), .B (n_18_8), .C1 (n_22_6), .C2 (n_28_3) );
AOI211_X1 g_6_12 (.ZN (n_6_12), .A (n_10_10), .B (n_16_9), .C1 (n_20_7), .C2 (n_26_4) );
AOI211_X1 g_4_13 (.ZN (n_4_13), .A (n_8_11), .B (n_14_8), .C1 (n_18_8), .C2 (n_24_5) );
AOI211_X1 g_6_14 (.ZN (n_6_14), .A (n_6_12), .B (n_12_9), .C1 (n_16_9), .C2 (n_22_6) );
AOI211_X1 g_8_13 (.ZN (n_8_13), .A (n_4_13), .B (n_10_10), .C1 (n_14_8), .C2 (n_20_7) );
AOI211_X1 g_10_12 (.ZN (n_10_12), .A (n_6_14), .B (n_8_11), .C1 (n_12_9), .C2 (n_18_8) );
AOI211_X1 g_12_11 (.ZN (n_12_11), .A (n_8_13), .B (n_6_12), .C1 (n_10_10), .C2 (n_16_9) );
AOI211_X1 g_14_10 (.ZN (n_14_10), .A (n_10_12), .B (n_4_13), .C1 (n_8_11), .C2 (n_14_8) );
AOI211_X1 g_13_12 (.ZN (n_13_12), .A (n_12_11), .B (n_6_14), .C1 (n_6_12), .C2 (n_12_9) );
AOI211_X1 g_11_11 (.ZN (n_11_11), .A (n_14_10), .B (n_8_13), .C1 (n_4_13), .C2 (n_10_10) );
AOI211_X1 g_13_10 (.ZN (n_13_10), .A (n_13_12), .B (n_10_12), .C1 (n_6_14), .C2 (n_8_11) );
AOI211_X1 g_15_9 (.ZN (n_15_9), .A (n_11_11), .B (n_12_11), .C1 (n_8_13), .C2 (n_6_12) );
AOI211_X1 g_17_8 (.ZN (n_17_8), .A (n_13_10), .B (n_14_10), .C1 (n_10_12), .C2 (n_4_13) );
AOI211_X1 g_19_7 (.ZN (n_19_7), .A (n_15_9), .B (n_13_12), .C1 (n_12_11), .C2 (n_6_14) );
AOI211_X1 g_21_6 (.ZN (n_21_6), .A (n_17_8), .B (n_11_11), .C1 (n_14_10), .C2 (n_8_13) );
AOI211_X1 g_23_5 (.ZN (n_23_5), .A (n_19_7), .B (n_13_10), .C1 (n_13_12), .C2 (n_10_12) );
AOI211_X1 g_25_4 (.ZN (n_25_4), .A (n_21_6), .B (n_15_9), .C1 (n_11_11), .C2 (n_12_11) );
AOI211_X1 g_24_6 (.ZN (n_24_6), .A (n_23_5), .B (n_17_8), .C1 (n_13_10), .C2 (n_14_10) );
AOI211_X1 g_22_7 (.ZN (n_22_7), .A (n_25_4), .B (n_19_7), .C1 (n_15_9), .C2 (n_13_12) );
AOI211_X1 g_20_8 (.ZN (n_20_8), .A (n_24_6), .B (n_21_6), .C1 (n_17_8), .C2 (n_11_11) );
AOI211_X1 g_18_9 (.ZN (n_18_9), .A (n_22_7), .B (n_23_5), .C1 (n_19_7), .C2 (n_13_10) );
AOI211_X1 g_16_10 (.ZN (n_16_10), .A (n_20_8), .B (n_25_4), .C1 (n_21_6), .C2 (n_15_9) );
AOI211_X1 g_14_11 (.ZN (n_14_11), .A (n_18_9), .B (n_24_6), .C1 (n_23_5), .C2 (n_17_8) );
AOI211_X1 g_12_12 (.ZN (n_12_12), .A (n_16_10), .B (n_22_7), .C1 (n_25_4), .C2 (n_19_7) );
AOI211_X1 g_10_11 (.ZN (n_10_11), .A (n_14_11), .B (n_20_8), .C1 (n_24_6), .C2 (n_21_6) );
AOI211_X1 g_8_12 (.ZN (n_8_12), .A (n_12_12), .B (n_18_9), .C1 (n_22_7), .C2 (n_23_5) );
AOI211_X1 g_10_13 (.ZN (n_10_13), .A (n_10_11), .B (n_16_10), .C1 (n_20_8), .C2 (n_25_4) );
AOI211_X1 g_8_14 (.ZN (n_8_14), .A (n_8_12), .B (n_14_11), .C1 (n_18_9), .C2 (n_24_6) );
AOI211_X1 g_9_12 (.ZN (n_9_12), .A (n_10_13), .B (n_12_12), .C1 (n_16_10), .C2 (n_22_7) );
AOI211_X1 g_7_13 (.ZN (n_7_13), .A (n_8_14), .B (n_10_11), .C1 (n_14_11), .C2 (n_20_8) );
AOI211_X1 g_5_14 (.ZN (n_5_14), .A (n_9_12), .B (n_8_12), .C1 (n_12_12), .C2 (n_18_9) );
AOI211_X1 g_4_12 (.ZN (n_4_12), .A (n_7_13), .B (n_10_13), .C1 (n_10_11), .C2 (n_16_10) );
AOI211_X1 g_2_13 (.ZN (n_2_13), .A (n_5_14), .B (n_8_14), .C1 (n_8_12), .C2 (n_14_11) );
AOI211_X1 g_1_15 (.ZN (n_1_15), .A (n_4_12), .B (n_9_12), .C1 (n_10_13), .C2 (n_12_12) );
AOI211_X1 g_3_14 (.ZN (n_3_14), .A (n_2_13), .B (n_7_13), .C1 (n_8_14), .C2 (n_10_11) );
AOI211_X1 g_4_16 (.ZN (n_4_16), .A (n_1_15), .B (n_5_14), .C1 (n_9_12), .C2 (n_8_12) );
AOI211_X1 g_6_15 (.ZN (n_6_15), .A (n_3_14), .B (n_4_12), .C1 (n_7_13), .C2 (n_10_13) );
AOI211_X1 g_4_14 (.ZN (n_4_14), .A (n_4_16), .B (n_2_13), .C1 (n_5_14), .C2 (n_8_14) );
AOI211_X1 g_6_13 (.ZN (n_6_13), .A (n_6_15), .B (n_1_15), .C1 (n_4_12), .C2 (n_9_12) );
AOI211_X1 g_5_15 (.ZN (n_5_15), .A (n_4_14), .B (n_3_14), .C1 (n_2_13), .C2 (n_7_13) );
AOI211_X1 g_3_16 (.ZN (n_3_16), .A (n_6_13), .B (n_4_16), .C1 (n_1_15), .C2 (n_5_14) );
AOI211_X1 g_2_18 (.ZN (n_2_18), .A (n_5_15), .B (n_6_15), .C1 (n_3_14), .C2 (n_4_12) );
AOI211_X1 g_1_20 (.ZN (n_1_20), .A (n_3_16), .B (n_4_14), .C1 (n_4_16), .C2 (n_2_13) );
AOI211_X1 g_3_21 (.ZN (n_3_21), .A (n_2_18), .B (n_6_13), .C1 (n_6_15), .C2 (n_1_15) );
AOI211_X1 g_4_19 (.ZN (n_4_19), .A (n_1_20), .B (n_5_15), .C1 (n_4_14), .C2 (n_3_14) );
AOI211_X1 g_5_17 (.ZN (n_5_17), .A (n_3_21), .B (n_3_16), .C1 (n_6_13), .C2 (n_4_16) );
AOI211_X1 g_3_18 (.ZN (n_3_18), .A (n_4_19), .B (n_2_18), .C1 (n_5_15), .C2 (n_6_15) );
AOI211_X1 g_1_19 (.ZN (n_1_19), .A (n_5_17), .B (n_1_20), .C1 (n_3_16), .C2 (n_4_14) );
AOI211_X1 g_2_17 (.ZN (n_2_17), .A (n_3_18), .B (n_3_21), .C1 (n_2_18), .C2 (n_6_13) );
AOI211_X1 g_3_15 (.ZN (n_3_15), .A (n_1_19), .B (n_4_19), .C1 (n_1_20), .C2 (n_5_15) );
AOI211_X1 g_4_17 (.ZN (n_4_17), .A (n_2_17), .B (n_5_17), .C1 (n_3_21), .C2 (n_3_16) );
AOI211_X1 g_3_19 (.ZN (n_3_19), .A (n_3_15), .B (n_3_18), .C1 (n_4_19), .C2 (n_2_18) );
AOI211_X1 g_2_21 (.ZN (n_2_21), .A (n_4_17), .B (n_1_19), .C1 (n_5_17), .C2 (n_1_20) );
AOI211_X1 g_1_23 (.ZN (n_1_23), .A (n_3_19), .B (n_2_17), .C1 (n_3_18), .C2 (n_3_21) );
AOI211_X1 g_3_22 (.ZN (n_3_22), .A (n_2_21), .B (n_3_15), .C1 (n_1_19), .C2 (n_4_19) );
AOI211_X1 g_4_20 (.ZN (n_4_20), .A (n_1_23), .B (n_4_17), .C1 (n_2_17), .C2 (n_5_17) );
AOI211_X1 g_5_18 (.ZN (n_5_18), .A (n_3_22), .B (n_3_19), .C1 (n_3_15), .C2 (n_3_18) );
AOI211_X1 g_6_16 (.ZN (n_6_16), .A (n_4_20), .B (n_2_21), .C1 (n_4_17), .C2 (n_1_19) );
AOI211_X1 g_7_14 (.ZN (n_7_14), .A (n_5_18), .B (n_1_23), .C1 (n_3_19), .C2 (n_2_17) );
AOI211_X1 g_9_13 (.ZN (n_9_13), .A (n_6_16), .B (n_3_22), .C1 (n_2_21), .C2 (n_3_15) );
AOI211_X1 g_11_12 (.ZN (n_11_12), .A (n_7_14), .B (n_4_20), .C1 (n_1_23), .C2 (n_4_17) );
AOI211_X1 g_13_11 (.ZN (n_13_11), .A (n_9_13), .B (n_5_18), .C1 (n_3_22), .C2 (n_3_19) );
AOI211_X1 g_15_10 (.ZN (n_15_10), .A (n_11_12), .B (n_6_16), .C1 (n_4_20), .C2 (n_2_21) );
AOI211_X1 g_14_12 (.ZN (n_14_12), .A (n_13_11), .B (n_7_14), .C1 (n_5_18), .C2 (n_1_23) );
AOI211_X1 g_16_11 (.ZN (n_16_11), .A (n_15_10), .B (n_9_13), .C1 (n_6_16), .C2 (n_3_22) );
AOI211_X1 g_18_10 (.ZN (n_18_10), .A (n_14_12), .B (n_11_12), .C1 (n_7_14), .C2 (n_4_20) );
AOI211_X1 g_20_9 (.ZN (n_20_9), .A (n_16_11), .B (n_13_11), .C1 (n_9_13), .C2 (n_5_18) );
AOI211_X1 g_22_8 (.ZN (n_22_8), .A (n_18_10), .B (n_15_10), .C1 (n_11_12), .C2 (n_6_16) );
AOI211_X1 g_24_7 (.ZN (n_24_7), .A (n_20_9), .B (n_14_12), .C1 (n_13_11), .C2 (n_7_14) );
AOI211_X1 g_26_6 (.ZN (n_26_6), .A (n_22_8), .B (n_16_11), .C1 (n_15_10), .C2 (n_9_13) );
AOI211_X1 g_28_5 (.ZN (n_28_5), .A (n_24_7), .B (n_18_10), .C1 (n_14_12), .C2 (n_11_12) );
AOI211_X1 g_30_4 (.ZN (n_30_4), .A (n_26_6), .B (n_20_9), .C1 (n_16_11), .C2 (n_13_11) );
AOI211_X1 g_32_3 (.ZN (n_32_3), .A (n_28_5), .B (n_22_8), .C1 (n_18_10), .C2 (n_15_10) );
AOI211_X1 g_34_2 (.ZN (n_34_2), .A (n_30_4), .B (n_24_7), .C1 (n_20_9), .C2 (n_14_12) );
AOI211_X1 g_36_1 (.ZN (n_36_1), .A (n_32_3), .B (n_26_6), .C1 (n_22_8), .C2 (n_16_11) );
AOI211_X1 g_35_3 (.ZN (n_35_3), .A (n_34_2), .B (n_28_5), .C1 (n_24_7), .C2 (n_18_10) );
AOI211_X1 g_33_4 (.ZN (n_33_4), .A (n_36_1), .B (n_30_4), .C1 (n_26_6), .C2 (n_20_9) );
AOI211_X1 g_31_5 (.ZN (n_31_5), .A (n_35_3), .B (n_32_3), .C1 (n_28_5), .C2 (n_22_8) );
AOI211_X1 g_29_4 (.ZN (n_29_4), .A (n_33_4), .B (n_34_2), .C1 (n_30_4), .C2 (n_24_7) );
AOI211_X1 g_27_5 (.ZN (n_27_5), .A (n_31_5), .B (n_36_1), .C1 (n_32_3), .C2 (n_26_6) );
AOI211_X1 g_25_6 (.ZN (n_25_6), .A (n_29_4), .B (n_35_3), .C1 (n_34_2), .C2 (n_28_5) );
AOI211_X1 g_23_7 (.ZN (n_23_7), .A (n_27_5), .B (n_33_4), .C1 (n_36_1), .C2 (n_30_4) );
AOI211_X1 g_21_8 (.ZN (n_21_8), .A (n_25_6), .B (n_31_5), .C1 (n_35_3), .C2 (n_32_3) );
AOI211_X1 g_19_9 (.ZN (n_19_9), .A (n_23_7), .B (n_29_4), .C1 (n_33_4), .C2 (n_34_2) );
AOI211_X1 g_17_10 (.ZN (n_17_10), .A (n_21_8), .B (n_27_5), .C1 (n_31_5), .C2 (n_36_1) );
AOI211_X1 g_15_11 (.ZN (n_15_11), .A (n_19_9), .B (n_25_6), .C1 (n_29_4), .C2 (n_35_3) );
AOI211_X1 g_14_13 (.ZN (n_14_13), .A (n_17_10), .B (n_23_7), .C1 (n_27_5), .C2 (n_33_4) );
AOI211_X1 g_16_12 (.ZN (n_16_12), .A (n_15_11), .B (n_21_8), .C1 (n_25_6), .C2 (n_31_5) );
AOI211_X1 g_18_11 (.ZN (n_18_11), .A (n_14_13), .B (n_19_9), .C1 (n_23_7), .C2 (n_29_4) );
AOI211_X1 g_20_10 (.ZN (n_20_10), .A (n_16_12), .B (n_17_10), .C1 (n_21_8), .C2 (n_27_5) );
AOI211_X1 g_22_9 (.ZN (n_22_9), .A (n_18_11), .B (n_15_11), .C1 (n_19_9), .C2 (n_25_6) );
AOI211_X1 g_24_8 (.ZN (n_24_8), .A (n_20_10), .B (n_14_13), .C1 (n_17_10), .C2 (n_23_7) );
AOI211_X1 g_26_7 (.ZN (n_26_7), .A (n_22_9), .B (n_16_12), .C1 (n_15_11), .C2 (n_21_8) );
AOI211_X1 g_28_6 (.ZN (n_28_6), .A (n_24_8), .B (n_18_11), .C1 (n_14_13), .C2 (n_19_9) );
AOI211_X1 g_27_8 (.ZN (n_27_8), .A (n_26_7), .B (n_20_10), .C1 (n_16_12), .C2 (n_17_10) );
AOI211_X1 g_25_7 (.ZN (n_25_7), .A (n_28_6), .B (n_22_9), .C1 (n_18_11), .C2 (n_15_11) );
AOI211_X1 g_27_6 (.ZN (n_27_6), .A (n_27_8), .B (n_24_8), .C1 (n_20_10), .C2 (n_14_13) );
AOI211_X1 g_29_5 (.ZN (n_29_5), .A (n_25_7), .B (n_26_7), .C1 (n_22_9), .C2 (n_16_12) );
AOI211_X1 g_31_4 (.ZN (n_31_4), .A (n_27_6), .B (n_28_6), .C1 (n_24_8), .C2 (n_18_11) );
AOI211_X1 g_33_3 (.ZN (n_33_3), .A (n_29_5), .B (n_27_8), .C1 (n_26_7), .C2 (n_20_10) );
AOI211_X1 g_35_2 (.ZN (n_35_2), .A (n_31_4), .B (n_25_7), .C1 (n_28_6), .C2 (n_22_9) );
AOI211_X1 g_37_1 (.ZN (n_37_1), .A (n_33_3), .B (n_27_6), .C1 (n_27_8), .C2 (n_24_8) );
AOI211_X1 g_38_3 (.ZN (n_38_3), .A (n_35_2), .B (n_29_5), .C1 (n_25_7), .C2 (n_26_7) );
AOI211_X1 g_36_4 (.ZN (n_36_4), .A (n_37_1), .B (n_31_4), .C1 (n_27_6), .C2 (n_28_6) );
AOI211_X1 g_34_5 (.ZN (n_34_5), .A (n_38_3), .B (n_33_3), .C1 (n_29_5), .C2 (n_27_8) );
AOI211_X1 g_32_6 (.ZN (n_32_6), .A (n_36_4), .B (n_35_2), .C1 (n_31_4), .C2 (n_25_7) );
AOI211_X1 g_30_7 (.ZN (n_30_7), .A (n_34_5), .B (n_37_1), .C1 (n_33_3), .C2 (n_27_6) );
AOI211_X1 g_28_8 (.ZN (n_28_8), .A (n_32_6), .B (n_38_3), .C1 (n_35_2), .C2 (n_29_5) );
AOI211_X1 g_29_6 (.ZN (n_29_6), .A (n_30_7), .B (n_36_4), .C1 (n_37_1), .C2 (n_31_4) );
AOI211_X1 g_27_7 (.ZN (n_27_7), .A (n_28_8), .B (n_34_5), .C1 (n_38_3), .C2 (n_33_3) );
AOI211_X1 g_25_8 (.ZN (n_25_8), .A (n_29_6), .B (n_32_6), .C1 (n_36_4), .C2 (n_35_2) );
AOI211_X1 g_23_9 (.ZN (n_23_9), .A (n_27_7), .B (n_30_7), .C1 (n_34_5), .C2 (n_37_1) );
AOI211_X1 g_21_10 (.ZN (n_21_10), .A (n_25_8), .B (n_28_8), .C1 (n_32_6), .C2 (n_38_3) );
AOI211_X1 g_19_11 (.ZN (n_19_11), .A (n_23_9), .B (n_29_6), .C1 (n_30_7), .C2 (n_36_4) );
AOI211_X1 g_17_12 (.ZN (n_17_12), .A (n_21_10), .B (n_27_7), .C1 (n_28_8), .C2 (n_34_5) );
AOI211_X1 g_15_13 (.ZN (n_15_13), .A (n_19_11), .B (n_25_8), .C1 (n_29_6), .C2 (n_32_6) );
AOI211_X1 g_13_14 (.ZN (n_13_14), .A (n_17_12), .B (n_23_9), .C1 (n_27_7), .C2 (n_30_7) );
AOI211_X1 g_11_13 (.ZN (n_11_13), .A (n_15_13), .B (n_21_10), .C1 (n_25_8), .C2 (n_28_8) );
AOI211_X1 g_9_14 (.ZN (n_9_14), .A (n_13_14), .B (n_19_11), .C1 (n_23_9), .C2 (n_29_6) );
AOI211_X1 g_7_15 (.ZN (n_7_15), .A (n_11_13), .B (n_17_12), .C1 (n_21_10), .C2 (n_27_7) );
AOI211_X1 g_5_16 (.ZN (n_5_16), .A (n_9_14), .B (n_15_13), .C1 (n_19_11), .C2 (n_25_8) );
AOI211_X1 g_4_18 (.ZN (n_4_18), .A (n_7_15), .B (n_13_14), .C1 (n_17_12), .C2 (n_23_9) );
AOI211_X1 g_6_17 (.ZN (n_6_17), .A (n_5_16), .B (n_11_13), .C1 (n_15_13), .C2 (n_21_10) );
AOI211_X1 g_8_16 (.ZN (n_8_16), .A (n_4_18), .B (n_9_14), .C1 (n_13_14), .C2 (n_19_11) );
AOI211_X1 g_10_15 (.ZN (n_10_15), .A (n_6_17), .B (n_7_15), .C1 (n_11_13), .C2 (n_17_12) );
AOI211_X1 g_12_14 (.ZN (n_12_14), .A (n_8_16), .B (n_5_16), .C1 (n_9_14), .C2 (n_15_13) );
AOI211_X1 g_14_15 (.ZN (n_14_15), .A (n_10_15), .B (n_4_18), .C1 (n_7_15), .C2 (n_13_14) );
AOI211_X1 g_13_13 (.ZN (n_13_13), .A (n_12_14), .B (n_6_17), .C1 (n_5_16), .C2 (n_11_13) );
AOI211_X1 g_15_12 (.ZN (n_15_12), .A (n_14_15), .B (n_8_16), .C1 (n_4_18), .C2 (n_9_14) );
AOI211_X1 g_17_11 (.ZN (n_17_11), .A (n_13_13), .B (n_10_15), .C1 (n_6_17), .C2 (n_7_15) );
AOI211_X1 g_19_10 (.ZN (n_19_10), .A (n_15_12), .B (n_12_14), .C1 (n_8_16), .C2 (n_5_16) );
AOI211_X1 g_21_9 (.ZN (n_21_9), .A (n_17_11), .B (n_14_15), .C1 (n_10_15), .C2 (n_4_18) );
AOI211_X1 g_23_8 (.ZN (n_23_8), .A (n_19_10), .B (n_13_13), .C1 (n_12_14), .C2 (n_6_17) );
AOI211_X1 g_25_9 (.ZN (n_25_9), .A (n_21_9), .B (n_15_12), .C1 (n_14_15), .C2 (n_8_16) );
AOI211_X1 g_23_10 (.ZN (n_23_10), .A (n_23_8), .B (n_17_11), .C1 (n_13_13), .C2 (n_10_15) );
AOI211_X1 g_21_11 (.ZN (n_21_11), .A (n_25_9), .B (n_19_10), .C1 (n_15_12), .C2 (n_12_14) );
AOI211_X1 g_19_12 (.ZN (n_19_12), .A (n_23_10), .B (n_21_9), .C1 (n_17_11), .C2 (n_14_15) );
AOI211_X1 g_17_13 (.ZN (n_17_13), .A (n_21_11), .B (n_23_8), .C1 (n_19_10), .C2 (n_13_13) );
AOI211_X1 g_15_14 (.ZN (n_15_14), .A (n_19_12), .B (n_25_9), .C1 (n_21_9), .C2 (n_15_12) );
AOI211_X1 g_13_15 (.ZN (n_13_15), .A (n_17_13), .B (n_23_10), .C1 (n_23_8), .C2 (n_17_11) );
AOI211_X1 g_12_13 (.ZN (n_12_13), .A (n_15_14), .B (n_21_11), .C1 (n_25_9), .C2 (n_19_10) );
AOI211_X1 g_10_14 (.ZN (n_10_14), .A (n_13_15), .B (n_19_12), .C1 (n_23_10), .C2 (n_21_9) );
AOI211_X1 g_8_15 (.ZN (n_8_15), .A (n_12_13), .B (n_17_13), .C1 (n_21_11), .C2 (n_23_8) );
AOI211_X1 g_7_17 (.ZN (n_7_17), .A (n_10_14), .B (n_15_14), .C1 (n_19_12), .C2 (n_25_9) );
AOI211_X1 g_9_16 (.ZN (n_9_16), .A (n_8_15), .B (n_13_15), .C1 (n_17_13), .C2 (n_23_10) );
AOI211_X1 g_11_15 (.ZN (n_11_15), .A (n_7_17), .B (n_12_13), .C1 (n_15_14), .C2 (n_21_11) );
AOI211_X1 g_10_17 (.ZN (n_10_17), .A (n_9_16), .B (n_10_14), .C1 (n_13_15), .C2 (n_19_12) );
AOI211_X1 g_12_16 (.ZN (n_12_16), .A (n_11_15), .B (n_8_15), .C1 (n_12_13), .C2 (n_17_13) );
AOI211_X1 g_11_14 (.ZN (n_11_14), .A (n_10_17), .B (n_7_17), .C1 (n_10_14), .C2 (n_15_14) );
AOI211_X1 g_9_15 (.ZN (n_9_15), .A (n_12_16), .B (n_9_16), .C1 (n_8_15), .C2 (n_13_15) );
AOI211_X1 g_7_16 (.ZN (n_7_16), .A (n_11_14), .B (n_11_15), .C1 (n_7_17), .C2 (n_12_13) );
AOI211_X1 g_6_18 (.ZN (n_6_18), .A (n_9_15), .B (n_10_17), .C1 (n_9_16), .C2 (n_10_14) );
AOI211_X1 g_8_17 (.ZN (n_8_17), .A (n_7_16), .B (n_12_16), .C1 (n_11_15), .C2 (n_8_15) );
AOI211_X1 g_10_16 (.ZN (n_10_16), .A (n_6_18), .B (n_11_14), .C1 (n_10_17), .C2 (n_7_17) );
AOI211_X1 g_12_15 (.ZN (n_12_15), .A (n_8_17), .B (n_9_15), .C1 (n_12_16), .C2 (n_9_16) );
AOI211_X1 g_14_14 (.ZN (n_14_14), .A (n_10_16), .B (n_7_16), .C1 (n_11_14), .C2 (n_11_15) );
AOI211_X1 g_16_13 (.ZN (n_16_13), .A (n_12_15), .B (n_6_18), .C1 (n_9_15), .C2 (n_10_17) );
AOI211_X1 g_18_12 (.ZN (n_18_12), .A (n_14_14), .B (n_8_17), .C1 (n_7_16), .C2 (n_12_16) );
AOI211_X1 g_20_11 (.ZN (n_20_11), .A (n_16_13), .B (n_10_16), .C1 (n_6_18), .C2 (n_11_14) );
AOI211_X1 g_22_10 (.ZN (n_22_10), .A (n_18_12), .B (n_12_15), .C1 (n_8_17), .C2 (n_9_15) );
AOI211_X1 g_24_9 (.ZN (n_24_9), .A (n_20_11), .B (n_14_14), .C1 (n_10_16), .C2 (n_7_16) );
AOI211_X1 g_26_8 (.ZN (n_26_8), .A (n_22_10), .B (n_16_13), .C1 (n_12_15), .C2 (n_6_18) );
AOI211_X1 g_28_7 (.ZN (n_28_7), .A (n_24_9), .B (n_18_12), .C1 (n_14_14), .C2 (n_8_17) );
AOI211_X1 g_30_6 (.ZN (n_30_6), .A (n_26_8), .B (n_20_11), .C1 (n_16_13), .C2 (n_10_16) );
AOI211_X1 g_32_5 (.ZN (n_32_5), .A (n_28_7), .B (n_22_10), .C1 (n_18_12), .C2 (n_12_15) );
AOI211_X1 g_34_4 (.ZN (n_34_4), .A (n_30_6), .B (n_24_9), .C1 (n_20_11), .C2 (n_14_14) );
AOI211_X1 g_36_3 (.ZN (n_36_3), .A (n_32_5), .B (n_26_8), .C1 (n_22_10), .C2 (n_16_13) );
AOI211_X1 g_38_2 (.ZN (n_38_2), .A (n_34_4), .B (n_28_7), .C1 (n_24_9), .C2 (n_18_12) );
AOI211_X1 g_40_1 (.ZN (n_40_1), .A (n_36_3), .B (n_30_6), .C1 (n_26_8), .C2 (n_20_11) );
AOI211_X1 g_39_3 (.ZN (n_39_3), .A (n_38_2), .B (n_32_5), .C1 (n_28_7), .C2 (n_22_10) );
AOI211_X1 g_37_4 (.ZN (n_37_4), .A (n_40_1), .B (n_34_4), .C1 (n_30_6), .C2 (n_24_9) );
AOI211_X1 g_35_5 (.ZN (n_35_5), .A (n_39_3), .B (n_36_3), .C1 (n_32_5), .C2 (n_26_8) );
AOI211_X1 g_33_6 (.ZN (n_33_6), .A (n_37_4), .B (n_38_2), .C1 (n_34_4), .C2 (n_28_7) );
AOI211_X1 g_31_7 (.ZN (n_31_7), .A (n_35_5), .B (n_40_1), .C1 (n_36_3), .C2 (n_30_6) );
AOI211_X1 g_29_8 (.ZN (n_29_8), .A (n_33_6), .B (n_39_3), .C1 (n_38_2), .C2 (n_32_5) );
AOI211_X1 g_27_9 (.ZN (n_27_9), .A (n_31_7), .B (n_37_4), .C1 (n_40_1), .C2 (n_34_4) );
AOI211_X1 g_25_10 (.ZN (n_25_10), .A (n_29_8), .B (n_35_5), .C1 (n_39_3), .C2 (n_36_3) );
AOI211_X1 g_23_11 (.ZN (n_23_11), .A (n_27_9), .B (n_33_6), .C1 (n_37_4), .C2 (n_38_2) );
AOI211_X1 g_21_12 (.ZN (n_21_12), .A (n_25_10), .B (n_31_7), .C1 (n_35_5), .C2 (n_40_1) );
AOI211_X1 g_19_13 (.ZN (n_19_13), .A (n_23_11), .B (n_29_8), .C1 (n_33_6), .C2 (n_39_3) );
AOI211_X1 g_17_14 (.ZN (n_17_14), .A (n_21_12), .B (n_27_9), .C1 (n_31_7), .C2 (n_37_4) );
AOI211_X1 g_15_15 (.ZN (n_15_15), .A (n_19_13), .B (n_25_10), .C1 (n_29_8), .C2 (n_35_5) );
AOI211_X1 g_13_16 (.ZN (n_13_16), .A (n_17_14), .B (n_23_11), .C1 (n_27_9), .C2 (n_33_6) );
AOI211_X1 g_11_17 (.ZN (n_11_17), .A (n_15_15), .B (n_21_12), .C1 (n_25_10), .C2 (n_31_7) );
AOI211_X1 g_9_18 (.ZN (n_9_18), .A (n_13_16), .B (n_19_13), .C1 (n_23_11), .C2 (n_29_8) );
AOI211_X1 g_7_19 (.ZN (n_7_19), .A (n_11_17), .B (n_17_14), .C1 (n_21_12), .C2 (n_27_9) );
AOI211_X1 g_5_20 (.ZN (n_5_20), .A (n_9_18), .B (n_15_15), .C1 (n_19_13), .C2 (n_25_10) );
AOI211_X1 g_4_22 (.ZN (n_4_22), .A (n_7_19), .B (n_13_16), .C1 (n_17_14), .C2 (n_23_11) );
AOI211_X1 g_3_20 (.ZN (n_3_20), .A (n_5_20), .B (n_11_17), .C1 (n_15_15), .C2 (n_21_12) );
AOI211_X1 g_5_19 (.ZN (n_5_19), .A (n_4_22), .B (n_9_18), .C1 (n_13_16), .C2 (n_19_13) );
AOI211_X1 g_7_18 (.ZN (n_7_18), .A (n_3_20), .B (n_7_19), .C1 (n_11_17), .C2 (n_17_14) );
AOI211_X1 g_9_17 (.ZN (n_9_17), .A (n_5_19), .B (n_5_20), .C1 (n_9_18), .C2 (n_15_15) );
AOI211_X1 g_11_16 (.ZN (n_11_16), .A (n_7_18), .B (n_4_22), .C1 (n_7_19), .C2 (n_13_16) );
AOI211_X1 g_10_18 (.ZN (n_10_18), .A (n_9_17), .B (n_3_20), .C1 (n_5_20), .C2 (n_11_17) );
AOI211_X1 g_12_17 (.ZN (n_12_17), .A (n_11_16), .B (n_5_19), .C1 (n_4_22), .C2 (n_9_18) );
AOI211_X1 g_14_16 (.ZN (n_14_16), .A (n_10_18), .B (n_7_18), .C1 (n_3_20), .C2 (n_7_19) );
AOI211_X1 g_16_15 (.ZN (n_16_15), .A (n_12_17), .B (n_9_17), .C1 (n_5_19), .C2 (n_5_20) );
AOI211_X1 g_18_14 (.ZN (n_18_14), .A (n_14_16), .B (n_11_16), .C1 (n_7_18), .C2 (n_4_22) );
AOI211_X1 g_20_13 (.ZN (n_20_13), .A (n_16_15), .B (n_10_18), .C1 (n_9_17), .C2 (n_3_20) );
AOI211_X1 g_22_12 (.ZN (n_22_12), .A (n_18_14), .B (n_12_17), .C1 (n_11_16), .C2 (n_5_19) );
AOI211_X1 g_24_11 (.ZN (n_24_11), .A (n_20_13), .B (n_14_16), .C1 (n_10_18), .C2 (n_7_18) );
AOI211_X1 g_26_10 (.ZN (n_26_10), .A (n_22_12), .B (n_16_15), .C1 (n_12_17), .C2 (n_9_17) );
AOI211_X1 g_28_9 (.ZN (n_28_9), .A (n_24_11), .B (n_18_14), .C1 (n_14_16), .C2 (n_11_16) );
AOI211_X1 g_29_7 (.ZN (n_29_7), .A (n_26_10), .B (n_20_13), .C1 (n_16_15), .C2 (n_10_18) );
AOI211_X1 g_31_6 (.ZN (n_31_6), .A (n_28_9), .B (n_22_12), .C1 (n_18_14), .C2 (n_12_17) );
AOI211_X1 g_33_5 (.ZN (n_33_5), .A (n_29_7), .B (n_24_11), .C1 (n_20_13), .C2 (n_14_16) );
AOI211_X1 g_35_4 (.ZN (n_35_4), .A (n_31_6), .B (n_26_10), .C1 (n_22_12), .C2 (n_16_15) );
AOI211_X1 g_37_3 (.ZN (n_37_3), .A (n_33_5), .B (n_28_9), .C1 (n_24_11), .C2 (n_18_14) );
AOI211_X1 g_39_2 (.ZN (n_39_2), .A (n_35_4), .B (n_29_7), .C1 (n_26_10), .C2 (n_20_13) );
AOI211_X1 g_41_1 (.ZN (n_41_1), .A (n_37_3), .B (n_31_6), .C1 (n_28_9), .C2 (n_22_12) );
AOI211_X1 g_42_3 (.ZN (n_42_3), .A (n_39_2), .B (n_33_5), .C1 (n_29_7), .C2 (n_24_11) );
AOI211_X1 g_40_4 (.ZN (n_40_4), .A (n_41_1), .B (n_35_4), .C1 (n_31_6), .C2 (n_26_10) );
AOI211_X1 g_38_5 (.ZN (n_38_5), .A (n_42_3), .B (n_37_3), .C1 (n_33_5), .C2 (n_28_9) );
AOI211_X1 g_36_6 (.ZN (n_36_6), .A (n_40_4), .B (n_39_2), .C1 (n_35_4), .C2 (n_29_7) );
AOI211_X1 g_34_7 (.ZN (n_34_7), .A (n_38_5), .B (n_41_1), .C1 (n_37_3), .C2 (n_31_6) );
AOI211_X1 g_32_8 (.ZN (n_32_8), .A (n_36_6), .B (n_42_3), .C1 (n_39_2), .C2 (n_33_5) );
AOI211_X1 g_30_9 (.ZN (n_30_9), .A (n_34_7), .B (n_40_4), .C1 (n_41_1), .C2 (n_35_4) );
AOI211_X1 g_28_10 (.ZN (n_28_10), .A (n_32_8), .B (n_38_5), .C1 (n_42_3), .C2 (n_37_3) );
AOI211_X1 g_26_9 (.ZN (n_26_9), .A (n_30_9), .B (n_36_6), .C1 (n_40_4), .C2 (n_39_2) );
AOI211_X1 g_24_10 (.ZN (n_24_10), .A (n_28_10), .B (n_34_7), .C1 (n_38_5), .C2 (n_41_1) );
AOI211_X1 g_22_11 (.ZN (n_22_11), .A (n_26_9), .B (n_32_8), .C1 (n_36_6), .C2 (n_42_3) );
AOI211_X1 g_20_12 (.ZN (n_20_12), .A (n_24_10), .B (n_30_9), .C1 (n_34_7), .C2 (n_40_4) );
AOI211_X1 g_18_13 (.ZN (n_18_13), .A (n_22_11), .B (n_28_10), .C1 (n_32_8), .C2 (n_38_5) );
AOI211_X1 g_16_14 (.ZN (n_16_14), .A (n_20_12), .B (n_26_9), .C1 (n_30_9), .C2 (n_36_6) );
AOI211_X1 g_15_16 (.ZN (n_15_16), .A (n_18_13), .B (n_24_10), .C1 (n_28_10), .C2 (n_34_7) );
AOI211_X1 g_17_15 (.ZN (n_17_15), .A (n_16_14), .B (n_22_11), .C1 (n_26_9), .C2 (n_32_8) );
AOI211_X1 g_19_14 (.ZN (n_19_14), .A (n_15_16), .B (n_20_12), .C1 (n_24_10), .C2 (n_30_9) );
AOI211_X1 g_21_13 (.ZN (n_21_13), .A (n_17_15), .B (n_18_13), .C1 (n_22_11), .C2 (n_28_10) );
AOI211_X1 g_23_12 (.ZN (n_23_12), .A (n_19_14), .B (n_16_14), .C1 (n_20_12), .C2 (n_26_9) );
AOI211_X1 g_25_11 (.ZN (n_25_11), .A (n_21_13), .B (n_15_16), .C1 (n_18_13), .C2 (n_24_10) );
AOI211_X1 g_27_10 (.ZN (n_27_10), .A (n_23_12), .B (n_17_15), .C1 (n_16_14), .C2 (n_22_11) );
AOI211_X1 g_29_9 (.ZN (n_29_9), .A (n_25_11), .B (n_19_14), .C1 (n_15_16), .C2 (n_20_12) );
AOI211_X1 g_31_8 (.ZN (n_31_8), .A (n_27_10), .B (n_21_13), .C1 (n_17_15), .C2 (n_18_13) );
AOI211_X1 g_33_7 (.ZN (n_33_7), .A (n_29_9), .B (n_23_12), .C1 (n_19_14), .C2 (n_16_14) );
AOI211_X1 g_35_6 (.ZN (n_35_6), .A (n_31_8), .B (n_25_11), .C1 (n_21_13), .C2 (n_15_16) );
AOI211_X1 g_37_5 (.ZN (n_37_5), .A (n_33_7), .B (n_27_10), .C1 (n_23_12), .C2 (n_17_15) );
AOI211_X1 g_39_4 (.ZN (n_39_4), .A (n_35_6), .B (n_29_9), .C1 (n_25_11), .C2 (n_19_14) );
AOI211_X1 g_41_3 (.ZN (n_41_3), .A (n_37_5), .B (n_31_8), .C1 (n_27_10), .C2 (n_21_13) );
AOI211_X1 g_43_2 (.ZN (n_43_2), .A (n_39_4), .B (n_33_7), .C1 (n_29_9), .C2 (n_23_12) );
AOI211_X1 g_45_1 (.ZN (n_45_1), .A (n_41_3), .B (n_35_6), .C1 (n_31_8), .C2 (n_25_11) );
AOI211_X1 g_46_3 (.ZN (n_46_3), .A (n_43_2), .B (n_37_5), .C1 (n_33_7), .C2 (n_27_10) );
AOI211_X1 g_44_4 (.ZN (n_44_4), .A (n_45_1), .B (n_39_4), .C1 (n_35_6), .C2 (n_29_9) );
AOI211_X1 g_42_5 (.ZN (n_42_5), .A (n_46_3), .B (n_41_3), .C1 (n_37_5), .C2 (n_31_8) );
AOI211_X1 g_43_3 (.ZN (n_43_3), .A (n_44_4), .B (n_43_2), .C1 (n_39_4), .C2 (n_33_7) );
AOI211_X1 g_44_1 (.ZN (n_44_1), .A (n_42_5), .B (n_45_1), .C1 (n_41_3), .C2 (n_35_6) );
AOI211_X1 g_42_2 (.ZN (n_42_2), .A (n_43_3), .B (n_46_3), .C1 (n_43_2), .C2 (n_37_5) );
AOI211_X1 g_40_3 (.ZN (n_40_3), .A (n_44_1), .B (n_44_4), .C1 (n_45_1), .C2 (n_39_4) );
AOI211_X1 g_38_4 (.ZN (n_38_4), .A (n_42_2), .B (n_42_5), .C1 (n_46_3), .C2 (n_41_3) );
AOI211_X1 g_36_5 (.ZN (n_36_5), .A (n_40_3), .B (n_43_3), .C1 (n_44_4), .C2 (n_43_2) );
AOI211_X1 g_34_6 (.ZN (n_34_6), .A (n_38_4), .B (n_44_1), .C1 (n_42_5), .C2 (n_45_1) );
AOI211_X1 g_32_7 (.ZN (n_32_7), .A (n_36_5), .B (n_42_2), .C1 (n_43_3), .C2 (n_46_3) );
AOI211_X1 g_30_8 (.ZN (n_30_8), .A (n_34_6), .B (n_40_3), .C1 (n_44_1), .C2 (n_44_4) );
AOI211_X1 g_29_10 (.ZN (n_29_10), .A (n_32_7), .B (n_38_4), .C1 (n_42_2), .C2 (n_42_5) );
AOI211_X1 g_31_9 (.ZN (n_31_9), .A (n_30_8), .B (n_36_5), .C1 (n_40_3), .C2 (n_43_3) );
AOI211_X1 g_33_8 (.ZN (n_33_8), .A (n_29_10), .B (n_34_6), .C1 (n_38_4), .C2 (n_44_1) );
AOI211_X1 g_35_7 (.ZN (n_35_7), .A (n_31_9), .B (n_32_7), .C1 (n_36_5), .C2 (n_42_2) );
AOI211_X1 g_37_6 (.ZN (n_37_6), .A (n_33_8), .B (n_30_8), .C1 (n_34_6), .C2 (n_40_3) );
AOI211_X1 g_39_5 (.ZN (n_39_5), .A (n_35_7), .B (n_29_10), .C1 (n_32_7), .C2 (n_38_4) );
AOI211_X1 g_41_4 (.ZN (n_41_4), .A (n_37_6), .B (n_31_9), .C1 (n_30_8), .C2 (n_36_5) );
AOI211_X1 g_40_6 (.ZN (n_40_6), .A (n_39_5), .B (n_33_8), .C1 (n_29_10), .C2 (n_34_6) );
AOI211_X1 g_38_7 (.ZN (n_38_7), .A (n_41_4), .B (n_35_7), .C1 (n_31_9), .C2 (n_32_7) );
AOI211_X1 g_36_8 (.ZN (n_36_8), .A (n_40_6), .B (n_37_6), .C1 (n_33_8), .C2 (n_30_8) );
AOI211_X1 g_34_9 (.ZN (n_34_9), .A (n_38_7), .B (n_39_5), .C1 (n_35_7), .C2 (n_29_10) );
AOI211_X1 g_32_10 (.ZN (n_32_10), .A (n_36_8), .B (n_41_4), .C1 (n_37_6), .C2 (n_31_9) );
AOI211_X1 g_30_11 (.ZN (n_30_11), .A (n_34_9), .B (n_40_6), .C1 (n_39_5), .C2 (n_33_8) );
AOI211_X1 g_28_12 (.ZN (n_28_12), .A (n_32_10), .B (n_38_7), .C1 (n_41_4), .C2 (n_35_7) );
AOI211_X1 g_26_11 (.ZN (n_26_11), .A (n_30_11), .B (n_36_8), .C1 (n_40_6), .C2 (n_37_6) );
AOI211_X1 g_24_12 (.ZN (n_24_12), .A (n_28_12), .B (n_34_9), .C1 (n_38_7), .C2 (n_39_5) );
AOI211_X1 g_22_13 (.ZN (n_22_13), .A (n_26_11), .B (n_32_10), .C1 (n_36_8), .C2 (n_41_4) );
AOI211_X1 g_20_14 (.ZN (n_20_14), .A (n_24_12), .B (n_30_11), .C1 (n_34_9), .C2 (n_40_6) );
AOI211_X1 g_18_15 (.ZN (n_18_15), .A (n_22_13), .B (n_28_12), .C1 (n_32_10), .C2 (n_38_7) );
AOI211_X1 g_16_16 (.ZN (n_16_16), .A (n_20_14), .B (n_26_11), .C1 (n_30_11), .C2 (n_36_8) );
AOI211_X1 g_14_17 (.ZN (n_14_17), .A (n_18_15), .B (n_24_12), .C1 (n_28_12), .C2 (n_34_9) );
AOI211_X1 g_12_18 (.ZN (n_12_18), .A (n_16_16), .B (n_22_13), .C1 (n_26_11), .C2 (n_32_10) );
AOI211_X1 g_10_19 (.ZN (n_10_19), .A (n_14_17), .B (n_20_14), .C1 (n_24_12), .C2 (n_30_11) );
AOI211_X1 g_8_18 (.ZN (n_8_18), .A (n_12_18), .B (n_18_15), .C1 (n_22_13), .C2 (n_28_12) );
AOI211_X1 g_6_19 (.ZN (n_6_19), .A (n_10_19), .B (n_16_16), .C1 (n_20_14), .C2 (n_26_11) );
AOI211_X1 g_5_21 (.ZN (n_5_21), .A (n_8_18), .B (n_14_17), .C1 (n_18_15), .C2 (n_24_12) );
AOI211_X1 g_7_20 (.ZN (n_7_20), .A (n_6_19), .B (n_12_18), .C1 (n_16_16), .C2 (n_22_13) );
AOI211_X1 g_9_19 (.ZN (n_9_19), .A (n_5_21), .B (n_10_19), .C1 (n_14_17), .C2 (n_20_14) );
AOI211_X1 g_11_18 (.ZN (n_11_18), .A (n_7_20), .B (n_8_18), .C1 (n_12_18), .C2 (n_18_15) );
AOI211_X1 g_13_17 (.ZN (n_13_17), .A (n_9_19), .B (n_6_19), .C1 (n_10_19), .C2 (n_16_16) );
AOI211_X1 g_12_19 (.ZN (n_12_19), .A (n_11_18), .B (n_5_21), .C1 (n_8_18), .C2 (n_14_17) );
AOI211_X1 g_14_18 (.ZN (n_14_18), .A (n_13_17), .B (n_7_20), .C1 (n_6_19), .C2 (n_12_18) );
AOI211_X1 g_16_17 (.ZN (n_16_17), .A (n_12_19), .B (n_9_19), .C1 (n_5_21), .C2 (n_10_19) );
AOI211_X1 g_18_16 (.ZN (n_18_16), .A (n_14_18), .B (n_11_18), .C1 (n_7_20), .C2 (n_8_18) );
AOI211_X1 g_20_15 (.ZN (n_20_15), .A (n_16_17), .B (n_13_17), .C1 (n_9_19), .C2 (n_6_19) );
AOI211_X1 g_22_14 (.ZN (n_22_14), .A (n_18_16), .B (n_12_19), .C1 (n_11_18), .C2 (n_5_21) );
AOI211_X1 g_24_13 (.ZN (n_24_13), .A (n_20_15), .B (n_14_18), .C1 (n_13_17), .C2 (n_7_20) );
AOI211_X1 g_26_12 (.ZN (n_26_12), .A (n_22_14), .B (n_16_17), .C1 (n_12_19), .C2 (n_9_19) );
AOI211_X1 g_28_11 (.ZN (n_28_11), .A (n_24_13), .B (n_18_16), .C1 (n_14_18), .C2 (n_11_18) );
AOI211_X1 g_30_10 (.ZN (n_30_10), .A (n_26_12), .B (n_20_15), .C1 (n_16_17), .C2 (n_13_17) );
AOI211_X1 g_32_9 (.ZN (n_32_9), .A (n_28_11), .B (n_22_14), .C1 (n_18_16), .C2 (n_12_19) );
AOI211_X1 g_34_8 (.ZN (n_34_8), .A (n_30_10), .B (n_24_13), .C1 (n_20_15), .C2 (n_14_18) );
AOI211_X1 g_36_7 (.ZN (n_36_7), .A (n_32_9), .B (n_26_12), .C1 (n_22_14), .C2 (n_16_17) );
AOI211_X1 g_38_6 (.ZN (n_38_6), .A (n_34_8), .B (n_28_11), .C1 (n_24_13), .C2 (n_18_16) );
AOI211_X1 g_40_5 (.ZN (n_40_5), .A (n_36_7), .B (n_30_10), .C1 (n_26_12), .C2 (n_20_15) );
AOI211_X1 g_42_4 (.ZN (n_42_4), .A (n_38_6), .B (n_32_9), .C1 (n_28_11), .C2 (n_22_14) );
AOI211_X1 g_44_3 (.ZN (n_44_3), .A (n_40_5), .B (n_34_8), .C1 (n_30_10), .C2 (n_24_13) );
AOI211_X1 g_46_2 (.ZN (n_46_2), .A (n_42_4), .B (n_36_7), .C1 (n_32_9), .C2 (n_26_12) );
AOI211_X1 g_48_1 (.ZN (n_48_1), .A (n_44_3), .B (n_38_6), .C1 (n_34_8), .C2 (n_28_11) );
AOI211_X1 g_47_3 (.ZN (n_47_3), .A (n_46_2), .B (n_40_5), .C1 (n_36_7), .C2 (n_30_10) );
AOI211_X1 g_45_4 (.ZN (n_45_4), .A (n_48_1), .B (n_42_4), .C1 (n_38_6), .C2 (n_32_9) );
AOI211_X1 g_43_5 (.ZN (n_43_5), .A (n_47_3), .B (n_44_3), .C1 (n_40_5), .C2 (n_34_8) );
AOI211_X1 g_41_6 (.ZN (n_41_6), .A (n_45_4), .B (n_46_2), .C1 (n_42_4), .C2 (n_36_7) );
AOI211_X1 g_39_7 (.ZN (n_39_7), .A (n_43_5), .B (n_48_1), .C1 (n_44_3), .C2 (n_38_6) );
AOI211_X1 g_37_8 (.ZN (n_37_8), .A (n_41_6), .B (n_47_3), .C1 (n_46_2), .C2 (n_40_5) );
AOI211_X1 g_35_9 (.ZN (n_35_9), .A (n_39_7), .B (n_45_4), .C1 (n_48_1), .C2 (n_42_4) );
AOI211_X1 g_33_10 (.ZN (n_33_10), .A (n_37_8), .B (n_43_5), .C1 (n_47_3), .C2 (n_44_3) );
AOI211_X1 g_31_11 (.ZN (n_31_11), .A (n_35_9), .B (n_41_6), .C1 (n_45_4), .C2 (n_46_2) );
AOI211_X1 g_29_12 (.ZN (n_29_12), .A (n_33_10), .B (n_39_7), .C1 (n_43_5), .C2 (n_48_1) );
AOI211_X1 g_27_11 (.ZN (n_27_11), .A (n_31_11), .B (n_37_8), .C1 (n_41_6), .C2 (n_47_3) );
AOI211_X1 g_25_12 (.ZN (n_25_12), .A (n_29_12), .B (n_35_9), .C1 (n_39_7), .C2 (n_45_4) );
AOI211_X1 g_23_13 (.ZN (n_23_13), .A (n_27_11), .B (n_33_10), .C1 (n_37_8), .C2 (n_43_5) );
AOI211_X1 g_21_14 (.ZN (n_21_14), .A (n_25_12), .B (n_31_11), .C1 (n_35_9), .C2 (n_41_6) );
AOI211_X1 g_19_15 (.ZN (n_19_15), .A (n_23_13), .B (n_29_12), .C1 (n_33_10), .C2 (n_39_7) );
AOI211_X1 g_17_16 (.ZN (n_17_16), .A (n_21_14), .B (n_27_11), .C1 (n_31_11), .C2 (n_37_8) );
AOI211_X1 g_15_17 (.ZN (n_15_17), .A (n_19_15), .B (n_25_12), .C1 (n_29_12), .C2 (n_35_9) );
AOI211_X1 g_13_18 (.ZN (n_13_18), .A (n_17_16), .B (n_23_13), .C1 (n_27_11), .C2 (n_33_10) );
AOI211_X1 g_11_19 (.ZN (n_11_19), .A (n_15_17), .B (n_21_14), .C1 (n_25_12), .C2 (n_31_11) );
AOI211_X1 g_9_20 (.ZN (n_9_20), .A (n_13_18), .B (n_19_15), .C1 (n_23_13), .C2 (n_29_12) );
AOI211_X1 g_7_21 (.ZN (n_7_21), .A (n_11_19), .B (n_17_16), .C1 (n_21_14), .C2 (n_27_11) );
AOI211_X1 g_8_19 (.ZN (n_8_19), .A (n_9_20), .B (n_15_17), .C1 (n_19_15), .C2 (n_25_12) );
AOI211_X1 g_6_20 (.ZN (n_6_20), .A (n_7_21), .B (n_13_18), .C1 (n_17_16), .C2 (n_23_13) );
AOI211_X1 g_4_21 (.ZN (n_4_21), .A (n_8_19), .B (n_11_19), .C1 (n_15_17), .C2 (n_21_14) );
AOI211_X1 g_2_22 (.ZN (n_2_22), .A (n_6_20), .B (n_9_20), .C1 (n_13_18), .C2 (n_19_15) );
AOI211_X1 g_1_24 (.ZN (n_1_24), .A (n_4_21), .B (n_7_21), .C1 (n_11_19), .C2 (n_17_16) );
AOI211_X1 g_3_23 (.ZN (n_3_23), .A (n_2_22), .B (n_8_19), .C1 (n_9_20), .C2 (n_15_17) );
AOI211_X1 g_5_22 (.ZN (n_5_22), .A (n_1_24), .B (n_6_20), .C1 (n_7_21), .C2 (n_13_18) );
AOI211_X1 g_4_24 (.ZN (n_4_24), .A (n_3_23), .B (n_4_21), .C1 (n_8_19), .C2 (n_11_19) );
AOI211_X1 g_2_25 (.ZN (n_2_25), .A (n_5_22), .B (n_2_22), .C1 (n_6_20), .C2 (n_9_20) );
AOI211_X1 g_1_27 (.ZN (n_1_27), .A (n_4_24), .B (n_1_24), .C1 (n_4_21), .C2 (n_7_21) );
AOI211_X1 g_3_26 (.ZN (n_3_26), .A (n_2_25), .B (n_3_23), .C1 (n_2_22), .C2 (n_8_19) );
AOI211_X1 g_4_28 (.ZN (n_4_28), .A (n_1_27), .B (n_5_22), .C1 (n_1_24), .C2 (n_6_20) );
AOI211_X1 g_2_29 (.ZN (n_2_29), .A (n_3_26), .B (n_4_24), .C1 (n_3_23), .C2 (n_4_21) );
AOI211_X1 g_1_31 (.ZN (n_1_31), .A (n_4_28), .B (n_2_25), .C1 (n_5_22), .C2 (n_2_22) );
AOI211_X1 g_3_30 (.ZN (n_3_30), .A (n_2_29), .B (n_1_27), .C1 (n_4_24), .C2 (n_1_24) );
AOI211_X1 g_4_32 (.ZN (n_4_32), .A (n_1_31), .B (n_3_26), .C1 (n_2_25), .C2 (n_3_23) );
AOI211_X1 g_2_33 (.ZN (n_2_33), .A (n_3_30), .B (n_4_28), .C1 (n_1_27), .C2 (n_5_22) );
AOI211_X1 g_1_35 (.ZN (n_1_35), .A (n_4_32), .B (n_2_29), .C1 (n_3_26), .C2 (n_4_24) );
AOI211_X1 g_3_34 (.ZN (n_3_34), .A (n_2_33), .B (n_1_31), .C1 (n_4_28), .C2 (n_2_25) );
AOI211_X1 g_4_36 (.ZN (n_4_36), .A (n_1_35), .B (n_3_30), .C1 (n_2_29), .C2 (n_1_27) );
AOI211_X1 g_2_37 (.ZN (n_2_37), .A (n_3_34), .B (n_4_32), .C1 (n_1_31), .C2 (n_3_26) );
AOI211_X1 g_1_39 (.ZN (n_1_39), .A (n_4_36), .B (n_2_33), .C1 (n_3_30), .C2 (n_4_28) );
AOI211_X1 g_3_38 (.ZN (n_3_38), .A (n_2_37), .B (n_1_35), .C1 (n_4_32), .C2 (n_2_29) );
AOI211_X1 g_4_40 (.ZN (n_4_40), .A (n_1_39), .B (n_3_34), .C1 (n_2_33), .C2 (n_1_31) );
AOI211_X1 g_2_41 (.ZN (n_2_41), .A (n_3_38), .B (n_4_36), .C1 (n_1_35), .C2 (n_3_30) );
AOI211_X1 g_1_43 (.ZN (n_1_43), .A (n_4_40), .B (n_2_37), .C1 (n_3_34), .C2 (n_4_32) );
AOI211_X1 g_3_42 (.ZN (n_3_42), .A (n_2_41), .B (n_1_39), .C1 (n_4_36), .C2 (n_2_33) );
AOI211_X1 g_4_44 (.ZN (n_4_44), .A (n_1_43), .B (n_3_38), .C1 (n_2_37), .C2 (n_1_35) );
AOI211_X1 g_2_45 (.ZN (n_2_45), .A (n_3_42), .B (n_4_40), .C1 (n_1_39), .C2 (n_3_34) );
AOI211_X1 g_1_47 (.ZN (n_1_47), .A (n_4_44), .B (n_2_41), .C1 (n_3_38), .C2 (n_4_36) );
AOI211_X1 g_3_46 (.ZN (n_3_46), .A (n_2_45), .B (n_1_43), .C1 (n_4_40), .C2 (n_2_37) );
AOI211_X1 g_4_48 (.ZN (n_4_48), .A (n_1_47), .B (n_3_42), .C1 (n_2_41), .C2 (n_1_39) );
AOI211_X1 g_2_49 (.ZN (n_2_49), .A (n_3_46), .B (n_4_44), .C1 (n_1_43), .C2 (n_3_38) );
AOI211_X1 g_1_51 (.ZN (n_1_51), .A (n_4_48), .B (n_2_45), .C1 (n_3_42), .C2 (n_4_40) );
AOI211_X1 g_3_50 (.ZN (n_3_50), .A (n_2_49), .B (n_1_47), .C1 (n_4_44), .C2 (n_2_41) );
AOI211_X1 g_4_52 (.ZN (n_4_52), .A (n_1_51), .B (n_3_46), .C1 (n_2_45), .C2 (n_1_43) );
AOI211_X1 g_2_53 (.ZN (n_2_53), .A (n_3_50), .B (n_4_48), .C1 (n_1_47), .C2 (n_3_42) );
AOI211_X1 g_1_55 (.ZN (n_1_55), .A (n_4_52), .B (n_2_49), .C1 (n_3_46), .C2 (n_4_44) );
AOI211_X1 g_3_54 (.ZN (n_3_54), .A (n_2_53), .B (n_1_51), .C1 (n_4_48), .C2 (n_2_45) );
AOI211_X1 g_4_56 (.ZN (n_4_56), .A (n_1_55), .B (n_3_50), .C1 (n_2_49), .C2 (n_1_47) );
AOI211_X1 g_2_57 (.ZN (n_2_57), .A (n_3_54), .B (n_4_52), .C1 (n_1_51), .C2 (n_3_46) );
AOI211_X1 g_1_59 (.ZN (n_1_59), .A (n_4_56), .B (n_2_53), .C1 (n_3_50), .C2 (n_4_48) );
AOI211_X1 g_3_58 (.ZN (n_3_58), .A (n_2_57), .B (n_1_55), .C1 (n_4_52), .C2 (n_2_49) );
AOI211_X1 g_4_60 (.ZN (n_4_60), .A (n_1_59), .B (n_3_54), .C1 (n_2_53), .C2 (n_1_51) );
AOI211_X1 g_2_61 (.ZN (n_2_61), .A (n_3_58), .B (n_4_56), .C1 (n_1_55), .C2 (n_3_50) );
AOI211_X1 g_1_63 (.ZN (n_1_63), .A (n_4_60), .B (n_2_57), .C1 (n_3_54), .C2 (n_4_52) );
AOI211_X1 g_3_62 (.ZN (n_3_62), .A (n_2_61), .B (n_1_59), .C1 (n_4_56), .C2 (n_2_53) );
AOI211_X1 g_4_64 (.ZN (n_4_64), .A (n_1_63), .B (n_3_58), .C1 (n_2_57), .C2 (n_1_55) );
AOI211_X1 g_2_65 (.ZN (n_2_65), .A (n_3_62), .B (n_4_60), .C1 (n_1_59), .C2 (n_3_54) );
AOI211_X1 g_1_67 (.ZN (n_1_67), .A (n_4_64), .B (n_2_61), .C1 (n_3_58), .C2 (n_4_56) );
AOI211_X1 g_3_66 (.ZN (n_3_66), .A (n_2_65), .B (n_1_63), .C1 (n_4_60), .C2 (n_2_57) );
AOI211_X1 g_4_68 (.ZN (n_4_68), .A (n_1_67), .B (n_3_62), .C1 (n_2_61), .C2 (n_1_59) );
AOI211_X1 g_2_69 (.ZN (n_2_69), .A (n_3_66), .B (n_4_64), .C1 (n_1_63), .C2 (n_3_58) );
AOI211_X1 g_1_71 (.ZN (n_1_71), .A (n_4_68), .B (n_2_65), .C1 (n_3_62), .C2 (n_4_60) );
AOI211_X1 g_3_70 (.ZN (n_3_70), .A (n_2_69), .B (n_1_67), .C1 (n_4_64), .C2 (n_2_61) );
AOI211_X1 g_4_72 (.ZN (n_4_72), .A (n_1_71), .B (n_3_66), .C1 (n_2_65), .C2 (n_1_63) );
AOI211_X1 g_2_73 (.ZN (n_2_73), .A (n_3_70), .B (n_4_68), .C1 (n_1_67), .C2 (n_3_62) );
AOI211_X1 g_1_75 (.ZN (n_1_75), .A (n_4_72), .B (n_2_69), .C1 (n_3_66), .C2 (n_4_64) );
AOI211_X1 g_3_74 (.ZN (n_3_74), .A (n_2_73), .B (n_1_71), .C1 (n_4_68), .C2 (n_2_65) );
AOI211_X1 g_4_76 (.ZN (n_4_76), .A (n_1_75), .B (n_3_70), .C1 (n_2_69), .C2 (n_1_67) );
AOI211_X1 g_2_77 (.ZN (n_2_77), .A (n_3_74), .B (n_4_72), .C1 (n_1_71), .C2 (n_3_66) );
AOI211_X1 g_1_79 (.ZN (n_1_79), .A (n_4_76), .B (n_2_73), .C1 (n_3_70), .C2 (n_4_68) );
AOI211_X1 g_3_78 (.ZN (n_3_78), .A (n_2_77), .B (n_1_75), .C1 (n_4_72), .C2 (n_2_69) );
AOI211_X1 g_4_80 (.ZN (n_4_80), .A (n_1_79), .B (n_3_74), .C1 (n_2_73), .C2 (n_1_71) );
AOI211_X1 g_2_81 (.ZN (n_2_81), .A (n_3_78), .B (n_4_76), .C1 (n_1_75), .C2 (n_3_70) );
AOI211_X1 g_1_83 (.ZN (n_1_83), .A (n_4_80), .B (n_2_77), .C1 (n_3_74), .C2 (n_4_72) );
AOI211_X1 g_3_82 (.ZN (n_3_82), .A (n_2_81), .B (n_1_79), .C1 (n_4_76), .C2 (n_2_73) );
AOI211_X1 g_4_84 (.ZN (n_4_84), .A (n_1_83), .B (n_3_78), .C1 (n_2_77), .C2 (n_1_75) );
AOI211_X1 g_2_85 (.ZN (n_2_85), .A (n_3_82), .B (n_4_80), .C1 (n_1_79), .C2 (n_3_74) );
AOI211_X1 g_1_87 (.ZN (n_1_87), .A (n_4_84), .B (n_2_81), .C1 (n_3_78), .C2 (n_4_76) );
AOI211_X1 g_3_86 (.ZN (n_3_86), .A (n_2_85), .B (n_1_83), .C1 (n_4_80), .C2 (n_2_77) );
AOI211_X1 g_4_88 (.ZN (n_4_88), .A (n_1_87), .B (n_3_82), .C1 (n_2_81), .C2 (n_1_79) );
AOI211_X1 g_2_89 (.ZN (n_2_89), .A (n_3_86), .B (n_4_84), .C1 (n_1_83), .C2 (n_3_78) );
AOI211_X1 g_1_91 (.ZN (n_1_91), .A (n_4_88), .B (n_2_85), .C1 (n_3_82), .C2 (n_4_80) );
AOI211_X1 g_3_90 (.ZN (n_3_90), .A (n_2_89), .B (n_1_87), .C1 (n_4_84), .C2 (n_2_81) );
AOI211_X1 g_4_92 (.ZN (n_4_92), .A (n_1_91), .B (n_3_86), .C1 (n_2_85), .C2 (n_1_83) );
AOI211_X1 g_2_93 (.ZN (n_2_93), .A (n_3_90), .B (n_4_88), .C1 (n_1_87), .C2 (n_3_82) );
AOI211_X1 g_1_95 (.ZN (n_1_95), .A (n_4_92), .B (n_2_89), .C1 (n_3_86), .C2 (n_4_84) );
AOI211_X1 g_3_94 (.ZN (n_3_94), .A (n_2_93), .B (n_1_91), .C1 (n_4_88), .C2 (n_2_85) );
AOI211_X1 g_4_96 (.ZN (n_4_96), .A (n_1_95), .B (n_3_90), .C1 (n_2_89), .C2 (n_1_87) );
AOI211_X1 g_2_97 (.ZN (n_2_97), .A (n_3_94), .B (n_4_92), .C1 (n_1_91), .C2 (n_3_86) );
AOI211_X1 g_1_99 (.ZN (n_1_99), .A (n_4_96), .B (n_2_93), .C1 (n_3_90), .C2 (n_4_88) );
AOI211_X1 g_3_98 (.ZN (n_3_98), .A (n_2_97), .B (n_1_95), .C1 (n_4_92), .C2 (n_2_89) );
AOI211_X1 g_4_100 (.ZN (n_4_100), .A (n_1_99), .B (n_3_94), .C1 (n_2_93), .C2 (n_1_91) );
AOI211_X1 g_2_101 (.ZN (n_2_101), .A (n_3_98), .B (n_4_96), .C1 (n_1_95), .C2 (n_3_90) );
AOI211_X1 g_1_103 (.ZN (n_1_103), .A (n_4_100), .B (n_2_97), .C1 (n_3_94), .C2 (n_4_92) );
AOI211_X1 g_3_102 (.ZN (n_3_102), .A (n_2_101), .B (n_1_99), .C1 (n_4_96), .C2 (n_2_93) );
AOI211_X1 g_4_104 (.ZN (n_4_104), .A (n_1_103), .B (n_3_98), .C1 (n_2_97), .C2 (n_1_95) );
AOI211_X1 g_2_105 (.ZN (n_2_105), .A (n_3_102), .B (n_4_100), .C1 (n_1_99), .C2 (n_3_94) );
AOI211_X1 g_1_107 (.ZN (n_1_107), .A (n_4_104), .B (n_2_101), .C1 (n_3_98), .C2 (n_4_96) );
AOI211_X1 g_3_106 (.ZN (n_3_106), .A (n_2_105), .B (n_1_103), .C1 (n_4_100), .C2 (n_2_97) );
AOI211_X1 g_4_108 (.ZN (n_4_108), .A (n_1_107), .B (n_3_102), .C1 (n_2_101), .C2 (n_1_99) );
AOI211_X1 g_2_109 (.ZN (n_2_109), .A (n_3_106), .B (n_4_104), .C1 (n_1_103), .C2 (n_3_98) );
AOI211_X1 g_1_111 (.ZN (n_1_111), .A (n_4_108), .B (n_2_105), .C1 (n_3_102), .C2 (n_4_100) );
AOI211_X1 g_3_110 (.ZN (n_3_110), .A (n_2_109), .B (n_1_107), .C1 (n_4_104), .C2 (n_2_101) );
AOI211_X1 g_4_112 (.ZN (n_4_112), .A (n_1_111), .B (n_3_106), .C1 (n_2_105), .C2 (n_1_103) );
AOI211_X1 g_2_113 (.ZN (n_2_113), .A (n_3_110), .B (n_4_108), .C1 (n_1_107), .C2 (n_3_102) );
AOI211_X1 g_1_115 (.ZN (n_1_115), .A (n_4_112), .B (n_2_109), .C1 (n_3_106), .C2 (n_4_104) );
AOI211_X1 g_3_114 (.ZN (n_3_114), .A (n_2_113), .B (n_1_111), .C1 (n_4_108), .C2 (n_2_105) );
AOI211_X1 g_4_116 (.ZN (n_4_116), .A (n_1_115), .B (n_3_110), .C1 (n_2_109), .C2 (n_1_107) );
AOI211_X1 g_2_117 (.ZN (n_2_117), .A (n_3_114), .B (n_4_112), .C1 (n_1_111), .C2 (n_3_106) );
AOI211_X1 g_1_119 (.ZN (n_1_119), .A (n_4_116), .B (n_2_113), .C1 (n_3_110), .C2 (n_4_108) );
AOI211_X1 g_3_118 (.ZN (n_3_118), .A (n_2_117), .B (n_1_115), .C1 (n_4_112), .C2 (n_2_109) );
AOI211_X1 g_4_120 (.ZN (n_4_120), .A (n_1_119), .B (n_3_114), .C1 (n_2_113), .C2 (n_1_111) );
AOI211_X1 g_2_121 (.ZN (n_2_121), .A (n_3_118), .B (n_4_116), .C1 (n_1_115), .C2 (n_3_110) );
AOI211_X1 g_1_123 (.ZN (n_1_123), .A (n_4_120), .B (n_2_117), .C1 (n_3_114), .C2 (n_4_112) );
AOI211_X1 g_3_122 (.ZN (n_3_122), .A (n_2_121), .B (n_1_119), .C1 (n_4_116), .C2 (n_2_113) );
AOI211_X1 g_4_124 (.ZN (n_4_124), .A (n_1_123), .B (n_3_118), .C1 (n_2_117), .C2 (n_1_115) );
AOI211_X1 g_2_125 (.ZN (n_2_125), .A (n_3_122), .B (n_4_120), .C1 (n_1_119), .C2 (n_3_114) );
AOI211_X1 g_1_127 (.ZN (n_1_127), .A (n_4_124), .B (n_2_121), .C1 (n_3_118), .C2 (n_4_116) );
AOI211_X1 g_3_126 (.ZN (n_3_126), .A (n_2_125), .B (n_1_123), .C1 (n_4_120), .C2 (n_2_117) );
AOI211_X1 g_4_128 (.ZN (n_4_128), .A (n_1_127), .B (n_3_122), .C1 (n_2_121), .C2 (n_1_119) );
AOI211_X1 g_2_129 (.ZN (n_2_129), .A (n_3_126), .B (n_4_124), .C1 (n_1_123), .C2 (n_3_118) );
AOI211_X1 g_1_131 (.ZN (n_1_131), .A (n_4_128), .B (n_2_125), .C1 (n_3_122), .C2 (n_4_120) );
AOI211_X1 g_3_130 (.ZN (n_3_130), .A (n_2_129), .B (n_1_127), .C1 (n_4_124), .C2 (n_2_121) );
AOI211_X1 g_4_132 (.ZN (n_4_132), .A (n_1_131), .B (n_3_126), .C1 (n_2_125), .C2 (n_1_123) );
AOI211_X1 g_2_133 (.ZN (n_2_133), .A (n_3_130), .B (n_4_128), .C1 (n_1_127), .C2 (n_3_122) );
AOI211_X1 g_1_135 (.ZN (n_1_135), .A (n_4_132), .B (n_2_129), .C1 (n_3_126), .C2 (n_4_124) );
AOI211_X1 g_3_134 (.ZN (n_3_134), .A (n_2_133), .B (n_1_131), .C1 (n_4_128), .C2 (n_2_125) );
AOI211_X1 g_4_136 (.ZN (n_4_136), .A (n_1_135), .B (n_3_130), .C1 (n_2_129), .C2 (n_1_127) );
AOI211_X1 g_2_137 (.ZN (n_2_137), .A (n_3_134), .B (n_4_132), .C1 (n_1_131), .C2 (n_3_126) );
AOI211_X1 g_1_139 (.ZN (n_1_139), .A (n_4_136), .B (n_2_133), .C1 (n_3_130), .C2 (n_4_128) );
AOI211_X1 g_3_138 (.ZN (n_3_138), .A (n_2_137), .B (n_1_135), .C1 (n_4_132), .C2 (n_2_129) );
AOI211_X1 g_4_140 (.ZN (n_4_140), .A (n_1_139), .B (n_3_134), .C1 (n_2_133), .C2 (n_1_131) );
AOI211_X1 g_2_141 (.ZN (n_2_141), .A (n_3_138), .B (n_4_136), .C1 (n_1_135), .C2 (n_3_130) );
AOI211_X1 g_1_143 (.ZN (n_1_143), .A (n_4_140), .B (n_2_137), .C1 (n_3_134), .C2 (n_4_132) );
AOI211_X1 g_3_142 (.ZN (n_3_142), .A (n_2_141), .B (n_1_139), .C1 (n_4_136), .C2 (n_2_133) );
AOI211_X1 g_4_144 (.ZN (n_4_144), .A (n_1_143), .B (n_3_138), .C1 (n_2_137), .C2 (n_1_135) );
AOI211_X1 g_2_145 (.ZN (n_2_145), .A (n_3_142), .B (n_4_140), .C1 (n_1_139), .C2 (n_3_134) );
AOI211_X1 g_1_147 (.ZN (n_1_147), .A (n_4_144), .B (n_2_141), .C1 (n_3_138), .C2 (n_4_136) );
AOI211_X1 g_3_146 (.ZN (n_3_146), .A (n_2_145), .B (n_1_143), .C1 (n_4_140), .C2 (n_2_137) );
AOI211_X1 g_4_148 (.ZN (n_4_148), .A (n_1_147), .B (n_3_142), .C1 (n_2_141), .C2 (n_1_139) );
AOI211_X1 g_2_149 (.ZN (n_2_149), .A (n_3_146), .B (n_4_144), .C1 (n_1_143), .C2 (n_3_138) );
AOI211_X1 g_4_150 (.ZN (n_4_150), .A (n_4_148), .B (n_2_145), .C1 (n_3_142), .C2 (n_4_140) );
AOI211_X1 g_6_149 (.ZN (n_6_149), .A (n_2_149), .B (n_1_147), .C1 (n_4_144), .C2 (n_2_141) );
AOI211_X1 g_8_150 (.ZN (n_8_150), .A (n_4_150), .B (n_3_146), .C1 (n_2_145), .C2 (n_1_143) );
AOI211_X1 g_10_149 (.ZN (n_10_149), .A (n_6_149), .B (n_4_148), .C1 (n_1_147), .C2 (n_3_142) );
AOI211_X1 g_12_150 (.ZN (n_12_150), .A (n_8_150), .B (n_2_149), .C1 (n_3_146), .C2 (n_4_144) );
AOI211_X1 g_14_149 (.ZN (n_14_149), .A (n_10_149), .B (n_4_150), .C1 (n_4_148), .C2 (n_2_145) );
AOI211_X1 g_16_150 (.ZN (n_16_150), .A (n_12_150), .B (n_6_149), .C1 (n_2_149), .C2 (n_1_147) );
AOI211_X1 g_18_149 (.ZN (n_18_149), .A (n_14_149), .B (n_8_150), .C1 (n_4_150), .C2 (n_3_146) );
AOI211_X1 g_20_150 (.ZN (n_20_150), .A (n_16_150), .B (n_10_149), .C1 (n_6_149), .C2 (n_4_148) );
AOI211_X1 g_22_149 (.ZN (n_22_149), .A (n_18_149), .B (n_12_150), .C1 (n_8_150), .C2 (n_2_149) );
AOI211_X1 g_24_150 (.ZN (n_24_150), .A (n_20_150), .B (n_14_149), .C1 (n_10_149), .C2 (n_4_150) );
AOI211_X1 g_26_149 (.ZN (n_26_149), .A (n_22_149), .B (n_16_150), .C1 (n_12_150), .C2 (n_6_149) );
AOI211_X1 g_28_150 (.ZN (n_28_150), .A (n_24_150), .B (n_18_149), .C1 (n_14_149), .C2 (n_8_150) );
AOI211_X1 g_30_149 (.ZN (n_30_149), .A (n_26_149), .B (n_20_150), .C1 (n_16_150), .C2 (n_10_149) );
AOI211_X1 g_32_150 (.ZN (n_32_150), .A (n_28_150), .B (n_22_149), .C1 (n_18_149), .C2 (n_12_150) );
AOI211_X1 g_34_149 (.ZN (n_34_149), .A (n_30_149), .B (n_24_150), .C1 (n_20_150), .C2 (n_14_149) );
AOI211_X1 g_36_150 (.ZN (n_36_150), .A (n_32_150), .B (n_26_149), .C1 (n_22_149), .C2 (n_16_150) );
AOI211_X1 g_38_149 (.ZN (n_38_149), .A (n_34_149), .B (n_28_150), .C1 (n_24_150), .C2 (n_18_149) );
AOI211_X1 g_40_150 (.ZN (n_40_150), .A (n_36_150), .B (n_30_149), .C1 (n_26_149), .C2 (n_20_150) );
AOI211_X1 g_42_149 (.ZN (n_42_149), .A (n_38_149), .B (n_32_150), .C1 (n_28_150), .C2 (n_22_149) );
AOI211_X1 g_44_150 (.ZN (n_44_150), .A (n_40_150), .B (n_34_149), .C1 (n_30_149), .C2 (n_24_150) );
AOI211_X1 g_46_149 (.ZN (n_46_149), .A (n_42_149), .B (n_36_150), .C1 (n_32_150), .C2 (n_26_149) );
AOI211_X1 g_48_150 (.ZN (n_48_150), .A (n_44_150), .B (n_38_149), .C1 (n_34_149), .C2 (n_28_150) );
AOI211_X1 g_50_149 (.ZN (n_50_149), .A (n_46_149), .B (n_40_150), .C1 (n_36_150), .C2 (n_30_149) );
AOI211_X1 g_52_150 (.ZN (n_52_150), .A (n_48_150), .B (n_42_149), .C1 (n_38_149), .C2 (n_32_150) );
AOI211_X1 g_54_149 (.ZN (n_54_149), .A (n_50_149), .B (n_44_150), .C1 (n_40_150), .C2 (n_34_149) );
AOI211_X1 g_56_150 (.ZN (n_56_150), .A (n_52_150), .B (n_46_149), .C1 (n_42_149), .C2 (n_36_150) );
AOI211_X1 g_58_149 (.ZN (n_58_149), .A (n_54_149), .B (n_48_150), .C1 (n_44_150), .C2 (n_38_149) );
AOI211_X1 g_60_150 (.ZN (n_60_150), .A (n_56_150), .B (n_50_149), .C1 (n_46_149), .C2 (n_40_150) );
AOI211_X1 g_62_149 (.ZN (n_62_149), .A (n_58_149), .B (n_52_150), .C1 (n_48_150), .C2 (n_42_149) );
AOI211_X1 g_64_150 (.ZN (n_64_150), .A (n_60_150), .B (n_54_149), .C1 (n_50_149), .C2 (n_44_150) );
AOI211_X1 g_66_149 (.ZN (n_66_149), .A (n_62_149), .B (n_56_150), .C1 (n_52_150), .C2 (n_46_149) );
AOI211_X1 g_68_150 (.ZN (n_68_150), .A (n_64_150), .B (n_58_149), .C1 (n_54_149), .C2 (n_48_150) );
AOI211_X1 g_70_149 (.ZN (n_70_149), .A (n_66_149), .B (n_60_150), .C1 (n_56_150), .C2 (n_50_149) );
AOI211_X1 g_72_150 (.ZN (n_72_150), .A (n_68_150), .B (n_62_149), .C1 (n_58_149), .C2 (n_52_150) );
AOI211_X1 g_74_149 (.ZN (n_74_149), .A (n_70_149), .B (n_64_150), .C1 (n_60_150), .C2 (n_54_149) );
AOI211_X1 g_76_150 (.ZN (n_76_150), .A (n_72_150), .B (n_66_149), .C1 (n_62_149), .C2 (n_56_150) );
AOI211_X1 g_78_149 (.ZN (n_78_149), .A (n_74_149), .B (n_68_150), .C1 (n_64_150), .C2 (n_58_149) );
AOI211_X1 g_80_150 (.ZN (n_80_150), .A (n_76_150), .B (n_70_149), .C1 (n_66_149), .C2 (n_60_150) );
AOI211_X1 g_82_149 (.ZN (n_82_149), .A (n_78_149), .B (n_72_150), .C1 (n_68_150), .C2 (n_62_149) );
AOI211_X1 g_84_150 (.ZN (n_84_150), .A (n_80_150), .B (n_74_149), .C1 (n_70_149), .C2 (n_64_150) );
AOI211_X1 g_86_149 (.ZN (n_86_149), .A (n_82_149), .B (n_76_150), .C1 (n_72_150), .C2 (n_66_149) );
AOI211_X1 g_88_150 (.ZN (n_88_150), .A (n_84_150), .B (n_78_149), .C1 (n_74_149), .C2 (n_68_150) );
AOI211_X1 g_90_149 (.ZN (n_90_149), .A (n_86_149), .B (n_80_150), .C1 (n_76_150), .C2 (n_70_149) );
AOI211_X1 g_92_150 (.ZN (n_92_150), .A (n_88_150), .B (n_82_149), .C1 (n_78_149), .C2 (n_72_150) );
AOI211_X1 g_94_149 (.ZN (n_94_149), .A (n_90_149), .B (n_84_150), .C1 (n_80_150), .C2 (n_74_149) );
AOI211_X1 g_96_150 (.ZN (n_96_150), .A (n_92_150), .B (n_86_149), .C1 (n_82_149), .C2 (n_76_150) );
AOI211_X1 g_98_149 (.ZN (n_98_149), .A (n_94_149), .B (n_88_150), .C1 (n_84_150), .C2 (n_78_149) );
AOI211_X1 g_100_150 (.ZN (n_100_150), .A (n_96_150), .B (n_90_149), .C1 (n_86_149), .C2 (n_80_150) );
AOI211_X1 g_102_149 (.ZN (n_102_149), .A (n_98_149), .B (n_92_150), .C1 (n_88_150), .C2 (n_82_149) );
AOI211_X1 g_104_150 (.ZN (n_104_150), .A (n_100_150), .B (n_94_149), .C1 (n_90_149), .C2 (n_84_150) );
AOI211_X1 g_106_149 (.ZN (n_106_149), .A (n_102_149), .B (n_96_150), .C1 (n_92_150), .C2 (n_86_149) );
AOI211_X1 g_108_150 (.ZN (n_108_150), .A (n_104_150), .B (n_98_149), .C1 (n_94_149), .C2 (n_88_150) );
AOI211_X1 g_110_149 (.ZN (n_110_149), .A (n_106_149), .B (n_100_150), .C1 (n_96_150), .C2 (n_90_149) );
AOI211_X1 g_112_150 (.ZN (n_112_150), .A (n_108_150), .B (n_102_149), .C1 (n_98_149), .C2 (n_92_150) );
AOI211_X1 g_114_149 (.ZN (n_114_149), .A (n_110_149), .B (n_104_150), .C1 (n_100_150), .C2 (n_94_149) );
AOI211_X1 g_116_150 (.ZN (n_116_150), .A (n_112_150), .B (n_106_149), .C1 (n_102_149), .C2 (n_96_150) );
AOI211_X1 g_118_149 (.ZN (n_118_149), .A (n_114_149), .B (n_108_150), .C1 (n_104_150), .C2 (n_98_149) );
AOI211_X1 g_120_150 (.ZN (n_120_150), .A (n_116_150), .B (n_110_149), .C1 (n_106_149), .C2 (n_100_150) );
AOI211_X1 g_122_149 (.ZN (n_122_149), .A (n_118_149), .B (n_112_150), .C1 (n_108_150), .C2 (n_102_149) );
AOI211_X1 g_124_150 (.ZN (n_124_150), .A (n_120_150), .B (n_114_149), .C1 (n_110_149), .C2 (n_104_150) );
AOI211_X1 g_126_149 (.ZN (n_126_149), .A (n_122_149), .B (n_116_150), .C1 (n_112_150), .C2 (n_106_149) );
AOI211_X1 g_128_150 (.ZN (n_128_150), .A (n_124_150), .B (n_118_149), .C1 (n_114_149), .C2 (n_108_150) );
AOI211_X1 g_130_149 (.ZN (n_130_149), .A (n_126_149), .B (n_120_150), .C1 (n_116_150), .C2 (n_110_149) );
AOI211_X1 g_132_150 (.ZN (n_132_150), .A (n_128_150), .B (n_122_149), .C1 (n_118_149), .C2 (n_112_150) );
AOI211_X1 g_134_149 (.ZN (n_134_149), .A (n_130_149), .B (n_124_150), .C1 (n_120_150), .C2 (n_114_149) );
AOI211_X1 g_136_150 (.ZN (n_136_150), .A (n_132_150), .B (n_126_149), .C1 (n_122_149), .C2 (n_116_150) );
AOI211_X1 g_138_149 (.ZN (n_138_149), .A (n_134_149), .B (n_128_150), .C1 (n_124_150), .C2 (n_118_149) );
AOI211_X1 g_140_150 (.ZN (n_140_150), .A (n_136_150), .B (n_130_149), .C1 (n_126_149), .C2 (n_120_150) );
AOI211_X1 g_142_149 (.ZN (n_142_149), .A (n_138_149), .B (n_132_150), .C1 (n_128_150), .C2 (n_122_149) );
AOI211_X1 g_140_148 (.ZN (n_140_148), .A (n_140_150), .B (n_134_149), .C1 (n_130_149), .C2 (n_124_150) );
AOI211_X1 g_142_147 (.ZN (n_142_147), .A (n_142_149), .B (n_136_150), .C1 (n_132_150), .C2 (n_126_149) );
AOI211_X1 g_144_146 (.ZN (n_144_146), .A (n_140_148), .B (n_138_149), .C1 (n_134_149), .C2 (n_128_150) );
AOI211_X1 g_143_148 (.ZN (n_143_148), .A (n_142_147), .B (n_140_150), .C1 (n_136_150), .C2 (n_130_149) );
AOI211_X1 g_142_150 (.ZN (n_142_150), .A (n_144_146), .B (n_142_149), .C1 (n_138_149), .C2 (n_132_150) );
AOI211_X1 g_144_149 (.ZN (n_144_149), .A (n_143_148), .B (n_140_148), .C1 (n_140_150), .C2 (n_134_149) );
AOI211_X1 g_146_148 (.ZN (n_146_148), .A (n_142_150), .B (n_142_147), .C1 (n_142_149), .C2 (n_136_150) );
AOI211_X1 g_148_147 (.ZN (n_148_147), .A (n_144_149), .B (n_144_146), .C1 (n_140_148), .C2 (n_138_149) );
AOI211_X1 g_149_145 (.ZN (n_149_145), .A (n_146_148), .B (n_143_148), .C1 (n_142_147), .C2 (n_140_150) );
AOI211_X1 g_150_143 (.ZN (n_150_143), .A (n_148_147), .B (n_142_150), .C1 (n_144_146), .C2 (n_142_149) );
AOI211_X1 g_148_144 (.ZN (n_148_144), .A (n_149_145), .B (n_144_149), .C1 (n_143_148), .C2 (n_140_148) );
AOI211_X1 g_147_146 (.ZN (n_147_146), .A (n_150_143), .B (n_146_148), .C1 (n_142_150), .C2 (n_142_147) );
AOI211_X1 g_145_147 (.ZN (n_145_147), .A (n_148_144), .B (n_148_147), .C1 (n_144_149), .C2 (n_144_146) );
AOI211_X1 g_146_145 (.ZN (n_146_145), .A (n_147_146), .B (n_149_145), .C1 (n_146_148), .C2 (n_143_148) );
AOI211_X1 g_147_143 (.ZN (n_147_143), .A (n_145_147), .B (n_150_143), .C1 (n_148_147), .C2 (n_142_150) );
AOI211_X1 g_148_141 (.ZN (n_148_141), .A (n_146_145), .B (n_148_144), .C1 (n_149_145), .C2 (n_144_149) );
AOI211_X1 g_149_143 (.ZN (n_149_143), .A (n_147_143), .B (n_147_146), .C1 (n_150_143), .C2 (n_146_148) );
AOI211_X1 g_150_141 (.ZN (n_150_141), .A (n_148_141), .B (n_145_147), .C1 (n_148_144), .C2 (n_148_147) );
AOI211_X1 g_149_139 (.ZN (n_149_139), .A (n_149_143), .B (n_146_145), .C1 (n_147_146), .C2 (n_149_145) );
AOI211_X1 g_150_137 (.ZN (n_150_137), .A (n_150_141), .B (n_147_143), .C1 (n_145_147), .C2 (n_150_143) );
AOI211_X1 g_149_135 (.ZN (n_149_135), .A (n_149_139), .B (n_148_141), .C1 (n_146_145), .C2 (n_148_144) );
AOI211_X1 g_150_133 (.ZN (n_150_133), .A (n_150_137), .B (n_149_143), .C1 (n_147_143), .C2 (n_147_146) );
AOI211_X1 g_149_131 (.ZN (n_149_131), .A (n_149_135), .B (n_150_141), .C1 (n_148_141), .C2 (n_145_147) );
AOI211_X1 g_150_129 (.ZN (n_150_129), .A (n_150_133), .B (n_149_139), .C1 (n_149_143), .C2 (n_146_145) );
AOI211_X1 g_149_127 (.ZN (n_149_127), .A (n_149_131), .B (n_150_137), .C1 (n_150_141), .C2 (n_147_143) );
AOI211_X1 g_150_125 (.ZN (n_150_125), .A (n_150_129), .B (n_149_135), .C1 (n_149_139), .C2 (n_148_141) );
AOI211_X1 g_149_123 (.ZN (n_149_123), .A (n_149_127), .B (n_150_133), .C1 (n_150_137), .C2 (n_149_143) );
AOI211_X1 g_150_121 (.ZN (n_150_121), .A (n_150_125), .B (n_149_131), .C1 (n_149_135), .C2 (n_150_141) );
AOI211_X1 g_149_119 (.ZN (n_149_119), .A (n_149_123), .B (n_150_129), .C1 (n_150_133), .C2 (n_149_139) );
AOI211_X1 g_150_117 (.ZN (n_150_117), .A (n_150_121), .B (n_149_127), .C1 (n_149_131), .C2 (n_150_137) );
AOI211_X1 g_149_115 (.ZN (n_149_115), .A (n_149_119), .B (n_150_125), .C1 (n_150_129), .C2 (n_149_135) );
AOI211_X1 g_150_113 (.ZN (n_150_113), .A (n_150_117), .B (n_149_123), .C1 (n_149_127), .C2 (n_150_133) );
AOI211_X1 g_149_111 (.ZN (n_149_111), .A (n_149_115), .B (n_150_121), .C1 (n_150_125), .C2 (n_149_131) );
AOI211_X1 g_150_109 (.ZN (n_150_109), .A (n_150_113), .B (n_149_119), .C1 (n_149_123), .C2 (n_150_129) );
AOI211_X1 g_149_107 (.ZN (n_149_107), .A (n_149_111), .B (n_150_117), .C1 (n_150_121), .C2 (n_149_127) );
AOI211_X1 g_150_105 (.ZN (n_150_105), .A (n_150_109), .B (n_149_115), .C1 (n_149_119), .C2 (n_150_125) );
AOI211_X1 g_149_103 (.ZN (n_149_103), .A (n_149_107), .B (n_150_113), .C1 (n_150_117), .C2 (n_149_123) );
AOI211_X1 g_150_101 (.ZN (n_150_101), .A (n_150_105), .B (n_149_111), .C1 (n_149_115), .C2 (n_150_121) );
AOI211_X1 g_149_99 (.ZN (n_149_99), .A (n_149_103), .B (n_150_109), .C1 (n_150_113), .C2 (n_149_119) );
AOI211_X1 g_150_97 (.ZN (n_150_97), .A (n_150_101), .B (n_149_107), .C1 (n_149_111), .C2 (n_150_117) );
AOI211_X1 g_149_95 (.ZN (n_149_95), .A (n_149_99), .B (n_150_105), .C1 (n_150_109), .C2 (n_149_115) );
AOI211_X1 g_150_93 (.ZN (n_150_93), .A (n_150_97), .B (n_149_103), .C1 (n_149_107), .C2 (n_150_113) );
AOI211_X1 g_149_91 (.ZN (n_149_91), .A (n_149_95), .B (n_150_101), .C1 (n_150_105), .C2 (n_149_111) );
AOI211_X1 g_150_89 (.ZN (n_150_89), .A (n_150_93), .B (n_149_99), .C1 (n_149_103), .C2 (n_150_109) );
AOI211_X1 g_149_87 (.ZN (n_149_87), .A (n_149_91), .B (n_150_97), .C1 (n_150_101), .C2 (n_149_107) );
AOI211_X1 g_150_85 (.ZN (n_150_85), .A (n_150_89), .B (n_149_95), .C1 (n_149_99), .C2 (n_150_105) );
AOI211_X1 g_149_83 (.ZN (n_149_83), .A (n_149_87), .B (n_150_93), .C1 (n_150_97), .C2 (n_149_103) );
AOI211_X1 g_150_81 (.ZN (n_150_81), .A (n_150_85), .B (n_149_91), .C1 (n_149_95), .C2 (n_150_101) );
AOI211_X1 g_149_79 (.ZN (n_149_79), .A (n_149_83), .B (n_150_89), .C1 (n_150_93), .C2 (n_149_99) );
AOI211_X1 g_150_77 (.ZN (n_150_77), .A (n_150_81), .B (n_149_87), .C1 (n_149_91), .C2 (n_150_97) );
AOI211_X1 g_149_75 (.ZN (n_149_75), .A (n_149_79), .B (n_150_85), .C1 (n_150_89), .C2 (n_149_95) );
AOI211_X1 g_150_73 (.ZN (n_150_73), .A (n_150_77), .B (n_149_83), .C1 (n_149_87), .C2 (n_150_93) );
AOI211_X1 g_149_71 (.ZN (n_149_71), .A (n_149_75), .B (n_150_81), .C1 (n_150_85), .C2 (n_149_91) );
AOI211_X1 g_150_69 (.ZN (n_150_69), .A (n_150_73), .B (n_149_79), .C1 (n_149_83), .C2 (n_150_89) );
AOI211_X1 g_149_67 (.ZN (n_149_67), .A (n_149_71), .B (n_150_77), .C1 (n_150_81), .C2 (n_149_87) );
AOI211_X1 g_150_65 (.ZN (n_150_65), .A (n_150_69), .B (n_149_75), .C1 (n_149_79), .C2 (n_150_85) );
AOI211_X1 g_149_63 (.ZN (n_149_63), .A (n_149_67), .B (n_150_73), .C1 (n_150_77), .C2 (n_149_83) );
AOI211_X1 g_150_61 (.ZN (n_150_61), .A (n_150_65), .B (n_149_71), .C1 (n_149_75), .C2 (n_150_81) );
AOI211_X1 g_149_59 (.ZN (n_149_59), .A (n_149_63), .B (n_150_69), .C1 (n_150_73), .C2 (n_149_79) );
AOI211_X1 g_150_57 (.ZN (n_150_57), .A (n_150_61), .B (n_149_67), .C1 (n_149_71), .C2 (n_150_77) );
AOI211_X1 g_149_55 (.ZN (n_149_55), .A (n_149_59), .B (n_150_65), .C1 (n_150_69), .C2 (n_149_75) );
AOI211_X1 g_150_53 (.ZN (n_150_53), .A (n_150_57), .B (n_149_63), .C1 (n_149_67), .C2 (n_150_73) );
AOI211_X1 g_149_51 (.ZN (n_149_51), .A (n_149_55), .B (n_150_61), .C1 (n_150_65), .C2 (n_149_71) );
AOI211_X1 g_150_49 (.ZN (n_150_49), .A (n_150_53), .B (n_149_59), .C1 (n_149_63), .C2 (n_150_69) );
AOI211_X1 g_149_47 (.ZN (n_149_47), .A (n_149_51), .B (n_150_57), .C1 (n_150_61), .C2 (n_149_67) );
AOI211_X1 g_150_45 (.ZN (n_150_45), .A (n_150_49), .B (n_149_55), .C1 (n_149_59), .C2 (n_150_65) );
AOI211_X1 g_149_43 (.ZN (n_149_43), .A (n_149_47), .B (n_150_53), .C1 (n_150_57), .C2 (n_149_63) );
AOI211_X1 g_150_41 (.ZN (n_150_41), .A (n_150_45), .B (n_149_51), .C1 (n_149_55), .C2 (n_150_61) );
AOI211_X1 g_149_39 (.ZN (n_149_39), .A (n_149_43), .B (n_150_49), .C1 (n_150_53), .C2 (n_149_59) );
AOI211_X1 g_150_37 (.ZN (n_150_37), .A (n_150_41), .B (n_149_47), .C1 (n_149_51), .C2 (n_150_57) );
AOI211_X1 g_149_35 (.ZN (n_149_35), .A (n_149_39), .B (n_150_45), .C1 (n_150_49), .C2 (n_149_55) );
AOI211_X1 g_150_33 (.ZN (n_150_33), .A (n_150_37), .B (n_149_43), .C1 (n_149_47), .C2 (n_150_53) );
AOI211_X1 g_149_31 (.ZN (n_149_31), .A (n_149_35), .B (n_150_41), .C1 (n_150_45), .C2 (n_149_51) );
AOI211_X1 g_150_29 (.ZN (n_150_29), .A (n_150_33), .B (n_149_39), .C1 (n_149_43), .C2 (n_150_49) );
AOI211_X1 g_149_27 (.ZN (n_149_27), .A (n_149_31), .B (n_150_37), .C1 (n_150_41), .C2 (n_149_47) );
AOI211_X1 g_150_25 (.ZN (n_150_25), .A (n_150_29), .B (n_149_35), .C1 (n_149_39), .C2 (n_150_45) );
AOI211_X1 g_149_23 (.ZN (n_149_23), .A (n_149_27), .B (n_150_33), .C1 (n_150_37), .C2 (n_149_43) );
AOI211_X1 g_150_21 (.ZN (n_150_21), .A (n_150_25), .B (n_149_31), .C1 (n_149_35), .C2 (n_150_41) );
AOI211_X1 g_149_19 (.ZN (n_149_19), .A (n_149_23), .B (n_150_29), .C1 (n_150_33), .C2 (n_149_39) );
AOI211_X1 g_150_17 (.ZN (n_150_17), .A (n_150_21), .B (n_149_27), .C1 (n_149_31), .C2 (n_150_37) );
AOI211_X1 g_149_15 (.ZN (n_149_15), .A (n_149_19), .B (n_150_25), .C1 (n_150_29), .C2 (n_149_35) );
AOI211_X1 g_150_13 (.ZN (n_150_13), .A (n_150_17), .B (n_149_23), .C1 (n_149_27), .C2 (n_150_33) );
AOI211_X1 g_149_11 (.ZN (n_149_11), .A (n_149_15), .B (n_150_21), .C1 (n_150_25), .C2 (n_149_31) );
AOI211_X1 g_150_9 (.ZN (n_150_9), .A (n_150_13), .B (n_149_19), .C1 (n_149_23), .C2 (n_150_29) );
AOI211_X1 g_149_7 (.ZN (n_149_7), .A (n_149_11), .B (n_150_17), .C1 (n_150_21), .C2 (n_149_27) );
AOI211_X1 g_148_5 (.ZN (n_148_5), .A (n_150_9), .B (n_149_15), .C1 (n_149_19), .C2 (n_150_25) );
AOI211_X1 g_146_4 (.ZN (n_146_4), .A (n_149_7), .B (n_150_13), .C1 (n_150_17), .C2 (n_149_23) );
AOI211_X1 g_148_3 (.ZN (n_148_3), .A (n_148_5), .B (n_149_11), .C1 (n_149_15), .C2 (n_150_21) );
AOI211_X1 g_146_2 (.ZN (n_146_2), .A (n_146_4), .B (n_150_9), .C1 (n_150_13), .C2 (n_149_19) );
AOI211_X1 g_144_1 (.ZN (n_144_1), .A (n_148_3), .B (n_149_7), .C1 (n_149_11), .C2 (n_150_17) );
AOI211_X1 g_143_3 (.ZN (n_143_3), .A (n_146_2), .B (n_148_5), .C1 (n_150_9), .C2 (n_149_15) );
AOI211_X1 g_145_4 (.ZN (n_145_4), .A (n_144_1), .B (n_146_4), .C1 (n_149_7), .C2 (n_150_13) );
AOI211_X1 g_147_5 (.ZN (n_147_5), .A (n_143_3), .B (n_148_3), .C1 (n_148_5), .C2 (n_149_11) );
AOI211_X1 g_148_7 (.ZN (n_148_7), .A (n_145_4), .B (n_146_2), .C1 (n_146_4), .C2 (n_150_9) );
AOI211_X1 g_149_5 (.ZN (n_149_5), .A (n_147_5), .B (n_144_1), .C1 (n_148_3), .C2 (n_149_7) );
AOI211_X1 g_150_7 (.ZN (n_150_7), .A (n_148_7), .B (n_143_3), .C1 (n_146_2), .C2 (n_148_5) );
AOI211_X1 g_148_6 (.ZN (n_148_6), .A (n_149_5), .B (n_145_4), .C1 (n_144_1), .C2 (n_146_4) );
AOI211_X1 g_147_4 (.ZN (n_147_4), .A (n_150_7), .B (n_147_5), .C1 (n_143_3), .C2 (n_148_3) );
AOI211_X1 g_145_3 (.ZN (n_145_3), .A (n_148_6), .B (n_148_7), .C1 (n_145_4), .C2 (n_146_2) );
AOI211_X1 g_143_2 (.ZN (n_143_2), .A (n_147_4), .B (n_149_5), .C1 (n_147_5), .C2 (n_144_1) );
AOI211_X1 g_141_1 (.ZN (n_141_1), .A (n_145_3), .B (n_150_7), .C1 (n_148_7), .C2 (n_143_3) );
AOI211_X1 g_142_3 (.ZN (n_142_3), .A (n_143_2), .B (n_148_6), .C1 (n_149_5), .C2 (n_145_4) );
AOI211_X1 g_144_4 (.ZN (n_144_4), .A (n_141_1), .B (n_147_4), .C1 (n_150_7), .C2 (n_147_5) );
AOI211_X1 g_146_5 (.ZN (n_146_5), .A (n_142_3), .B (n_145_3), .C1 (n_148_6), .C2 (n_148_7) );
AOI211_X1 g_147_7 (.ZN (n_147_7), .A (n_144_4), .B (n_143_2), .C1 (n_147_4), .C2 (n_149_5) );
AOI211_X1 g_148_9 (.ZN (n_148_9), .A (n_146_5), .B (n_141_1), .C1 (n_145_3), .C2 (n_150_7) );
AOI211_X1 g_147_11 (.ZN (n_147_11), .A (n_147_7), .B (n_142_3), .C1 (n_143_2), .C2 (n_148_6) );
AOI211_X1 g_148_13 (.ZN (n_148_13), .A (n_148_9), .B (n_144_4), .C1 (n_141_1), .C2 (n_147_4) );
AOI211_X1 g_147_15 (.ZN (n_147_15), .A (n_147_11), .B (n_146_5), .C1 (n_142_3), .C2 (n_145_3) );
AOI211_X1 g_148_17 (.ZN (n_148_17), .A (n_148_13), .B (n_147_7), .C1 (n_144_4), .C2 (n_143_2) );
AOI211_X1 g_147_19 (.ZN (n_147_19), .A (n_147_15), .B (n_148_9), .C1 (n_146_5), .C2 (n_141_1) );
AOI211_X1 g_148_21 (.ZN (n_148_21), .A (n_148_17), .B (n_147_11), .C1 (n_147_7), .C2 (n_142_3) );
AOI211_X1 g_147_23 (.ZN (n_147_23), .A (n_147_19), .B (n_148_13), .C1 (n_148_9), .C2 (n_144_4) );
AOI211_X1 g_148_25 (.ZN (n_148_25), .A (n_148_21), .B (n_147_15), .C1 (n_147_11), .C2 (n_146_5) );
AOI211_X1 g_147_27 (.ZN (n_147_27), .A (n_147_23), .B (n_148_17), .C1 (n_148_13), .C2 (n_147_7) );
AOI211_X1 g_148_29 (.ZN (n_148_29), .A (n_148_25), .B (n_147_19), .C1 (n_147_15), .C2 (n_148_9) );
AOI211_X1 g_147_31 (.ZN (n_147_31), .A (n_147_27), .B (n_148_21), .C1 (n_148_17), .C2 (n_147_11) );
AOI211_X1 g_148_33 (.ZN (n_148_33), .A (n_148_29), .B (n_147_23), .C1 (n_147_19), .C2 (n_148_13) );
AOI211_X1 g_147_35 (.ZN (n_147_35), .A (n_147_31), .B (n_148_25), .C1 (n_148_21), .C2 (n_147_15) );
AOI211_X1 g_148_37 (.ZN (n_148_37), .A (n_148_33), .B (n_147_27), .C1 (n_147_23), .C2 (n_148_17) );
AOI211_X1 g_147_39 (.ZN (n_147_39), .A (n_147_35), .B (n_148_29), .C1 (n_148_25), .C2 (n_147_19) );
AOI211_X1 g_148_41 (.ZN (n_148_41), .A (n_148_37), .B (n_147_31), .C1 (n_147_27), .C2 (n_148_21) );
AOI211_X1 g_147_43 (.ZN (n_147_43), .A (n_147_39), .B (n_148_33), .C1 (n_148_29), .C2 (n_147_23) );
AOI211_X1 g_148_45 (.ZN (n_148_45), .A (n_148_41), .B (n_147_35), .C1 (n_147_31), .C2 (n_148_25) );
AOI211_X1 g_147_47 (.ZN (n_147_47), .A (n_147_43), .B (n_148_37), .C1 (n_148_33), .C2 (n_147_27) );
AOI211_X1 g_148_49 (.ZN (n_148_49), .A (n_148_45), .B (n_147_39), .C1 (n_147_35), .C2 (n_148_29) );
AOI211_X1 g_147_51 (.ZN (n_147_51), .A (n_147_47), .B (n_148_41), .C1 (n_148_37), .C2 (n_147_31) );
AOI211_X1 g_148_53 (.ZN (n_148_53), .A (n_148_49), .B (n_147_43), .C1 (n_147_39), .C2 (n_148_33) );
AOI211_X1 g_147_55 (.ZN (n_147_55), .A (n_147_51), .B (n_148_45), .C1 (n_148_41), .C2 (n_147_35) );
AOI211_X1 g_148_57 (.ZN (n_148_57), .A (n_148_53), .B (n_147_47), .C1 (n_147_43), .C2 (n_148_37) );
AOI211_X1 g_147_59 (.ZN (n_147_59), .A (n_147_55), .B (n_148_49), .C1 (n_148_45), .C2 (n_147_39) );
AOI211_X1 g_148_61 (.ZN (n_148_61), .A (n_148_57), .B (n_147_51), .C1 (n_147_47), .C2 (n_148_41) );
AOI211_X1 g_147_63 (.ZN (n_147_63), .A (n_147_59), .B (n_148_53), .C1 (n_148_49), .C2 (n_147_43) );
AOI211_X1 g_148_65 (.ZN (n_148_65), .A (n_148_61), .B (n_147_55), .C1 (n_147_51), .C2 (n_148_45) );
AOI211_X1 g_147_67 (.ZN (n_147_67), .A (n_147_63), .B (n_148_57), .C1 (n_148_53), .C2 (n_147_47) );
AOI211_X1 g_148_69 (.ZN (n_148_69), .A (n_148_65), .B (n_147_59), .C1 (n_147_55), .C2 (n_148_49) );
AOI211_X1 g_147_71 (.ZN (n_147_71), .A (n_147_67), .B (n_148_61), .C1 (n_148_57), .C2 (n_147_51) );
AOI211_X1 g_148_73 (.ZN (n_148_73), .A (n_148_69), .B (n_147_63), .C1 (n_147_59), .C2 (n_148_53) );
AOI211_X1 g_147_75 (.ZN (n_147_75), .A (n_147_71), .B (n_148_65), .C1 (n_148_61), .C2 (n_147_55) );
AOI211_X1 g_148_77 (.ZN (n_148_77), .A (n_148_73), .B (n_147_67), .C1 (n_147_63), .C2 (n_148_57) );
AOI211_X1 g_147_79 (.ZN (n_147_79), .A (n_147_75), .B (n_148_69), .C1 (n_148_65), .C2 (n_147_59) );
AOI211_X1 g_148_81 (.ZN (n_148_81), .A (n_148_77), .B (n_147_71), .C1 (n_147_67), .C2 (n_148_61) );
AOI211_X1 g_147_83 (.ZN (n_147_83), .A (n_147_79), .B (n_148_73), .C1 (n_148_69), .C2 (n_147_63) );
AOI211_X1 g_148_85 (.ZN (n_148_85), .A (n_148_81), .B (n_147_75), .C1 (n_147_71), .C2 (n_148_65) );
AOI211_X1 g_147_87 (.ZN (n_147_87), .A (n_147_83), .B (n_148_77), .C1 (n_148_73), .C2 (n_147_67) );
AOI211_X1 g_148_89 (.ZN (n_148_89), .A (n_148_85), .B (n_147_79), .C1 (n_147_75), .C2 (n_148_69) );
AOI211_X1 g_147_91 (.ZN (n_147_91), .A (n_147_87), .B (n_148_81), .C1 (n_148_77), .C2 (n_147_71) );
AOI211_X1 g_148_93 (.ZN (n_148_93), .A (n_148_89), .B (n_147_83), .C1 (n_147_79), .C2 (n_148_73) );
AOI211_X1 g_147_95 (.ZN (n_147_95), .A (n_147_91), .B (n_148_85), .C1 (n_148_81), .C2 (n_147_75) );
AOI211_X1 g_148_97 (.ZN (n_148_97), .A (n_148_93), .B (n_147_87), .C1 (n_147_83), .C2 (n_148_77) );
AOI211_X1 g_147_99 (.ZN (n_147_99), .A (n_147_95), .B (n_148_89), .C1 (n_148_85), .C2 (n_147_79) );
AOI211_X1 g_148_101 (.ZN (n_148_101), .A (n_148_97), .B (n_147_91), .C1 (n_147_87), .C2 (n_148_81) );
AOI211_X1 g_147_103 (.ZN (n_147_103), .A (n_147_99), .B (n_148_93), .C1 (n_148_89), .C2 (n_147_83) );
AOI211_X1 g_148_105 (.ZN (n_148_105), .A (n_148_101), .B (n_147_95), .C1 (n_147_91), .C2 (n_148_85) );
AOI211_X1 g_147_107 (.ZN (n_147_107), .A (n_147_103), .B (n_148_97), .C1 (n_148_93), .C2 (n_147_87) );
AOI211_X1 g_148_109 (.ZN (n_148_109), .A (n_148_105), .B (n_147_99), .C1 (n_147_95), .C2 (n_148_89) );
AOI211_X1 g_147_111 (.ZN (n_147_111), .A (n_147_107), .B (n_148_101), .C1 (n_148_97), .C2 (n_147_91) );
AOI211_X1 g_148_113 (.ZN (n_148_113), .A (n_148_109), .B (n_147_103), .C1 (n_147_99), .C2 (n_148_93) );
AOI211_X1 g_147_115 (.ZN (n_147_115), .A (n_147_111), .B (n_148_105), .C1 (n_148_101), .C2 (n_147_95) );
AOI211_X1 g_148_117 (.ZN (n_148_117), .A (n_148_113), .B (n_147_107), .C1 (n_147_103), .C2 (n_148_97) );
AOI211_X1 g_147_119 (.ZN (n_147_119), .A (n_147_115), .B (n_148_109), .C1 (n_148_105), .C2 (n_147_99) );
AOI211_X1 g_148_121 (.ZN (n_148_121), .A (n_148_117), .B (n_147_111), .C1 (n_147_107), .C2 (n_148_101) );
AOI211_X1 g_147_123 (.ZN (n_147_123), .A (n_147_119), .B (n_148_113), .C1 (n_148_109), .C2 (n_147_103) );
AOI211_X1 g_148_125 (.ZN (n_148_125), .A (n_148_121), .B (n_147_115), .C1 (n_147_111), .C2 (n_148_105) );
AOI211_X1 g_147_127 (.ZN (n_147_127), .A (n_147_123), .B (n_148_117), .C1 (n_148_113), .C2 (n_147_107) );
AOI211_X1 g_148_129 (.ZN (n_148_129), .A (n_148_125), .B (n_147_119), .C1 (n_147_115), .C2 (n_148_109) );
AOI211_X1 g_147_131 (.ZN (n_147_131), .A (n_147_127), .B (n_148_121), .C1 (n_148_117), .C2 (n_147_111) );
AOI211_X1 g_148_133 (.ZN (n_148_133), .A (n_148_129), .B (n_147_123), .C1 (n_147_119), .C2 (n_148_113) );
AOI211_X1 g_147_135 (.ZN (n_147_135), .A (n_147_131), .B (n_148_125), .C1 (n_148_121), .C2 (n_147_115) );
AOI211_X1 g_148_137 (.ZN (n_148_137), .A (n_148_133), .B (n_147_127), .C1 (n_147_123), .C2 (n_148_117) );
AOI211_X1 g_147_139 (.ZN (n_147_139), .A (n_147_135), .B (n_148_129), .C1 (n_148_125), .C2 (n_147_119) );
AOI211_X1 g_146_137 (.ZN (n_146_137), .A (n_148_137), .B (n_147_131), .C1 (n_147_127), .C2 (n_148_121) );
AOI211_X1 g_148_136 (.ZN (n_148_136), .A (n_147_139), .B (n_148_133), .C1 (n_148_129), .C2 (n_147_123) );
AOI211_X1 g_150_135 (.ZN (n_150_135), .A (n_146_137), .B (n_147_135), .C1 (n_147_131), .C2 (n_148_125) );
AOI211_X1 g_148_134 (.ZN (n_148_134), .A (n_148_136), .B (n_148_137), .C1 (n_148_133), .C2 (n_147_127) );
AOI211_X1 g_146_133 (.ZN (n_146_133), .A (n_150_135), .B (n_147_139), .C1 (n_147_135), .C2 (n_148_129) );
AOI211_X1 g_148_132 (.ZN (n_148_132), .A (n_148_134), .B (n_146_137), .C1 (n_148_137), .C2 (n_147_131) );
AOI211_X1 g_150_131 (.ZN (n_150_131), .A (n_146_133), .B (n_148_136), .C1 (n_147_139), .C2 (n_148_133) );
AOI211_X1 g_148_130 (.ZN (n_148_130), .A (n_148_132), .B (n_150_135), .C1 (n_146_137), .C2 (n_147_135) );
AOI211_X1 g_146_129 (.ZN (n_146_129), .A (n_150_131), .B (n_148_134), .C1 (n_148_136), .C2 (n_148_137) );
AOI211_X1 g_148_128 (.ZN (n_148_128), .A (n_148_130), .B (n_146_133), .C1 (n_150_135), .C2 (n_147_139) );
AOI211_X1 g_150_127 (.ZN (n_150_127), .A (n_146_129), .B (n_148_132), .C1 (n_148_134), .C2 (n_146_137) );
AOI211_X1 g_148_126 (.ZN (n_148_126), .A (n_148_128), .B (n_150_131), .C1 (n_146_133), .C2 (n_148_136) );
AOI211_X1 g_146_125 (.ZN (n_146_125), .A (n_150_127), .B (n_148_130), .C1 (n_148_132), .C2 (n_150_135) );
AOI211_X1 g_148_124 (.ZN (n_148_124), .A (n_148_126), .B (n_146_129), .C1 (n_150_131), .C2 (n_148_134) );
AOI211_X1 g_150_123 (.ZN (n_150_123), .A (n_146_125), .B (n_148_128), .C1 (n_148_130), .C2 (n_146_133) );
AOI211_X1 g_148_122 (.ZN (n_148_122), .A (n_148_124), .B (n_150_127), .C1 (n_146_129), .C2 (n_148_132) );
AOI211_X1 g_146_121 (.ZN (n_146_121), .A (n_150_123), .B (n_148_126), .C1 (n_148_128), .C2 (n_150_131) );
AOI211_X1 g_148_120 (.ZN (n_148_120), .A (n_148_122), .B (n_146_125), .C1 (n_150_127), .C2 (n_148_130) );
AOI211_X1 g_150_119 (.ZN (n_150_119), .A (n_146_121), .B (n_148_124), .C1 (n_148_126), .C2 (n_146_129) );
AOI211_X1 g_148_118 (.ZN (n_148_118), .A (n_148_120), .B (n_150_123), .C1 (n_146_125), .C2 (n_148_128) );
AOI211_X1 g_146_117 (.ZN (n_146_117), .A (n_150_119), .B (n_148_122), .C1 (n_148_124), .C2 (n_150_127) );
AOI211_X1 g_148_116 (.ZN (n_148_116), .A (n_148_118), .B (n_146_121), .C1 (n_150_123), .C2 (n_148_126) );
AOI211_X1 g_150_115 (.ZN (n_150_115), .A (n_146_117), .B (n_148_120), .C1 (n_148_122), .C2 (n_146_125) );
AOI211_X1 g_148_114 (.ZN (n_148_114), .A (n_148_116), .B (n_150_119), .C1 (n_146_121), .C2 (n_148_124) );
AOI211_X1 g_146_113 (.ZN (n_146_113), .A (n_150_115), .B (n_148_118), .C1 (n_148_120), .C2 (n_150_123) );
AOI211_X1 g_148_112 (.ZN (n_148_112), .A (n_148_114), .B (n_146_117), .C1 (n_150_119), .C2 (n_148_122) );
AOI211_X1 g_150_111 (.ZN (n_150_111), .A (n_146_113), .B (n_148_116), .C1 (n_148_118), .C2 (n_146_121) );
AOI211_X1 g_148_110 (.ZN (n_148_110), .A (n_148_112), .B (n_150_115), .C1 (n_146_117), .C2 (n_148_120) );
AOI211_X1 g_146_109 (.ZN (n_146_109), .A (n_150_111), .B (n_148_114), .C1 (n_148_116), .C2 (n_150_119) );
AOI211_X1 g_148_108 (.ZN (n_148_108), .A (n_148_110), .B (n_146_113), .C1 (n_150_115), .C2 (n_148_118) );
AOI211_X1 g_150_107 (.ZN (n_150_107), .A (n_146_109), .B (n_148_112), .C1 (n_148_114), .C2 (n_146_117) );
AOI211_X1 g_148_106 (.ZN (n_148_106), .A (n_148_108), .B (n_150_111), .C1 (n_146_113), .C2 (n_148_116) );
AOI211_X1 g_146_105 (.ZN (n_146_105), .A (n_150_107), .B (n_148_110), .C1 (n_148_112), .C2 (n_150_115) );
AOI211_X1 g_148_104 (.ZN (n_148_104), .A (n_148_106), .B (n_146_109), .C1 (n_150_111), .C2 (n_148_114) );
AOI211_X1 g_150_103 (.ZN (n_150_103), .A (n_146_105), .B (n_148_108), .C1 (n_148_110), .C2 (n_146_113) );
AOI211_X1 g_148_102 (.ZN (n_148_102), .A (n_148_104), .B (n_150_107), .C1 (n_146_109), .C2 (n_148_112) );
AOI211_X1 g_146_101 (.ZN (n_146_101), .A (n_150_103), .B (n_148_106), .C1 (n_148_108), .C2 (n_150_111) );
AOI211_X1 g_148_100 (.ZN (n_148_100), .A (n_148_102), .B (n_146_105), .C1 (n_150_107), .C2 (n_148_110) );
AOI211_X1 g_150_99 (.ZN (n_150_99), .A (n_146_101), .B (n_148_104), .C1 (n_148_106), .C2 (n_146_109) );
AOI211_X1 g_148_98 (.ZN (n_148_98), .A (n_148_100), .B (n_150_103), .C1 (n_146_105), .C2 (n_148_108) );
AOI211_X1 g_146_97 (.ZN (n_146_97), .A (n_150_99), .B (n_148_102), .C1 (n_148_104), .C2 (n_150_107) );
AOI211_X1 g_148_96 (.ZN (n_148_96), .A (n_148_98), .B (n_146_101), .C1 (n_150_103), .C2 (n_148_106) );
AOI211_X1 g_150_95 (.ZN (n_150_95), .A (n_146_97), .B (n_148_100), .C1 (n_148_102), .C2 (n_146_105) );
AOI211_X1 g_148_94 (.ZN (n_148_94), .A (n_148_96), .B (n_150_99), .C1 (n_146_101), .C2 (n_148_104) );
AOI211_X1 g_146_93 (.ZN (n_146_93), .A (n_150_95), .B (n_148_98), .C1 (n_148_100), .C2 (n_150_103) );
AOI211_X1 g_148_92 (.ZN (n_148_92), .A (n_148_94), .B (n_146_97), .C1 (n_150_99), .C2 (n_148_102) );
AOI211_X1 g_150_91 (.ZN (n_150_91), .A (n_146_93), .B (n_148_96), .C1 (n_148_98), .C2 (n_146_101) );
AOI211_X1 g_148_90 (.ZN (n_148_90), .A (n_148_92), .B (n_150_95), .C1 (n_146_97), .C2 (n_148_100) );
AOI211_X1 g_146_89 (.ZN (n_146_89), .A (n_150_91), .B (n_148_94), .C1 (n_148_96), .C2 (n_150_99) );
AOI211_X1 g_148_88 (.ZN (n_148_88), .A (n_148_90), .B (n_146_93), .C1 (n_150_95), .C2 (n_148_98) );
AOI211_X1 g_150_87 (.ZN (n_150_87), .A (n_146_89), .B (n_148_92), .C1 (n_148_94), .C2 (n_146_97) );
AOI211_X1 g_148_86 (.ZN (n_148_86), .A (n_148_88), .B (n_150_91), .C1 (n_146_93), .C2 (n_148_96) );
AOI211_X1 g_146_85 (.ZN (n_146_85), .A (n_150_87), .B (n_148_90), .C1 (n_148_92), .C2 (n_150_95) );
AOI211_X1 g_148_84 (.ZN (n_148_84), .A (n_148_86), .B (n_146_89), .C1 (n_150_91), .C2 (n_148_94) );
AOI211_X1 g_150_83 (.ZN (n_150_83), .A (n_146_85), .B (n_148_88), .C1 (n_148_90), .C2 (n_146_93) );
AOI211_X1 g_148_82 (.ZN (n_148_82), .A (n_148_84), .B (n_150_87), .C1 (n_146_89), .C2 (n_148_92) );
AOI211_X1 g_146_81 (.ZN (n_146_81), .A (n_150_83), .B (n_148_86), .C1 (n_148_88), .C2 (n_150_91) );
AOI211_X1 g_148_80 (.ZN (n_148_80), .A (n_148_82), .B (n_146_85), .C1 (n_150_87), .C2 (n_148_90) );
AOI211_X1 g_150_79 (.ZN (n_150_79), .A (n_146_81), .B (n_148_84), .C1 (n_148_86), .C2 (n_146_89) );
AOI211_X1 g_148_78 (.ZN (n_148_78), .A (n_148_80), .B (n_150_83), .C1 (n_146_85), .C2 (n_148_88) );
AOI211_X1 g_146_77 (.ZN (n_146_77), .A (n_150_79), .B (n_148_82), .C1 (n_148_84), .C2 (n_150_87) );
AOI211_X1 g_148_76 (.ZN (n_148_76), .A (n_148_78), .B (n_146_81), .C1 (n_150_83), .C2 (n_148_86) );
AOI211_X1 g_150_75 (.ZN (n_150_75), .A (n_146_77), .B (n_148_80), .C1 (n_148_82), .C2 (n_146_85) );
AOI211_X1 g_148_74 (.ZN (n_148_74), .A (n_148_76), .B (n_150_79), .C1 (n_146_81), .C2 (n_148_84) );
AOI211_X1 g_146_73 (.ZN (n_146_73), .A (n_150_75), .B (n_148_78), .C1 (n_148_80), .C2 (n_150_83) );
AOI211_X1 g_148_72 (.ZN (n_148_72), .A (n_148_74), .B (n_146_77), .C1 (n_150_79), .C2 (n_148_82) );
AOI211_X1 g_150_71 (.ZN (n_150_71), .A (n_146_73), .B (n_148_76), .C1 (n_148_78), .C2 (n_146_81) );
AOI211_X1 g_148_70 (.ZN (n_148_70), .A (n_148_72), .B (n_150_75), .C1 (n_146_77), .C2 (n_148_80) );
AOI211_X1 g_146_69 (.ZN (n_146_69), .A (n_150_71), .B (n_148_74), .C1 (n_148_76), .C2 (n_150_79) );
AOI211_X1 g_148_68 (.ZN (n_148_68), .A (n_148_70), .B (n_146_73), .C1 (n_150_75), .C2 (n_148_78) );
AOI211_X1 g_150_67 (.ZN (n_150_67), .A (n_146_69), .B (n_148_72), .C1 (n_148_74), .C2 (n_146_77) );
AOI211_X1 g_148_66 (.ZN (n_148_66), .A (n_148_68), .B (n_150_71), .C1 (n_146_73), .C2 (n_148_76) );
AOI211_X1 g_146_65 (.ZN (n_146_65), .A (n_150_67), .B (n_148_70), .C1 (n_148_72), .C2 (n_150_75) );
AOI211_X1 g_148_64 (.ZN (n_148_64), .A (n_148_66), .B (n_146_69), .C1 (n_150_71), .C2 (n_148_74) );
AOI211_X1 g_150_63 (.ZN (n_150_63), .A (n_146_65), .B (n_148_68), .C1 (n_148_70), .C2 (n_146_73) );
AOI211_X1 g_148_62 (.ZN (n_148_62), .A (n_148_64), .B (n_150_67), .C1 (n_146_69), .C2 (n_148_72) );
AOI211_X1 g_146_61 (.ZN (n_146_61), .A (n_150_63), .B (n_148_66), .C1 (n_148_68), .C2 (n_150_71) );
AOI211_X1 g_148_60 (.ZN (n_148_60), .A (n_148_62), .B (n_146_65), .C1 (n_150_67), .C2 (n_148_70) );
AOI211_X1 g_150_59 (.ZN (n_150_59), .A (n_146_61), .B (n_148_64), .C1 (n_148_66), .C2 (n_146_69) );
AOI211_X1 g_148_58 (.ZN (n_148_58), .A (n_148_60), .B (n_150_63), .C1 (n_146_65), .C2 (n_148_68) );
AOI211_X1 g_146_57 (.ZN (n_146_57), .A (n_150_59), .B (n_148_62), .C1 (n_148_64), .C2 (n_150_67) );
AOI211_X1 g_148_56 (.ZN (n_148_56), .A (n_148_58), .B (n_146_61), .C1 (n_150_63), .C2 (n_148_66) );
AOI211_X1 g_150_55 (.ZN (n_150_55), .A (n_146_57), .B (n_148_60), .C1 (n_148_62), .C2 (n_146_65) );
AOI211_X1 g_148_54 (.ZN (n_148_54), .A (n_148_56), .B (n_150_59), .C1 (n_146_61), .C2 (n_148_64) );
AOI211_X1 g_146_53 (.ZN (n_146_53), .A (n_150_55), .B (n_148_58), .C1 (n_148_60), .C2 (n_150_63) );
AOI211_X1 g_148_52 (.ZN (n_148_52), .A (n_148_54), .B (n_146_57), .C1 (n_150_59), .C2 (n_148_62) );
AOI211_X1 g_150_51 (.ZN (n_150_51), .A (n_146_53), .B (n_148_56), .C1 (n_148_58), .C2 (n_146_61) );
AOI211_X1 g_148_50 (.ZN (n_148_50), .A (n_148_52), .B (n_150_55), .C1 (n_146_57), .C2 (n_148_60) );
AOI211_X1 g_146_49 (.ZN (n_146_49), .A (n_150_51), .B (n_148_54), .C1 (n_148_56), .C2 (n_150_59) );
AOI211_X1 g_148_48 (.ZN (n_148_48), .A (n_148_50), .B (n_146_53), .C1 (n_150_55), .C2 (n_148_58) );
AOI211_X1 g_150_47 (.ZN (n_150_47), .A (n_146_49), .B (n_148_52), .C1 (n_148_54), .C2 (n_146_57) );
AOI211_X1 g_148_46 (.ZN (n_148_46), .A (n_148_48), .B (n_150_51), .C1 (n_146_53), .C2 (n_148_56) );
AOI211_X1 g_146_45 (.ZN (n_146_45), .A (n_150_47), .B (n_148_50), .C1 (n_148_52), .C2 (n_150_55) );
AOI211_X1 g_148_44 (.ZN (n_148_44), .A (n_148_46), .B (n_146_49), .C1 (n_150_51), .C2 (n_148_54) );
AOI211_X1 g_150_43 (.ZN (n_150_43), .A (n_146_45), .B (n_148_48), .C1 (n_148_50), .C2 (n_146_53) );
AOI211_X1 g_148_42 (.ZN (n_148_42), .A (n_148_44), .B (n_150_47), .C1 (n_146_49), .C2 (n_148_52) );
AOI211_X1 g_146_41 (.ZN (n_146_41), .A (n_150_43), .B (n_148_46), .C1 (n_148_48), .C2 (n_150_51) );
AOI211_X1 g_148_40 (.ZN (n_148_40), .A (n_148_42), .B (n_146_45), .C1 (n_150_47), .C2 (n_148_50) );
AOI211_X1 g_150_39 (.ZN (n_150_39), .A (n_146_41), .B (n_148_44), .C1 (n_148_46), .C2 (n_146_49) );
AOI211_X1 g_148_38 (.ZN (n_148_38), .A (n_148_40), .B (n_150_43), .C1 (n_146_45), .C2 (n_148_48) );
AOI211_X1 g_146_37 (.ZN (n_146_37), .A (n_150_39), .B (n_148_42), .C1 (n_148_44), .C2 (n_150_47) );
AOI211_X1 g_148_36 (.ZN (n_148_36), .A (n_148_38), .B (n_146_41), .C1 (n_150_43), .C2 (n_148_46) );
AOI211_X1 g_150_35 (.ZN (n_150_35), .A (n_146_37), .B (n_148_40), .C1 (n_148_42), .C2 (n_146_45) );
AOI211_X1 g_148_34 (.ZN (n_148_34), .A (n_148_36), .B (n_150_39), .C1 (n_146_41), .C2 (n_148_44) );
AOI211_X1 g_146_33 (.ZN (n_146_33), .A (n_150_35), .B (n_148_38), .C1 (n_148_40), .C2 (n_150_43) );
AOI211_X1 g_148_32 (.ZN (n_148_32), .A (n_148_34), .B (n_146_37), .C1 (n_150_39), .C2 (n_148_42) );
AOI211_X1 g_150_31 (.ZN (n_150_31), .A (n_146_33), .B (n_148_36), .C1 (n_148_38), .C2 (n_146_41) );
AOI211_X1 g_148_30 (.ZN (n_148_30), .A (n_148_32), .B (n_150_35), .C1 (n_146_37), .C2 (n_148_40) );
AOI211_X1 g_146_29 (.ZN (n_146_29), .A (n_150_31), .B (n_148_34), .C1 (n_148_36), .C2 (n_150_39) );
AOI211_X1 g_148_28 (.ZN (n_148_28), .A (n_148_30), .B (n_146_33), .C1 (n_150_35), .C2 (n_148_38) );
AOI211_X1 g_150_27 (.ZN (n_150_27), .A (n_146_29), .B (n_148_32), .C1 (n_148_34), .C2 (n_146_37) );
AOI211_X1 g_148_26 (.ZN (n_148_26), .A (n_148_28), .B (n_150_31), .C1 (n_146_33), .C2 (n_148_36) );
AOI211_X1 g_146_25 (.ZN (n_146_25), .A (n_150_27), .B (n_148_30), .C1 (n_148_32), .C2 (n_150_35) );
AOI211_X1 g_148_24 (.ZN (n_148_24), .A (n_148_26), .B (n_146_29), .C1 (n_150_31), .C2 (n_148_34) );
AOI211_X1 g_150_23 (.ZN (n_150_23), .A (n_146_25), .B (n_148_28), .C1 (n_148_30), .C2 (n_146_33) );
AOI211_X1 g_148_22 (.ZN (n_148_22), .A (n_148_24), .B (n_150_27), .C1 (n_146_29), .C2 (n_148_32) );
AOI211_X1 g_146_21 (.ZN (n_146_21), .A (n_150_23), .B (n_148_26), .C1 (n_148_28), .C2 (n_150_31) );
AOI211_X1 g_148_20 (.ZN (n_148_20), .A (n_148_22), .B (n_146_25), .C1 (n_150_27), .C2 (n_148_30) );
AOI211_X1 g_150_19 (.ZN (n_150_19), .A (n_146_21), .B (n_148_24), .C1 (n_148_26), .C2 (n_146_29) );
AOI211_X1 g_148_18 (.ZN (n_148_18), .A (n_148_20), .B (n_150_23), .C1 (n_146_25), .C2 (n_148_28) );
AOI211_X1 g_146_17 (.ZN (n_146_17), .A (n_150_19), .B (n_148_22), .C1 (n_148_24), .C2 (n_150_27) );
AOI211_X1 g_148_16 (.ZN (n_148_16), .A (n_148_18), .B (n_146_21), .C1 (n_150_23), .C2 (n_148_26) );
AOI211_X1 g_150_15 (.ZN (n_150_15), .A (n_146_17), .B (n_148_20), .C1 (n_148_22), .C2 (n_146_25) );
AOI211_X1 g_148_14 (.ZN (n_148_14), .A (n_148_16), .B (n_150_19), .C1 (n_146_21), .C2 (n_148_24) );
AOI211_X1 g_146_13 (.ZN (n_146_13), .A (n_150_15), .B (n_148_18), .C1 (n_148_20), .C2 (n_150_23) );
AOI211_X1 g_148_12 (.ZN (n_148_12), .A (n_148_14), .B (n_146_17), .C1 (n_150_19), .C2 (n_148_22) );
AOI211_X1 g_150_11 (.ZN (n_150_11), .A (n_146_13), .B (n_148_16), .C1 (n_148_18), .C2 (n_146_21) );
AOI211_X1 g_149_9 (.ZN (n_149_9), .A (n_148_12), .B (n_150_15), .C1 (n_146_17), .C2 (n_148_20) );
AOI211_X1 g_147_8 (.ZN (n_147_8), .A (n_150_11), .B (n_148_14), .C1 (n_148_16), .C2 (n_150_19) );
AOI211_X1 g_146_6 (.ZN (n_146_6), .A (n_149_9), .B (n_146_13), .C1 (n_150_15), .C2 (n_148_18) );
AOI211_X1 g_144_5 (.ZN (n_144_5), .A (n_147_8), .B (n_148_12), .C1 (n_148_14), .C2 (n_146_17) );
AOI211_X1 g_142_4 (.ZN (n_142_4), .A (n_146_6), .B (n_150_11), .C1 (n_146_13), .C2 (n_148_16) );
AOI211_X1 g_144_3 (.ZN (n_144_3), .A (n_144_5), .B (n_149_9), .C1 (n_148_12), .C2 (n_150_15) );
AOI211_X1 g_142_2 (.ZN (n_142_2), .A (n_142_4), .B (n_147_8), .C1 (n_150_11), .C2 (n_148_14) );
AOI211_X1 g_140_1 (.ZN (n_140_1), .A (n_144_3), .B (n_146_6), .C1 (n_149_9), .C2 (n_146_13) );
AOI211_X1 g_139_3 (.ZN (n_139_3), .A (n_142_2), .B (n_144_5), .C1 (n_147_8), .C2 (n_148_12) );
AOI211_X1 g_141_4 (.ZN (n_141_4), .A (n_140_1), .B (n_142_4), .C1 (n_146_6), .C2 (n_150_11) );
AOI211_X1 g_143_5 (.ZN (n_143_5), .A (n_139_3), .B (n_144_3), .C1 (n_144_5), .C2 (n_149_9) );
AOI211_X1 g_145_6 (.ZN (n_145_6), .A (n_141_4), .B (n_142_2), .C1 (n_142_4), .C2 (n_147_8) );
AOI211_X1 g_146_8 (.ZN (n_146_8), .A (n_143_5), .B (n_140_1), .C1 (n_144_3), .C2 (n_146_6) );
AOI211_X1 g_147_6 (.ZN (n_147_6), .A (n_145_6), .B (n_139_3), .C1 (n_142_2), .C2 (n_144_5) );
AOI211_X1 g_148_8 (.ZN (n_148_8), .A (n_146_8), .B (n_141_4), .C1 (n_140_1), .C2 (n_142_4) );
AOI211_X1 g_147_10 (.ZN (n_147_10), .A (n_147_6), .B (n_143_5), .C1 (n_139_3), .C2 (n_144_3) );
AOI211_X1 g_145_9 (.ZN (n_145_9), .A (n_148_8), .B (n_145_6), .C1 (n_141_4), .C2 (n_142_2) );
AOI211_X1 g_146_7 (.ZN (n_146_7), .A (n_147_10), .B (n_146_8), .C1 (n_143_5), .C2 (n_140_1) );
AOI211_X1 g_145_5 (.ZN (n_145_5), .A (n_145_9), .B (n_147_6), .C1 (n_145_6), .C2 (n_139_3) );
AOI211_X1 g_144_7 (.ZN (n_144_7), .A (n_146_7), .B (n_148_8), .C1 (n_146_8), .C2 (n_141_4) );
AOI211_X1 g_142_6 (.ZN (n_142_6), .A (n_145_5), .B (n_147_10), .C1 (n_147_6), .C2 (n_143_5) );
AOI211_X1 g_143_4 (.ZN (n_143_4), .A (n_144_7), .B (n_145_9), .C1 (n_148_8), .C2 (n_145_6) );
AOI211_X1 g_141_3 (.ZN (n_141_3), .A (n_142_6), .B (n_146_7), .C1 (n_147_10), .C2 (n_146_8) );
AOI211_X1 g_139_2 (.ZN (n_139_2), .A (n_143_4), .B (n_145_5), .C1 (n_145_9), .C2 (n_147_6) );
AOI211_X1 g_137_1 (.ZN (n_137_1), .A (n_141_3), .B (n_144_7), .C1 (n_146_7), .C2 (n_148_8) );
AOI211_X1 g_138_3 (.ZN (n_138_3), .A (n_139_2), .B (n_142_6), .C1 (n_145_5), .C2 (n_147_10) );
AOI211_X1 g_140_4 (.ZN (n_140_4), .A (n_137_1), .B (n_143_4), .C1 (n_144_7), .C2 (n_145_9) );
AOI211_X1 g_142_5 (.ZN (n_142_5), .A (n_138_3), .B (n_141_3), .C1 (n_142_6), .C2 (n_146_7) );
AOI211_X1 g_144_6 (.ZN (n_144_6), .A (n_140_4), .B (n_139_2), .C1 (n_143_4), .C2 (n_145_5) );
AOI211_X1 g_143_8 (.ZN (n_143_8), .A (n_142_5), .B (n_137_1), .C1 (n_141_3), .C2 (n_144_7) );
AOI211_X1 g_145_7 (.ZN (n_145_7), .A (n_144_6), .B (n_138_3), .C1 (n_139_2), .C2 (n_142_6) );
AOI211_X1 g_143_6 (.ZN (n_143_6), .A (n_143_8), .B (n_140_4), .C1 (n_137_1), .C2 (n_143_4) );
AOI211_X1 g_141_5 (.ZN (n_141_5), .A (n_145_7), .B (n_142_5), .C1 (n_138_3), .C2 (n_141_3) );
AOI211_X1 g_140_3 (.ZN (n_140_3), .A (n_143_6), .B (n_144_6), .C1 (n_140_4), .C2 (n_139_2) );
AOI211_X1 g_138_2 (.ZN (n_138_2), .A (n_141_5), .B (n_143_8), .C1 (n_142_5), .C2 (n_137_1) );
AOI211_X1 g_136_1 (.ZN (n_136_1), .A (n_140_3), .B (n_145_7), .C1 (n_144_6), .C2 (n_138_3) );
AOI211_X1 g_135_3 (.ZN (n_135_3), .A (n_138_2), .B (n_143_6), .C1 (n_143_8), .C2 (n_140_4) );
AOI211_X1 g_137_4 (.ZN (n_137_4), .A (n_136_1), .B (n_141_5), .C1 (n_145_7), .C2 (n_142_5) );
AOI211_X1 g_139_5 (.ZN (n_139_5), .A (n_135_3), .B (n_140_3), .C1 (n_143_6), .C2 (n_144_6) );
AOI211_X1 g_141_6 (.ZN (n_141_6), .A (n_137_4), .B (n_138_2), .C1 (n_141_5), .C2 (n_143_8) );
AOI211_X1 g_143_7 (.ZN (n_143_7), .A (n_139_5), .B (n_136_1), .C1 (n_140_3), .C2 (n_145_7) );
AOI211_X1 g_145_8 (.ZN (n_145_8), .A (n_141_6), .B (n_135_3), .C1 (n_138_2), .C2 (n_143_6) );
AOI211_X1 g_147_9 (.ZN (n_147_9), .A (n_143_7), .B (n_137_4), .C1 (n_136_1), .C2 (n_141_5) );
AOI211_X1 g_148_11 (.ZN (n_148_11), .A (n_145_8), .B (n_139_5), .C1 (n_135_3), .C2 (n_140_3) );
AOI211_X1 g_149_13 (.ZN (n_149_13), .A (n_147_9), .B (n_141_6), .C1 (n_137_4), .C2 (n_138_2) );
AOI211_X1 g_147_14 (.ZN (n_147_14), .A (n_148_11), .B (n_143_7), .C1 (n_139_5), .C2 (n_136_1) );
AOI211_X1 g_146_12 (.ZN (n_146_12), .A (n_149_13), .B (n_145_8), .C1 (n_141_6), .C2 (n_135_3) );
AOI211_X1 g_145_10 (.ZN (n_145_10), .A (n_147_14), .B (n_147_9), .C1 (n_143_7), .C2 (n_137_4) );
AOI211_X1 g_144_8 (.ZN (n_144_8), .A (n_146_12), .B (n_148_11), .C1 (n_145_8), .C2 (n_139_5) );
AOI211_X1 g_146_9 (.ZN (n_146_9), .A (n_145_10), .B (n_149_13), .C1 (n_147_9), .C2 (n_141_6) );
AOI211_X1 g_148_10 (.ZN (n_148_10), .A (n_144_8), .B (n_147_14), .C1 (n_148_11), .C2 (n_143_7) );
AOI211_X1 g_146_11 (.ZN (n_146_11), .A (n_146_9), .B (n_146_12), .C1 (n_149_13), .C2 (n_145_8) );
AOI211_X1 g_144_10 (.ZN (n_144_10), .A (n_148_10), .B (n_145_10), .C1 (n_147_14), .C2 (n_147_9) );
AOI211_X1 g_142_9 (.ZN (n_142_9), .A (n_146_11), .B (n_144_8), .C1 (n_146_12), .C2 (n_148_11) );
AOI211_X1 g_141_7 (.ZN (n_141_7), .A (n_144_10), .B (n_146_9), .C1 (n_145_10), .C2 (n_149_13) );
AOI211_X1 g_140_5 (.ZN (n_140_5), .A (n_142_9), .B (n_148_10), .C1 (n_144_8), .C2 (n_147_14) );
AOI211_X1 g_138_4 (.ZN (n_138_4), .A (n_141_7), .B (n_146_11), .C1 (n_146_9), .C2 (n_146_12) );
AOI211_X1 g_136_3 (.ZN (n_136_3), .A (n_140_5), .B (n_144_10), .C1 (n_148_10), .C2 (n_145_10) );
AOI211_X1 g_134_2 (.ZN (n_134_2), .A (n_138_4), .B (n_142_9), .C1 (n_146_11), .C2 (n_144_8) );
AOI211_X1 g_132_1 (.ZN (n_132_1), .A (n_136_3), .B (n_141_7), .C1 (n_144_10), .C2 (n_146_9) );
AOI211_X1 g_131_3 (.ZN (n_131_3), .A (n_134_2), .B (n_140_5), .C1 (n_142_9), .C2 (n_148_10) );
AOI211_X1 g_133_4 (.ZN (n_133_4), .A (n_132_1), .B (n_138_4), .C1 (n_141_7), .C2 (n_146_11) );
AOI211_X1 g_135_5 (.ZN (n_135_5), .A (n_131_3), .B (n_136_3), .C1 (n_140_5), .C2 (n_144_10) );
AOI211_X1 g_134_3 (.ZN (n_134_3), .A (n_133_4), .B (n_134_2), .C1 (n_138_4), .C2 (n_142_9) );
AOI211_X1 g_133_1 (.ZN (n_133_1), .A (n_135_5), .B (n_132_1), .C1 (n_136_3), .C2 (n_141_7) );
AOI211_X1 g_135_2 (.ZN (n_135_2), .A (n_134_3), .B (n_131_3), .C1 (n_134_2), .C2 (n_140_5) );
AOI211_X1 g_136_4 (.ZN (n_136_4), .A (n_133_1), .B (n_133_4), .C1 (n_132_1), .C2 (n_138_4) );
AOI211_X1 g_137_6 (.ZN (n_137_6), .A (n_135_2), .B (n_135_5), .C1 (n_131_3), .C2 (n_136_3) );
AOI211_X1 g_139_7 (.ZN (n_139_7), .A (n_136_4), .B (n_134_3), .C1 (n_133_4), .C2 (n_134_2) );
AOI211_X1 g_138_5 (.ZN (n_138_5), .A (n_137_6), .B (n_133_1), .C1 (n_135_5), .C2 (n_132_1) );
AOI211_X1 g_137_3 (.ZN (n_137_3), .A (n_139_7), .B (n_135_2), .C1 (n_134_3), .C2 (n_131_3) );
AOI211_X1 g_139_4 (.ZN (n_139_4), .A (n_138_5), .B (n_136_4), .C1 (n_133_1), .C2 (n_133_4) );
AOI211_X1 g_140_6 (.ZN (n_140_6), .A (n_137_3), .B (n_137_6), .C1 (n_135_2), .C2 (n_135_5) );
AOI211_X1 g_142_7 (.ZN (n_142_7), .A (n_139_4), .B (n_139_7), .C1 (n_136_4), .C2 (n_134_3) );
AOI211_X1 g_143_9 (.ZN (n_143_9), .A (n_140_6), .B (n_138_5), .C1 (n_137_6), .C2 (n_133_1) );
AOI211_X1 g_141_8 (.ZN (n_141_8), .A (n_142_7), .B (n_137_3), .C1 (n_139_7), .C2 (n_135_2) );
AOI211_X1 g_140_10 (.ZN (n_140_10), .A (n_143_9), .B (n_139_4), .C1 (n_138_5), .C2 (n_136_4) );
AOI211_X1 g_139_8 (.ZN (n_139_8), .A (n_141_8), .B (n_140_6), .C1 (n_137_3), .C2 (n_137_6) );
AOI211_X1 g_138_6 (.ZN (n_138_6), .A (n_140_10), .B (n_142_7), .C1 (n_139_4), .C2 (n_139_7) );
AOI211_X1 g_136_5 (.ZN (n_136_5), .A (n_139_8), .B (n_143_9), .C1 (n_140_6), .C2 (n_138_5) );
AOI211_X1 g_134_4 (.ZN (n_134_4), .A (n_138_6), .B (n_141_8), .C1 (n_142_7), .C2 (n_137_3) );
AOI211_X1 g_132_3 (.ZN (n_132_3), .A (n_136_5), .B (n_140_10), .C1 (n_143_9), .C2 (n_139_4) );
AOI211_X1 g_130_2 (.ZN (n_130_2), .A (n_134_4), .B (n_139_8), .C1 (n_141_8), .C2 (n_140_6) );
AOI211_X1 g_128_1 (.ZN (n_128_1), .A (n_132_3), .B (n_138_6), .C1 (n_140_10), .C2 (n_142_7) );
AOI211_X1 g_127_3 (.ZN (n_127_3), .A (n_130_2), .B (n_136_5), .C1 (n_139_8), .C2 (n_143_9) );
AOI211_X1 g_129_4 (.ZN (n_129_4), .A (n_128_1), .B (n_134_4), .C1 (n_138_6), .C2 (n_141_8) );
AOI211_X1 g_131_5 (.ZN (n_131_5), .A (n_127_3), .B (n_132_3), .C1 (n_136_5), .C2 (n_140_10) );
AOI211_X1 g_130_3 (.ZN (n_130_3), .A (n_129_4), .B (n_130_2), .C1 (n_134_4), .C2 (n_139_8) );
AOI211_X1 g_129_1 (.ZN (n_129_1), .A (n_131_5), .B (n_128_1), .C1 (n_132_3), .C2 (n_138_6) );
AOI211_X1 g_131_2 (.ZN (n_131_2), .A (n_130_3), .B (n_127_3), .C1 (n_130_2), .C2 (n_136_5) );
AOI211_X1 g_132_4 (.ZN (n_132_4), .A (n_129_1), .B (n_129_4), .C1 (n_128_1), .C2 (n_134_4) );
AOI211_X1 g_133_6 (.ZN (n_133_6), .A (n_131_2), .B (n_131_5), .C1 (n_127_3), .C2 (n_132_3) );
AOI211_X1 g_135_7 (.ZN (n_135_7), .A (n_132_4), .B (n_130_3), .C1 (n_129_4), .C2 (n_130_2) );
AOI211_X1 g_134_5 (.ZN (n_134_5), .A (n_133_6), .B (n_129_1), .C1 (n_131_5), .C2 (n_128_1) );
AOI211_X1 g_133_3 (.ZN (n_133_3), .A (n_135_7), .B (n_131_2), .C1 (n_130_3), .C2 (n_127_3) );
AOI211_X1 g_135_4 (.ZN (n_135_4), .A (n_134_5), .B (n_132_4), .C1 (n_129_1), .C2 (n_129_4) );
AOI211_X1 g_136_6 (.ZN (n_136_6), .A (n_133_3), .B (n_133_6), .C1 (n_131_2), .C2 (n_131_5) );
AOI211_X1 g_137_8 (.ZN (n_137_8), .A (n_135_4), .B (n_135_7), .C1 (n_132_4), .C2 (n_130_3) );
AOI211_X1 g_138_10 (.ZN (n_138_10), .A (n_136_6), .B (n_134_5), .C1 (n_133_6), .C2 (n_129_1) );
AOI211_X1 g_140_9 (.ZN (n_140_9), .A (n_137_8), .B (n_133_3), .C1 (n_135_7), .C2 (n_131_2) );
AOI211_X1 g_142_8 (.ZN (n_142_8), .A (n_138_10), .B (n_135_4), .C1 (n_134_5), .C2 (n_132_4) );
AOI211_X1 g_140_7 (.ZN (n_140_7), .A (n_140_9), .B (n_136_6), .C1 (n_133_3), .C2 (n_133_6) );
AOI211_X1 g_141_9 (.ZN (n_141_9), .A (n_142_8), .B (n_137_8), .C1 (n_135_4), .C2 (n_135_7) );
AOI211_X1 g_142_11 (.ZN (n_142_11), .A (n_140_7), .B (n_138_10), .C1 (n_136_6), .C2 (n_134_5) );
AOI211_X1 g_144_12 (.ZN (n_144_12), .A (n_141_9), .B (n_140_9), .C1 (n_137_8), .C2 (n_133_3) );
AOI211_X1 g_143_10 (.ZN (n_143_10), .A (n_142_11), .B (n_142_8), .C1 (n_138_10), .C2 (n_135_4) );
AOI211_X1 g_145_11 (.ZN (n_145_11), .A (n_144_12), .B (n_140_7), .C1 (n_140_9), .C2 (n_136_6) );
AOI211_X1 g_144_9 (.ZN (n_144_9), .A (n_143_10), .B (n_141_9), .C1 (n_142_8), .C2 (n_137_8) );
AOI211_X1 g_146_10 (.ZN (n_146_10), .A (n_145_11), .B (n_142_11), .C1 (n_140_7), .C2 (n_138_10) );
AOI211_X1 g_147_12 (.ZN (n_147_12), .A (n_144_9), .B (n_144_12), .C1 (n_141_9), .C2 (n_140_9) );
AOI211_X1 g_145_13 (.ZN (n_145_13), .A (n_146_10), .B (n_143_10), .C1 (n_142_11), .C2 (n_142_8) );
AOI211_X1 g_144_11 (.ZN (n_144_11), .A (n_147_12), .B (n_145_11), .C1 (n_144_12), .C2 (n_140_7) );
AOI211_X1 g_142_10 (.ZN (n_142_10), .A (n_145_13), .B (n_144_9), .C1 (n_143_10), .C2 (n_141_9) );
AOI211_X1 g_143_12 (.ZN (n_143_12), .A (n_144_11), .B (n_146_10), .C1 (n_145_11), .C2 (n_142_11) );
AOI211_X1 g_141_11 (.ZN (n_141_11), .A (n_142_10), .B (n_147_12), .C1 (n_144_9), .C2 (n_144_12) );
AOI211_X1 g_139_12 (.ZN (n_139_12), .A (n_143_12), .B (n_145_13), .C1 (n_146_10), .C2 (n_143_10) );
AOI211_X1 g_141_13 (.ZN (n_141_13), .A (n_141_11), .B (n_144_11), .C1 (n_147_12), .C2 (n_145_11) );
AOI211_X1 g_140_11 (.ZN (n_140_11), .A (n_139_12), .B (n_142_10), .C1 (n_145_13), .C2 (n_144_9) );
AOI211_X1 g_139_9 (.ZN (n_139_9), .A (n_141_13), .B (n_143_12), .C1 (n_144_11), .C2 (n_146_10) );
AOI211_X1 g_138_7 (.ZN (n_138_7), .A (n_140_11), .B (n_141_11), .C1 (n_142_10), .C2 (n_147_12) );
AOI211_X1 g_137_5 (.ZN (n_137_5), .A (n_139_9), .B (n_139_12), .C1 (n_143_12), .C2 (n_145_13) );
AOI211_X1 g_139_6 (.ZN (n_139_6), .A (n_138_7), .B (n_141_13), .C1 (n_141_11), .C2 (n_144_11) );
AOI211_X1 g_140_8 (.ZN (n_140_8), .A (n_137_5), .B (n_140_11), .C1 (n_139_12), .C2 (n_142_10) );
AOI211_X1 g_141_10 (.ZN (n_141_10), .A (n_139_6), .B (n_139_9), .C1 (n_141_13), .C2 (n_143_12) );
AOI211_X1 g_142_12 (.ZN (n_142_12), .A (n_140_8), .B (n_138_7), .C1 (n_140_11), .C2 (n_141_11) );
AOI211_X1 g_143_14 (.ZN (n_143_14), .A (n_141_10), .B (n_137_5), .C1 (n_139_9), .C2 (n_139_12) );
AOI211_X1 g_145_15 (.ZN (n_145_15), .A (n_142_12), .B (n_139_6), .C1 (n_138_7), .C2 (n_141_13) );
AOI211_X1 g_144_13 (.ZN (n_144_13), .A (n_143_14), .B (n_140_8), .C1 (n_137_5), .C2 (n_140_11) );
AOI211_X1 g_143_11 (.ZN (n_143_11), .A (n_145_15), .B (n_141_10), .C1 (n_139_6), .C2 (n_139_9) );
AOI211_X1 g_145_12 (.ZN (n_145_12), .A (n_144_13), .B (n_142_12), .C1 (n_140_8), .C2 (n_138_7) );
AOI211_X1 g_147_13 (.ZN (n_147_13), .A (n_143_11), .B (n_143_14), .C1 (n_141_10), .C2 (n_137_5) );
AOI211_X1 g_145_14 (.ZN (n_145_14), .A (n_145_12), .B (n_145_15), .C1 (n_142_12), .C2 (n_139_6) );
AOI211_X1 g_143_13 (.ZN (n_143_13), .A (n_147_13), .B (n_144_13), .C1 (n_143_14), .C2 (n_140_8) );
AOI211_X1 g_141_12 (.ZN (n_141_12), .A (n_145_14), .B (n_143_11), .C1 (n_145_15), .C2 (n_141_10) );
AOI211_X1 g_139_11 (.ZN (n_139_11), .A (n_143_13), .B (n_145_12), .C1 (n_144_13), .C2 (n_142_12) );
AOI211_X1 g_138_9 (.ZN (n_138_9), .A (n_141_12), .B (n_147_13), .C1 (n_143_11), .C2 (n_143_14) );
AOI211_X1 g_137_7 (.ZN (n_137_7), .A (n_139_11), .B (n_145_14), .C1 (n_145_12), .C2 (n_145_15) );
AOI211_X1 g_135_6 (.ZN (n_135_6), .A (n_138_9), .B (n_143_13), .C1 (n_147_13), .C2 (n_144_13) );
AOI211_X1 g_133_5 (.ZN (n_133_5), .A (n_137_7), .B (n_141_12), .C1 (n_145_14), .C2 (n_143_11) );
AOI211_X1 g_131_4 (.ZN (n_131_4), .A (n_135_6), .B (n_139_11), .C1 (n_143_13), .C2 (n_145_12) );
AOI211_X1 g_129_3 (.ZN (n_129_3), .A (n_133_5), .B (n_138_9), .C1 (n_141_12), .C2 (n_147_13) );
AOI211_X1 g_127_2 (.ZN (n_127_2), .A (n_131_4), .B (n_137_7), .C1 (n_139_11), .C2 (n_145_14) );
AOI211_X1 g_125_1 (.ZN (n_125_1), .A (n_129_3), .B (n_135_6), .C1 (n_138_9), .C2 (n_143_13) );
AOI211_X1 g_126_3 (.ZN (n_126_3), .A (n_127_2), .B (n_133_5), .C1 (n_137_7), .C2 (n_141_12) );
AOI211_X1 g_128_4 (.ZN (n_128_4), .A (n_125_1), .B (n_131_4), .C1 (n_135_6), .C2 (n_139_11) );
AOI211_X1 g_130_5 (.ZN (n_130_5), .A (n_126_3), .B (n_129_3), .C1 (n_133_5), .C2 (n_138_9) );
AOI211_X1 g_132_6 (.ZN (n_132_6), .A (n_128_4), .B (n_127_2), .C1 (n_131_4), .C2 (n_137_7) );
AOI211_X1 g_134_7 (.ZN (n_134_7), .A (n_130_5), .B (n_125_1), .C1 (n_129_3), .C2 (n_135_6) );
AOI211_X1 g_136_8 (.ZN (n_136_8), .A (n_132_6), .B (n_126_3), .C1 (n_127_2), .C2 (n_133_5) );
AOI211_X1 g_137_10 (.ZN (n_137_10), .A (n_134_7), .B (n_128_4), .C1 (n_125_1), .C2 (n_131_4) );
AOI211_X1 g_138_8 (.ZN (n_138_8), .A (n_136_8), .B (n_130_5), .C1 (n_126_3), .C2 (n_129_3) );
AOI211_X1 g_136_7 (.ZN (n_136_7), .A (n_137_10), .B (n_132_6), .C1 (n_128_4), .C2 (n_127_2) );
AOI211_X1 g_134_6 (.ZN (n_134_6), .A (n_138_8), .B (n_134_7), .C1 (n_130_5), .C2 (n_125_1) );
AOI211_X1 g_132_5 (.ZN (n_132_5), .A (n_136_7), .B (n_136_8), .C1 (n_132_6), .C2 (n_126_3) );
AOI211_X1 g_130_4 (.ZN (n_130_4), .A (n_134_6), .B (n_137_10), .C1 (n_134_7), .C2 (n_128_4) );
AOI211_X1 g_128_3 (.ZN (n_128_3), .A (n_132_5), .B (n_138_8), .C1 (n_136_8), .C2 (n_130_5) );
AOI211_X1 g_126_2 (.ZN (n_126_2), .A (n_130_4), .B (n_136_7), .C1 (n_137_10), .C2 (n_132_6) );
AOI211_X1 g_124_1 (.ZN (n_124_1), .A (n_128_3), .B (n_134_6), .C1 (n_138_8), .C2 (n_134_7) );
AOI211_X1 g_123_3 (.ZN (n_123_3), .A (n_126_2), .B (n_132_5), .C1 (n_136_7), .C2 (n_136_8) );
AOI211_X1 g_125_4 (.ZN (n_125_4), .A (n_124_1), .B (n_130_4), .C1 (n_134_6), .C2 (n_137_10) );
AOI211_X1 g_127_5 (.ZN (n_127_5), .A (n_123_3), .B (n_128_3), .C1 (n_132_5), .C2 (n_138_8) );
AOI211_X1 g_129_6 (.ZN (n_129_6), .A (n_125_4), .B (n_126_2), .C1 (n_130_4), .C2 (n_136_7) );
AOI211_X1 g_131_7 (.ZN (n_131_7), .A (n_127_5), .B (n_124_1), .C1 (n_128_3), .C2 (n_134_6) );
AOI211_X1 g_133_8 (.ZN (n_133_8), .A (n_129_6), .B (n_123_3), .C1 (n_126_2), .C2 (n_132_5) );
AOI211_X1 g_135_9 (.ZN (n_135_9), .A (n_131_7), .B (n_125_4), .C1 (n_124_1), .C2 (n_130_4) );
AOI211_X1 g_136_11 (.ZN (n_136_11), .A (n_133_8), .B (n_127_5), .C1 (n_123_3), .C2 (n_128_3) );
AOI211_X1 g_137_9 (.ZN (n_137_9), .A (n_135_9), .B (n_129_6), .C1 (n_125_4), .C2 (n_126_2) );
AOI211_X1 g_139_10 (.ZN (n_139_10), .A (n_136_11), .B (n_131_7), .C1 (n_127_5), .C2 (n_124_1) );
AOI211_X1 g_138_12 (.ZN (n_138_12), .A (n_137_9), .B (n_133_8), .C1 (n_129_6), .C2 (n_123_3) );
AOI211_X1 g_140_13 (.ZN (n_140_13), .A (n_139_10), .B (n_135_9), .C1 (n_131_7), .C2 (n_125_4) );
AOI211_X1 g_142_14 (.ZN (n_142_14), .A (n_138_12), .B (n_136_11), .C1 (n_133_8), .C2 (n_127_5) );
AOI211_X1 g_144_15 (.ZN (n_144_15), .A (n_140_13), .B (n_137_9), .C1 (n_135_9), .C2 (n_129_6) );
AOI211_X1 g_146_14 (.ZN (n_146_14), .A (n_142_14), .B (n_139_10), .C1 (n_136_11), .C2 (n_131_7) );
AOI211_X1 g_147_16 (.ZN (n_147_16), .A (n_144_15), .B (n_138_12), .C1 (n_137_9), .C2 (n_133_8) );
AOI211_X1 g_149_17 (.ZN (n_149_17), .A (n_146_14), .B (n_140_13), .C1 (n_139_10), .C2 (n_135_9) );
AOI211_X1 g_148_15 (.ZN (n_148_15), .A (n_147_16), .B (n_142_14), .C1 (n_138_12), .C2 (n_136_11) );
AOI211_X1 g_146_16 (.ZN (n_146_16), .A (n_149_17), .B (n_144_15), .C1 (n_140_13), .C2 (n_137_9) );
AOI211_X1 g_147_18 (.ZN (n_147_18), .A (n_148_15), .B (n_146_14), .C1 (n_142_14), .C2 (n_139_10) );
AOI211_X1 g_145_17 (.ZN (n_145_17), .A (n_146_16), .B (n_147_16), .C1 (n_144_15), .C2 (n_138_12) );
AOI211_X1 g_146_15 (.ZN (n_146_15), .A (n_147_18), .B (n_149_17), .C1 (n_146_14), .C2 (n_140_13) );
AOI211_X1 g_144_14 (.ZN (n_144_14), .A (n_145_17), .B (n_148_15), .C1 (n_147_16), .C2 (n_142_14) );
AOI211_X1 g_142_13 (.ZN (n_142_13), .A (n_146_15), .B (n_146_16), .C1 (n_149_17), .C2 (n_144_15) );
AOI211_X1 g_140_12 (.ZN (n_140_12), .A (n_144_14), .B (n_147_18), .C1 (n_148_15), .C2 (n_146_14) );
AOI211_X1 g_138_11 (.ZN (n_138_11), .A (n_142_13), .B (n_145_17), .C1 (n_146_16), .C2 (n_147_16) );
AOI211_X1 g_136_10 (.ZN (n_136_10), .A (n_140_12), .B (n_146_15), .C1 (n_147_18), .C2 (n_149_17) );
AOI211_X1 g_135_8 (.ZN (n_135_8), .A (n_138_11), .B (n_144_14), .C1 (n_145_17), .C2 (n_148_15) );
AOI211_X1 g_133_7 (.ZN (n_133_7), .A (n_136_10), .B (n_142_13), .C1 (n_146_15), .C2 (n_146_16) );
AOI211_X1 g_131_6 (.ZN (n_131_6), .A (n_135_8), .B (n_140_12), .C1 (n_144_14), .C2 (n_147_18) );
AOI211_X1 g_129_5 (.ZN (n_129_5), .A (n_133_7), .B (n_138_11), .C1 (n_142_13), .C2 (n_145_17) );
AOI211_X1 g_127_4 (.ZN (n_127_4), .A (n_131_6), .B (n_136_10), .C1 (n_140_12), .C2 (n_146_15) );
AOI211_X1 g_125_3 (.ZN (n_125_3), .A (n_129_5), .B (n_135_8), .C1 (n_138_11), .C2 (n_144_14) );
AOI211_X1 g_123_2 (.ZN (n_123_2), .A (n_127_4), .B (n_133_7), .C1 (n_136_10), .C2 (n_142_13) );
AOI211_X1 g_121_1 (.ZN (n_121_1), .A (n_125_3), .B (n_131_6), .C1 (n_135_8), .C2 (n_140_12) );
AOI211_X1 g_122_3 (.ZN (n_122_3), .A (n_123_2), .B (n_129_5), .C1 (n_133_7), .C2 (n_138_11) );
AOI211_X1 g_124_4 (.ZN (n_124_4), .A (n_121_1), .B (n_127_4), .C1 (n_131_6), .C2 (n_136_10) );
AOI211_X1 g_126_5 (.ZN (n_126_5), .A (n_122_3), .B (n_125_3), .C1 (n_129_5), .C2 (n_135_8) );
AOI211_X1 g_128_6 (.ZN (n_128_6), .A (n_124_4), .B (n_123_2), .C1 (n_127_4), .C2 (n_133_7) );
AOI211_X1 g_130_7 (.ZN (n_130_7), .A (n_126_5), .B (n_121_1), .C1 (n_125_3), .C2 (n_131_6) );
AOI211_X1 g_132_8 (.ZN (n_132_8), .A (n_128_6), .B (n_122_3), .C1 (n_123_2), .C2 (n_129_5) );
AOI211_X1 g_134_9 (.ZN (n_134_9), .A (n_130_7), .B (n_124_4), .C1 (n_121_1), .C2 (n_127_4) );
AOI211_X1 g_132_10 (.ZN (n_132_10), .A (n_132_8), .B (n_126_5), .C1 (n_122_3), .C2 (n_125_3) );
AOI211_X1 g_131_8 (.ZN (n_131_8), .A (n_134_9), .B (n_128_6), .C1 (n_124_4), .C2 (n_123_2) );
AOI211_X1 g_130_6 (.ZN (n_130_6), .A (n_132_10), .B (n_130_7), .C1 (n_126_5), .C2 (n_121_1) );
AOI211_X1 g_128_5 (.ZN (n_128_5), .A (n_131_8), .B (n_132_8), .C1 (n_128_6), .C2 (n_122_3) );
AOI211_X1 g_126_4 (.ZN (n_126_4), .A (n_130_6), .B (n_134_9), .C1 (n_130_7), .C2 (n_124_4) );
AOI211_X1 g_124_3 (.ZN (n_124_3), .A (n_128_5), .B (n_132_10), .C1 (n_132_8), .C2 (n_126_5) );
AOI211_X1 g_122_2 (.ZN (n_122_2), .A (n_126_4), .B (n_131_8), .C1 (n_134_9), .C2 (n_128_6) );
AOI211_X1 g_120_1 (.ZN (n_120_1), .A (n_124_3), .B (n_130_6), .C1 (n_132_10), .C2 (n_130_7) );
AOI211_X1 g_119_3 (.ZN (n_119_3), .A (n_122_2), .B (n_128_5), .C1 (n_131_8), .C2 (n_132_8) );
AOI211_X1 g_121_4 (.ZN (n_121_4), .A (n_120_1), .B (n_126_4), .C1 (n_130_6), .C2 (n_134_9) );
AOI211_X1 g_123_5 (.ZN (n_123_5), .A (n_119_3), .B (n_124_3), .C1 (n_128_5), .C2 (n_132_10) );
AOI211_X1 g_125_6 (.ZN (n_125_6), .A (n_121_4), .B (n_122_2), .C1 (n_126_4), .C2 (n_131_8) );
AOI211_X1 g_127_7 (.ZN (n_127_7), .A (n_123_5), .B (n_120_1), .C1 (n_124_3), .C2 (n_130_6) );
AOI211_X1 g_129_8 (.ZN (n_129_8), .A (n_125_6), .B (n_119_3), .C1 (n_122_2), .C2 (n_128_5) );
AOI211_X1 g_131_9 (.ZN (n_131_9), .A (n_127_7), .B (n_121_4), .C1 (n_120_1), .C2 (n_126_4) );
AOI211_X1 g_132_7 (.ZN (n_132_7), .A (n_129_8), .B (n_123_5), .C1 (n_119_3), .C2 (n_124_3) );
AOI211_X1 g_133_9 (.ZN (n_133_9), .A (n_131_9), .B (n_125_6), .C1 (n_121_4), .C2 (n_122_2) );
AOI211_X1 g_134_11 (.ZN (n_134_11), .A (n_132_7), .B (n_127_7), .C1 (n_123_5), .C2 (n_120_1) );
AOI211_X1 g_136_12 (.ZN (n_136_12), .A (n_133_9), .B (n_129_8), .C1 (n_125_6), .C2 (n_119_3) );
AOI211_X1 g_135_10 (.ZN (n_135_10), .A (n_134_11), .B (n_131_9), .C1 (n_127_7), .C2 (n_121_4) );
AOI211_X1 g_134_8 (.ZN (n_134_8), .A (n_136_12), .B (n_132_7), .C1 (n_129_8), .C2 (n_123_5) );
AOI211_X1 g_136_9 (.ZN (n_136_9), .A (n_135_10), .B (n_133_9), .C1 (n_131_9), .C2 (n_125_6) );
AOI211_X1 g_137_11 (.ZN (n_137_11), .A (n_134_8), .B (n_134_11), .C1 (n_132_7), .C2 (n_127_7) );
AOI211_X1 g_138_13 (.ZN (n_138_13), .A (n_136_9), .B (n_136_12), .C1 (n_133_9), .C2 (n_129_8) );
AOI211_X1 g_140_14 (.ZN (n_140_14), .A (n_137_11), .B (n_135_10), .C1 (n_134_11), .C2 (n_131_9) );
AOI211_X1 g_142_15 (.ZN (n_142_15), .A (n_138_13), .B (n_134_8), .C1 (n_136_12), .C2 (n_132_7) );
AOI211_X1 g_144_16 (.ZN (n_144_16), .A (n_140_14), .B (n_136_9), .C1 (n_135_10), .C2 (n_133_9) );
AOI211_X1 g_145_18 (.ZN (n_145_18), .A (n_142_15), .B (n_137_11), .C1 (n_134_8), .C2 (n_134_11) );
AOI211_X1 g_147_17 (.ZN (n_147_17), .A (n_144_16), .B (n_138_13), .C1 (n_136_9), .C2 (n_136_12) );
AOI211_X1 g_145_16 (.ZN (n_145_16), .A (n_145_18), .B (n_140_14), .C1 (n_137_11), .C2 (n_135_10) );
AOI211_X1 g_143_15 (.ZN (n_143_15), .A (n_147_17), .B (n_142_15), .C1 (n_138_13), .C2 (n_134_8) );
AOI211_X1 g_141_14 (.ZN (n_141_14), .A (n_145_16), .B (n_144_16), .C1 (n_140_14), .C2 (n_136_9) );
AOI211_X1 g_139_13 (.ZN (n_139_13), .A (n_143_15), .B (n_145_18), .C1 (n_142_15), .C2 (n_137_11) );
AOI211_X1 g_137_12 (.ZN (n_137_12), .A (n_141_14), .B (n_147_17), .C1 (n_144_16), .C2 (n_138_13) );
AOI211_X1 g_135_11 (.ZN (n_135_11), .A (n_139_13), .B (n_145_16), .C1 (n_145_18), .C2 (n_140_14) );
AOI211_X1 g_133_10 (.ZN (n_133_10), .A (n_137_12), .B (n_143_15), .C1 (n_147_17), .C2 (n_142_15) );
AOI211_X1 g_134_12 (.ZN (n_134_12), .A (n_135_11), .B (n_141_14), .C1 (n_145_16), .C2 (n_144_16) );
AOI211_X1 g_136_13 (.ZN (n_136_13), .A (n_133_10), .B (n_139_13), .C1 (n_143_15), .C2 (n_145_18) );
AOI211_X1 g_138_14 (.ZN (n_138_14), .A (n_134_12), .B (n_137_12), .C1 (n_141_14), .C2 (n_147_17) );
AOI211_X1 g_140_15 (.ZN (n_140_15), .A (n_136_13), .B (n_135_11), .C1 (n_139_13), .C2 (n_145_16) );
AOI211_X1 g_142_16 (.ZN (n_142_16), .A (n_138_14), .B (n_133_10), .C1 (n_137_12), .C2 (n_143_15) );
AOI211_X1 g_144_17 (.ZN (n_144_17), .A (n_140_15), .B (n_134_12), .C1 (n_135_11), .C2 (n_141_14) );
AOI211_X1 g_145_19 (.ZN (n_145_19), .A (n_142_16), .B (n_136_13), .C1 (n_133_10), .C2 (n_139_13) );
AOI211_X1 g_143_18 (.ZN (n_143_18), .A (n_144_17), .B (n_138_14), .C1 (n_134_12), .C2 (n_137_12) );
AOI211_X1 g_141_17 (.ZN (n_141_17), .A (n_145_19), .B (n_140_15), .C1 (n_136_13), .C2 (n_135_11) );
AOI211_X1 g_143_16 (.ZN (n_143_16), .A (n_143_18), .B (n_142_16), .C1 (n_138_14), .C2 (n_133_10) );
AOI211_X1 g_141_15 (.ZN (n_141_15), .A (n_141_17), .B (n_144_17), .C1 (n_140_15), .C2 (n_134_12) );
AOI211_X1 g_139_14 (.ZN (n_139_14), .A (n_143_16), .B (n_145_19), .C1 (n_142_16), .C2 (n_136_13) );
AOI211_X1 g_137_13 (.ZN (n_137_13), .A (n_141_15), .B (n_143_18), .C1 (n_144_17), .C2 (n_138_14) );
AOI211_X1 g_135_12 (.ZN (n_135_12), .A (n_139_14), .B (n_141_17), .C1 (n_145_19), .C2 (n_140_15) );
AOI211_X1 g_134_10 (.ZN (n_134_10), .A (n_137_13), .B (n_143_16), .C1 (n_143_18), .C2 (n_142_16) );
AOI211_X1 g_132_9 (.ZN (n_132_9), .A (n_135_12), .B (n_141_15), .C1 (n_141_17), .C2 (n_144_17) );
AOI211_X1 g_130_8 (.ZN (n_130_8), .A (n_134_10), .B (n_139_14), .C1 (n_143_16), .C2 (n_145_19) );
AOI211_X1 g_128_7 (.ZN (n_128_7), .A (n_132_9), .B (n_137_13), .C1 (n_141_15), .C2 (n_143_18) );
AOI211_X1 g_126_6 (.ZN (n_126_6), .A (n_130_8), .B (n_135_12), .C1 (n_139_14), .C2 (n_141_17) );
AOI211_X1 g_124_5 (.ZN (n_124_5), .A (n_128_7), .B (n_134_10), .C1 (n_137_13), .C2 (n_143_16) );
AOI211_X1 g_122_4 (.ZN (n_122_4), .A (n_126_6), .B (n_132_9), .C1 (n_135_12), .C2 (n_141_15) );
AOI211_X1 g_120_3 (.ZN (n_120_3), .A (n_124_5), .B (n_130_8), .C1 (n_134_10), .C2 (n_139_14) );
AOI211_X1 g_118_2 (.ZN (n_118_2), .A (n_122_4), .B (n_128_7), .C1 (n_132_9), .C2 (n_137_13) );
AOI211_X1 g_116_1 (.ZN (n_116_1), .A (n_120_3), .B (n_126_6), .C1 (n_130_8), .C2 (n_135_12) );
AOI211_X1 g_115_3 (.ZN (n_115_3), .A (n_118_2), .B (n_124_5), .C1 (n_128_7), .C2 (n_134_10) );
AOI211_X1 g_117_4 (.ZN (n_117_4), .A (n_116_1), .B (n_122_4), .C1 (n_126_6), .C2 (n_132_9) );
AOI211_X1 g_119_5 (.ZN (n_119_5), .A (n_115_3), .B (n_120_3), .C1 (n_124_5), .C2 (n_130_8) );
AOI211_X1 g_118_3 (.ZN (n_118_3), .A (n_117_4), .B (n_118_2), .C1 (n_122_4), .C2 (n_128_7) );
AOI211_X1 g_117_1 (.ZN (n_117_1), .A (n_119_5), .B (n_116_1), .C1 (n_120_3), .C2 (n_126_6) );
AOI211_X1 g_119_2 (.ZN (n_119_2), .A (n_118_3), .B (n_115_3), .C1 (n_118_2), .C2 (n_124_5) );
AOI211_X1 g_120_4 (.ZN (n_120_4), .A (n_117_1), .B (n_117_4), .C1 (n_116_1), .C2 (n_122_4) );
AOI211_X1 g_121_6 (.ZN (n_121_6), .A (n_119_2), .B (n_119_5), .C1 (n_115_3), .C2 (n_120_3) );
AOI211_X1 g_123_7 (.ZN (n_123_7), .A (n_120_4), .B (n_118_3), .C1 (n_117_4), .C2 (n_118_2) );
AOI211_X1 g_122_5 (.ZN (n_122_5), .A (n_121_6), .B (n_117_1), .C1 (n_119_5), .C2 (n_116_1) );
AOI211_X1 g_121_3 (.ZN (n_121_3), .A (n_123_7), .B (n_119_2), .C1 (n_118_3), .C2 (n_115_3) );
AOI211_X1 g_123_4 (.ZN (n_123_4), .A (n_122_5), .B (n_120_4), .C1 (n_117_1), .C2 (n_117_4) );
AOI211_X1 g_124_6 (.ZN (n_124_6), .A (n_121_3), .B (n_121_6), .C1 (n_119_2), .C2 (n_119_5) );
AOI211_X1 g_125_8 (.ZN (n_125_8), .A (n_123_4), .B (n_123_7), .C1 (n_120_4), .C2 (n_118_3) );
AOI211_X1 g_127_9 (.ZN (n_127_9), .A (n_124_6), .B (n_122_5), .C1 (n_121_6), .C2 (n_117_1) );
AOI211_X1 g_126_7 (.ZN (n_126_7), .A (n_125_8), .B (n_121_3), .C1 (n_123_7), .C2 (n_119_2) );
AOI211_X1 g_125_5 (.ZN (n_125_5), .A (n_127_9), .B (n_123_4), .C1 (n_122_5), .C2 (n_120_4) );
AOI211_X1 g_127_6 (.ZN (n_127_6), .A (n_126_7), .B (n_124_6), .C1 (n_121_3), .C2 (n_121_6) );
AOI211_X1 g_129_7 (.ZN (n_129_7), .A (n_125_5), .B (n_125_8), .C1 (n_123_4), .C2 (n_123_7) );
AOI211_X1 g_130_9 (.ZN (n_130_9), .A (n_127_6), .B (n_127_9), .C1 (n_124_6), .C2 (n_122_5) );
AOI211_X1 g_128_8 (.ZN (n_128_8), .A (n_129_7), .B (n_126_7), .C1 (n_125_8), .C2 (n_121_3) );
AOI211_X1 g_129_10 (.ZN (n_129_10), .A (n_130_9), .B (n_125_5), .C1 (n_127_9), .C2 (n_123_4) );
AOI211_X1 g_131_11 (.ZN (n_131_11), .A (n_128_8), .B (n_127_6), .C1 (n_126_7), .C2 (n_124_6) );
AOI211_X1 g_133_12 (.ZN (n_133_12), .A (n_129_10), .B (n_129_7), .C1 (n_125_5), .C2 (n_125_8) );
AOI211_X1 g_135_13 (.ZN (n_135_13), .A (n_131_11), .B (n_130_9), .C1 (n_127_6), .C2 (n_127_9) );
AOI211_X1 g_137_14 (.ZN (n_137_14), .A (n_133_12), .B (n_128_8), .C1 (n_129_7), .C2 (n_126_7) );
AOI211_X1 g_139_15 (.ZN (n_139_15), .A (n_135_13), .B (n_129_10), .C1 (n_130_9), .C2 (n_125_5) );
AOI211_X1 g_141_16 (.ZN (n_141_16), .A (n_137_14), .B (n_131_11), .C1 (n_128_8), .C2 (n_127_6) );
AOI211_X1 g_143_17 (.ZN (n_143_17), .A (n_139_15), .B (n_133_12), .C1 (n_129_10), .C2 (n_129_7) );
AOI211_X1 g_141_18 (.ZN (n_141_18), .A (n_141_16), .B (n_135_13), .C1 (n_131_11), .C2 (n_130_9) );
AOI211_X1 g_140_16 (.ZN (n_140_16), .A (n_143_17), .B (n_137_14), .C1 (n_133_12), .C2 (n_128_8) );
AOI211_X1 g_138_15 (.ZN (n_138_15), .A (n_141_18), .B (n_139_15), .C1 (n_135_13), .C2 (n_129_10) );
AOI211_X1 g_136_14 (.ZN (n_136_14), .A (n_140_16), .B (n_141_16), .C1 (n_137_14), .C2 (n_131_11) );
AOI211_X1 g_134_13 (.ZN (n_134_13), .A (n_138_15), .B (n_143_17), .C1 (n_139_15), .C2 (n_133_12) );
AOI211_X1 g_133_11 (.ZN (n_133_11), .A (n_136_14), .B (n_141_18), .C1 (n_141_16), .C2 (n_135_13) );
AOI211_X1 g_131_10 (.ZN (n_131_10), .A (n_134_13), .B (n_140_16), .C1 (n_143_17), .C2 (n_137_14) );
AOI211_X1 g_129_9 (.ZN (n_129_9), .A (n_133_11), .B (n_138_15), .C1 (n_141_18), .C2 (n_139_15) );
AOI211_X1 g_127_8 (.ZN (n_127_8), .A (n_131_10), .B (n_136_14), .C1 (n_140_16), .C2 (n_141_16) );
AOI211_X1 g_125_7 (.ZN (n_125_7), .A (n_129_9), .B (n_134_13), .C1 (n_138_15), .C2 (n_143_17) );
AOI211_X1 g_123_6 (.ZN (n_123_6), .A (n_127_8), .B (n_133_11), .C1 (n_136_14), .C2 (n_141_18) );
AOI211_X1 g_121_5 (.ZN (n_121_5), .A (n_125_7), .B (n_131_10), .C1 (n_134_13), .C2 (n_140_16) );
AOI211_X1 g_119_4 (.ZN (n_119_4), .A (n_123_6), .B (n_129_9), .C1 (n_133_11), .C2 (n_138_15) );
AOI211_X1 g_117_3 (.ZN (n_117_3), .A (n_121_5), .B (n_127_8), .C1 (n_131_10), .C2 (n_136_14) );
AOI211_X1 g_115_2 (.ZN (n_115_2), .A (n_119_4), .B (n_125_7), .C1 (n_129_9), .C2 (n_134_13) );
AOI211_X1 g_113_1 (.ZN (n_113_1), .A (n_117_3), .B (n_123_6), .C1 (n_127_8), .C2 (n_133_11) );
AOI211_X1 g_114_3 (.ZN (n_114_3), .A (n_115_2), .B (n_121_5), .C1 (n_125_7), .C2 (n_131_10) );
AOI211_X1 g_116_4 (.ZN (n_116_4), .A (n_113_1), .B (n_119_4), .C1 (n_123_6), .C2 (n_129_9) );
AOI211_X1 g_118_5 (.ZN (n_118_5), .A (n_114_3), .B (n_117_3), .C1 (n_121_5), .C2 (n_127_8) );
AOI211_X1 g_120_6 (.ZN (n_120_6), .A (n_116_4), .B (n_115_2), .C1 (n_119_4), .C2 (n_125_7) );
AOI211_X1 g_122_7 (.ZN (n_122_7), .A (n_118_5), .B (n_113_1), .C1 (n_117_3), .C2 (n_123_6) );
AOI211_X1 g_124_8 (.ZN (n_124_8), .A (n_120_6), .B (n_114_3), .C1 (n_115_2), .C2 (n_121_5) );
AOI211_X1 g_126_9 (.ZN (n_126_9), .A (n_122_7), .B (n_116_4), .C1 (n_113_1), .C2 (n_119_4) );
AOI211_X1 g_128_10 (.ZN (n_128_10), .A (n_124_8), .B (n_118_5), .C1 (n_114_3), .C2 (n_117_3) );
AOI211_X1 g_130_11 (.ZN (n_130_11), .A (n_126_9), .B (n_120_6), .C1 (n_116_4), .C2 (n_115_2) );
AOI211_X1 g_132_12 (.ZN (n_132_12), .A (n_128_10), .B (n_122_7), .C1 (n_118_5), .C2 (n_113_1) );
AOI211_X1 g_133_14 (.ZN (n_133_14), .A (n_130_11), .B (n_124_8), .C1 (n_120_6), .C2 (n_114_3) );
AOI211_X1 g_135_15 (.ZN (n_135_15), .A (n_132_12), .B (n_126_9), .C1 (n_122_7), .C2 (n_116_4) );
AOI211_X1 g_137_16 (.ZN (n_137_16), .A (n_133_14), .B (n_128_10), .C1 (n_124_8), .C2 (n_118_5) );
AOI211_X1 g_139_17 (.ZN (n_139_17), .A (n_135_15), .B (n_130_11), .C1 (n_126_9), .C2 (n_120_6) );
AOI211_X1 g_140_19 (.ZN (n_140_19), .A (n_137_16), .B (n_132_12), .C1 (n_128_10), .C2 (n_122_7) );
AOI211_X1 g_142_18 (.ZN (n_142_18), .A (n_139_17), .B (n_133_14), .C1 (n_130_11), .C2 (n_124_8) );
AOI211_X1 g_140_17 (.ZN (n_140_17), .A (n_140_19), .B (n_135_15), .C1 (n_132_12), .C2 (n_126_9) );
AOI211_X1 g_138_16 (.ZN (n_138_16), .A (n_142_18), .B (n_137_16), .C1 (n_133_14), .C2 (n_128_10) );
AOI211_X1 g_136_15 (.ZN (n_136_15), .A (n_140_17), .B (n_139_17), .C1 (n_135_15), .C2 (n_130_11) );
AOI211_X1 g_134_14 (.ZN (n_134_14), .A (n_138_16), .B (n_140_19), .C1 (n_137_16), .C2 (n_132_12) );
AOI211_X1 g_132_13 (.ZN (n_132_13), .A (n_136_15), .B (n_142_18), .C1 (n_139_17), .C2 (n_133_14) );
AOI211_X1 g_130_12 (.ZN (n_130_12), .A (n_134_14), .B (n_140_17), .C1 (n_140_19), .C2 (n_135_15) );
AOI211_X1 g_132_11 (.ZN (n_132_11), .A (n_132_13), .B (n_138_16), .C1 (n_142_18), .C2 (n_137_16) );
AOI211_X1 g_130_10 (.ZN (n_130_10), .A (n_130_12), .B (n_136_15), .C1 (n_140_17), .C2 (n_139_17) );
AOI211_X1 g_128_9 (.ZN (n_128_9), .A (n_132_11), .B (n_134_14), .C1 (n_138_16), .C2 (n_140_19) );
AOI211_X1 g_126_8 (.ZN (n_126_8), .A (n_130_10), .B (n_132_13), .C1 (n_136_15), .C2 (n_142_18) );
AOI211_X1 g_124_7 (.ZN (n_124_7), .A (n_128_9), .B (n_130_12), .C1 (n_134_14), .C2 (n_140_17) );
AOI211_X1 g_122_6 (.ZN (n_122_6), .A (n_126_8), .B (n_132_11), .C1 (n_132_13), .C2 (n_138_16) );
AOI211_X1 g_120_5 (.ZN (n_120_5), .A (n_124_7), .B (n_130_10), .C1 (n_130_12), .C2 (n_136_15) );
AOI211_X1 g_118_4 (.ZN (n_118_4), .A (n_122_6), .B (n_128_9), .C1 (n_132_11), .C2 (n_134_14) );
AOI211_X1 g_116_3 (.ZN (n_116_3), .A (n_120_5), .B (n_126_8), .C1 (n_130_10), .C2 (n_132_13) );
AOI211_X1 g_114_2 (.ZN (n_114_2), .A (n_118_4), .B (n_124_7), .C1 (n_128_9), .C2 (n_130_12) );
AOI211_X1 g_112_1 (.ZN (n_112_1), .A (n_116_3), .B (n_122_6), .C1 (n_126_8), .C2 (n_132_11) );
AOI211_X1 g_111_3 (.ZN (n_111_3), .A (n_114_2), .B (n_120_5), .C1 (n_124_7), .C2 (n_130_10) );
AOI211_X1 g_113_4 (.ZN (n_113_4), .A (n_112_1), .B (n_118_4), .C1 (n_122_6), .C2 (n_128_9) );
AOI211_X1 g_115_5 (.ZN (n_115_5), .A (n_111_3), .B (n_116_3), .C1 (n_120_5), .C2 (n_126_8) );
AOI211_X1 g_117_6 (.ZN (n_117_6), .A (n_113_4), .B (n_114_2), .C1 (n_118_4), .C2 (n_124_7) );
AOI211_X1 g_119_7 (.ZN (n_119_7), .A (n_115_5), .B (n_112_1), .C1 (n_116_3), .C2 (n_122_6) );
AOI211_X1 g_121_8 (.ZN (n_121_8), .A (n_117_6), .B (n_111_3), .C1 (n_114_2), .C2 (n_120_5) );
AOI211_X1 g_123_9 (.ZN (n_123_9), .A (n_119_7), .B (n_113_4), .C1 (n_112_1), .C2 (n_118_4) );
AOI211_X1 g_125_10 (.ZN (n_125_10), .A (n_121_8), .B (n_115_5), .C1 (n_111_3), .C2 (n_116_3) );
AOI211_X1 g_127_11 (.ZN (n_127_11), .A (n_123_9), .B (n_117_6), .C1 (n_113_4), .C2 (n_114_2) );
AOI211_X1 g_129_12 (.ZN (n_129_12), .A (n_125_10), .B (n_119_7), .C1 (n_115_5), .C2 (n_112_1) );
AOI211_X1 g_131_13 (.ZN (n_131_13), .A (n_127_11), .B (n_121_8), .C1 (n_117_6), .C2 (n_111_3) );
AOI211_X1 g_129_14 (.ZN (n_129_14), .A (n_129_12), .B (n_123_9), .C1 (n_119_7), .C2 (n_113_4) );
AOI211_X1 g_128_12 (.ZN (n_128_12), .A (n_131_13), .B (n_125_10), .C1 (n_121_8), .C2 (n_115_5) );
AOI211_X1 g_127_10 (.ZN (n_127_10), .A (n_129_14), .B (n_127_11), .C1 (n_123_9), .C2 (n_117_6) );
AOI211_X1 g_125_9 (.ZN (n_125_9), .A (n_128_12), .B (n_129_12), .C1 (n_125_10), .C2 (n_119_7) );
AOI211_X1 g_123_8 (.ZN (n_123_8), .A (n_127_10), .B (n_131_13), .C1 (n_127_11), .C2 (n_121_8) );
AOI211_X1 g_121_7 (.ZN (n_121_7), .A (n_125_9), .B (n_129_14), .C1 (n_129_12), .C2 (n_123_9) );
AOI211_X1 g_119_6 (.ZN (n_119_6), .A (n_123_8), .B (n_128_12), .C1 (n_131_13), .C2 (n_125_10) );
AOI211_X1 g_117_5 (.ZN (n_117_5), .A (n_121_7), .B (n_127_10), .C1 (n_129_14), .C2 (n_127_11) );
AOI211_X1 g_115_4 (.ZN (n_115_4), .A (n_119_6), .B (n_125_9), .C1 (n_128_12), .C2 (n_129_12) );
AOI211_X1 g_113_3 (.ZN (n_113_3), .A (n_117_5), .B (n_123_8), .C1 (n_127_10), .C2 (n_131_13) );
AOI211_X1 g_111_2 (.ZN (n_111_2), .A (n_115_4), .B (n_121_7), .C1 (n_125_9), .C2 (n_129_14) );
AOI211_X1 g_109_1 (.ZN (n_109_1), .A (n_113_3), .B (n_119_6), .C1 (n_123_8), .C2 (n_128_12) );
AOI211_X1 g_110_3 (.ZN (n_110_3), .A (n_111_2), .B (n_117_5), .C1 (n_121_7), .C2 (n_127_10) );
AOI211_X1 g_112_4 (.ZN (n_112_4), .A (n_109_1), .B (n_115_4), .C1 (n_119_6), .C2 (n_125_9) );
AOI211_X1 g_114_5 (.ZN (n_114_5), .A (n_110_3), .B (n_113_3), .C1 (n_117_5), .C2 (n_123_8) );
AOI211_X1 g_116_6 (.ZN (n_116_6), .A (n_112_4), .B (n_111_2), .C1 (n_115_4), .C2 (n_121_7) );
AOI211_X1 g_118_7 (.ZN (n_118_7), .A (n_114_5), .B (n_109_1), .C1 (n_113_3), .C2 (n_119_6) );
AOI211_X1 g_120_8 (.ZN (n_120_8), .A (n_116_6), .B (n_110_3), .C1 (n_111_2), .C2 (n_117_5) );
AOI211_X1 g_122_9 (.ZN (n_122_9), .A (n_118_7), .B (n_112_4), .C1 (n_109_1), .C2 (n_115_4) );
AOI211_X1 g_124_10 (.ZN (n_124_10), .A (n_120_8), .B (n_114_5), .C1 (n_110_3), .C2 (n_113_3) );
AOI211_X1 g_126_11 (.ZN (n_126_11), .A (n_122_9), .B (n_116_6), .C1 (n_112_4), .C2 (n_111_2) );
AOI211_X1 g_127_13 (.ZN (n_127_13), .A (n_124_10), .B (n_118_7), .C1 (n_114_5), .C2 (n_109_1) );
AOI211_X1 g_128_11 (.ZN (n_128_11), .A (n_126_11), .B (n_120_8), .C1 (n_116_6), .C2 (n_110_3) );
AOI211_X1 g_126_10 (.ZN (n_126_10), .A (n_127_13), .B (n_122_9), .C1 (n_118_7), .C2 (n_112_4) );
AOI211_X1 g_124_9 (.ZN (n_124_9), .A (n_128_11), .B (n_124_10), .C1 (n_120_8), .C2 (n_114_5) );
AOI211_X1 g_122_8 (.ZN (n_122_8), .A (n_126_10), .B (n_126_11), .C1 (n_122_9), .C2 (n_116_6) );
AOI211_X1 g_120_7 (.ZN (n_120_7), .A (n_124_9), .B (n_127_13), .C1 (n_124_10), .C2 (n_118_7) );
AOI211_X1 g_118_6 (.ZN (n_118_6), .A (n_122_8), .B (n_128_11), .C1 (n_126_11), .C2 (n_120_8) );
AOI211_X1 g_116_5 (.ZN (n_116_5), .A (n_120_7), .B (n_126_10), .C1 (n_127_13), .C2 (n_122_9) );
AOI211_X1 g_114_4 (.ZN (n_114_4), .A (n_118_6), .B (n_124_9), .C1 (n_128_11), .C2 (n_124_10) );
AOI211_X1 g_112_3 (.ZN (n_112_3), .A (n_116_5), .B (n_122_8), .C1 (n_126_10), .C2 (n_126_11) );
AOI211_X1 g_110_2 (.ZN (n_110_2), .A (n_114_4), .B (n_120_7), .C1 (n_124_9), .C2 (n_127_13) );
AOI211_X1 g_108_1 (.ZN (n_108_1), .A (n_112_3), .B (n_118_6), .C1 (n_122_8), .C2 (n_128_11) );
AOI211_X1 g_107_3 (.ZN (n_107_3), .A (n_110_2), .B (n_116_5), .C1 (n_120_7), .C2 (n_126_10) );
AOI211_X1 g_109_4 (.ZN (n_109_4), .A (n_108_1), .B (n_114_4), .C1 (n_118_6), .C2 (n_124_9) );
AOI211_X1 g_111_5 (.ZN (n_111_5), .A (n_107_3), .B (n_112_3), .C1 (n_116_5), .C2 (n_122_8) );
AOI211_X1 g_113_6 (.ZN (n_113_6), .A (n_109_4), .B (n_110_2), .C1 (n_114_4), .C2 (n_120_7) );
AOI211_X1 g_115_7 (.ZN (n_115_7), .A (n_111_5), .B (n_108_1), .C1 (n_112_3), .C2 (n_118_6) );
AOI211_X1 g_117_8 (.ZN (n_117_8), .A (n_113_6), .B (n_107_3), .C1 (n_110_2), .C2 (n_116_5) );
AOI211_X1 g_119_9 (.ZN (n_119_9), .A (n_115_7), .B (n_109_4), .C1 (n_108_1), .C2 (n_114_4) );
AOI211_X1 g_121_10 (.ZN (n_121_10), .A (n_117_8), .B (n_111_5), .C1 (n_107_3), .C2 (n_112_3) );
AOI211_X1 g_123_11 (.ZN (n_123_11), .A (n_119_9), .B (n_113_6), .C1 (n_109_4), .C2 (n_110_2) );
AOI211_X1 g_125_12 (.ZN (n_125_12), .A (n_121_10), .B (n_115_7), .C1 (n_111_5), .C2 (n_108_1) );
AOI211_X1 g_123_13 (.ZN (n_123_13), .A (n_123_11), .B (n_117_8), .C1 (n_113_6), .C2 (n_107_3) );
AOI211_X1 g_124_11 (.ZN (n_124_11), .A (n_125_12), .B (n_119_9), .C1 (n_115_7), .C2 (n_109_4) );
AOI211_X1 g_122_10 (.ZN (n_122_10), .A (n_123_13), .B (n_121_10), .C1 (n_117_8), .C2 (n_111_5) );
AOI211_X1 g_120_9 (.ZN (n_120_9), .A (n_124_11), .B (n_123_11), .C1 (n_119_9), .C2 (n_113_6) );
AOI211_X1 g_118_8 (.ZN (n_118_8), .A (n_122_10), .B (n_125_12), .C1 (n_121_10), .C2 (n_115_7) );
AOI211_X1 g_116_7 (.ZN (n_116_7), .A (n_120_9), .B (n_123_13), .C1 (n_123_11), .C2 (n_117_8) );
AOI211_X1 g_114_6 (.ZN (n_114_6), .A (n_118_8), .B (n_124_11), .C1 (n_125_12), .C2 (n_119_9) );
AOI211_X1 g_112_5 (.ZN (n_112_5), .A (n_116_7), .B (n_122_10), .C1 (n_123_13), .C2 (n_121_10) );
AOI211_X1 g_110_4 (.ZN (n_110_4), .A (n_114_6), .B (n_120_9), .C1 (n_124_11), .C2 (n_123_11) );
AOI211_X1 g_108_3 (.ZN (n_108_3), .A (n_112_5), .B (n_118_8), .C1 (n_122_10), .C2 (n_125_12) );
AOI211_X1 g_106_2 (.ZN (n_106_2), .A (n_110_4), .B (n_116_7), .C1 (n_120_9), .C2 (n_123_13) );
AOI211_X1 g_104_1 (.ZN (n_104_1), .A (n_108_3), .B (n_114_6), .C1 (n_118_8), .C2 (n_124_11) );
AOI211_X1 g_103_3 (.ZN (n_103_3), .A (n_106_2), .B (n_112_5), .C1 (n_116_7), .C2 (n_122_10) );
AOI211_X1 g_105_4 (.ZN (n_105_4), .A (n_104_1), .B (n_110_4), .C1 (n_114_6), .C2 (n_120_9) );
AOI211_X1 g_107_5 (.ZN (n_107_5), .A (n_103_3), .B (n_108_3), .C1 (n_112_5), .C2 (n_118_8) );
AOI211_X1 g_106_3 (.ZN (n_106_3), .A (n_105_4), .B (n_106_2), .C1 (n_110_4), .C2 (n_116_7) );
AOI211_X1 g_105_1 (.ZN (n_105_1), .A (n_107_5), .B (n_104_1), .C1 (n_108_3), .C2 (n_114_6) );
AOI211_X1 g_107_2 (.ZN (n_107_2), .A (n_106_3), .B (n_103_3), .C1 (n_106_2), .C2 (n_112_5) );
AOI211_X1 g_108_4 (.ZN (n_108_4), .A (n_105_1), .B (n_105_4), .C1 (n_104_1), .C2 (n_110_4) );
AOI211_X1 g_109_6 (.ZN (n_109_6), .A (n_107_2), .B (n_107_5), .C1 (n_103_3), .C2 (n_108_3) );
AOI211_X1 g_111_7 (.ZN (n_111_7), .A (n_108_4), .B (n_106_3), .C1 (n_105_4), .C2 (n_106_2) );
AOI211_X1 g_110_5 (.ZN (n_110_5), .A (n_109_6), .B (n_105_1), .C1 (n_107_5), .C2 (n_104_1) );
AOI211_X1 g_109_3 (.ZN (n_109_3), .A (n_111_7), .B (n_107_2), .C1 (n_106_3), .C2 (n_103_3) );
AOI211_X1 g_111_4 (.ZN (n_111_4), .A (n_110_5), .B (n_108_4), .C1 (n_105_1), .C2 (n_105_4) );
AOI211_X1 g_112_6 (.ZN (n_112_6), .A (n_109_3), .B (n_109_6), .C1 (n_107_2), .C2 (n_107_5) );
AOI211_X1 g_113_8 (.ZN (n_113_8), .A (n_111_4), .B (n_111_7), .C1 (n_108_4), .C2 (n_106_3) );
AOI211_X1 g_115_9 (.ZN (n_115_9), .A (n_112_6), .B (n_110_5), .C1 (n_109_6), .C2 (n_105_1) );
AOI211_X1 g_114_7 (.ZN (n_114_7), .A (n_113_8), .B (n_109_3), .C1 (n_111_7), .C2 (n_107_2) );
AOI211_X1 g_113_5 (.ZN (n_113_5), .A (n_115_9), .B (n_111_4), .C1 (n_110_5), .C2 (n_108_4) );
AOI211_X1 g_115_6 (.ZN (n_115_6), .A (n_114_7), .B (n_112_6), .C1 (n_109_3), .C2 (n_109_6) );
AOI211_X1 g_116_8 (.ZN (n_116_8), .A (n_113_5), .B (n_113_8), .C1 (n_111_4), .C2 (n_111_7) );
AOI211_X1 g_117_10 (.ZN (n_117_10), .A (n_115_6), .B (n_115_9), .C1 (n_112_6), .C2 (n_110_5) );
AOI211_X1 g_119_11 (.ZN (n_119_11), .A (n_116_8), .B (n_114_7), .C1 (n_113_8), .C2 (n_109_3) );
AOI211_X1 g_118_9 (.ZN (n_118_9), .A (n_117_10), .B (n_113_5), .C1 (n_115_9), .C2 (n_111_4) );
AOI211_X1 g_117_7 (.ZN (n_117_7), .A (n_119_11), .B (n_115_6), .C1 (n_114_7), .C2 (n_112_6) );
AOI211_X1 g_119_8 (.ZN (n_119_8), .A (n_118_9), .B (n_116_8), .C1 (n_113_5), .C2 (n_113_8) );
AOI211_X1 g_120_10 (.ZN (n_120_10), .A (n_117_7), .B (n_117_10), .C1 (n_115_6), .C2 (n_115_9) );
AOI211_X1 g_121_12 (.ZN (n_121_12), .A (n_119_8), .B (n_119_11), .C1 (n_116_8), .C2 (n_114_7) );
AOI211_X1 g_119_13 (.ZN (n_119_13), .A (n_120_10), .B (n_118_9), .C1 (n_117_10), .C2 (n_113_5) );
AOI211_X1 g_120_11 (.ZN (n_120_11), .A (n_121_12), .B (n_117_7), .C1 (n_119_11), .C2 (n_115_6) );
AOI211_X1 g_121_9 (.ZN (n_121_9), .A (n_119_13), .B (n_119_8), .C1 (n_118_9), .C2 (n_116_8) );
AOI211_X1 g_122_11 (.ZN (n_122_11), .A (n_120_11), .B (n_120_10), .C1 (n_117_7), .C2 (n_117_10) );
AOI211_X1 g_124_12 (.ZN (n_124_12), .A (n_121_9), .B (n_121_12), .C1 (n_119_8), .C2 (n_119_11) );
AOI211_X1 g_123_10 (.ZN (n_123_10), .A (n_122_11), .B (n_119_13), .C1 (n_120_10), .C2 (n_118_9) );
AOI211_X1 g_122_12 (.ZN (n_122_12), .A (n_124_12), .B (n_120_11), .C1 (n_121_12), .C2 (n_117_7) );
AOI211_X1 g_121_14 (.ZN (n_121_14), .A (n_123_10), .B (n_121_9), .C1 (n_119_13), .C2 (n_119_8) );
AOI211_X1 g_120_12 (.ZN (n_120_12), .A (n_122_12), .B (n_122_11), .C1 (n_120_11), .C2 (n_120_10) );
AOI211_X1 g_119_10 (.ZN (n_119_10), .A (n_121_14), .B (n_124_12), .C1 (n_121_9), .C2 (n_121_12) );
AOI211_X1 g_117_9 (.ZN (n_117_9), .A (n_120_12), .B (n_123_10), .C1 (n_122_11), .C2 (n_119_13) );
AOI211_X1 g_118_11 (.ZN (n_118_11), .A (n_119_10), .B (n_122_12), .C1 (n_124_12), .C2 (n_120_11) );
AOI211_X1 g_116_10 (.ZN (n_116_10), .A (n_117_9), .B (n_121_14), .C1 (n_123_10), .C2 (n_121_9) );
AOI211_X1 g_115_8 (.ZN (n_115_8), .A (n_118_11), .B (n_120_12), .C1 (n_122_12), .C2 (n_122_11) );
AOI211_X1 g_113_7 (.ZN (n_113_7), .A (n_116_10), .B (n_119_10), .C1 (n_121_14), .C2 (n_124_12) );
AOI211_X1 g_111_6 (.ZN (n_111_6), .A (n_115_8), .B (n_117_9), .C1 (n_120_12), .C2 (n_123_10) );
AOI211_X1 g_109_5 (.ZN (n_109_5), .A (n_113_7), .B (n_118_11), .C1 (n_119_10), .C2 (n_122_12) );
AOI211_X1 g_107_4 (.ZN (n_107_4), .A (n_111_6), .B (n_116_10), .C1 (n_117_9), .C2 (n_121_14) );
AOI211_X1 g_105_3 (.ZN (n_105_3), .A (n_109_5), .B (n_115_8), .C1 (n_118_11), .C2 (n_120_12) );
AOI211_X1 g_103_2 (.ZN (n_103_2), .A (n_107_4), .B (n_113_7), .C1 (n_116_10), .C2 (n_119_10) );
AOI211_X1 g_101_1 (.ZN (n_101_1), .A (n_105_3), .B (n_111_6), .C1 (n_115_8), .C2 (n_117_9) );
AOI211_X1 g_102_3 (.ZN (n_102_3), .A (n_103_2), .B (n_109_5), .C1 (n_113_7), .C2 (n_118_11) );
AOI211_X1 g_104_4 (.ZN (n_104_4), .A (n_101_1), .B (n_107_4), .C1 (n_111_6), .C2 (n_116_10) );
AOI211_X1 g_106_5 (.ZN (n_106_5), .A (n_102_3), .B (n_105_3), .C1 (n_109_5), .C2 (n_115_8) );
AOI211_X1 g_108_6 (.ZN (n_108_6), .A (n_104_4), .B (n_103_2), .C1 (n_107_4), .C2 (n_113_7) );
AOI211_X1 g_110_7 (.ZN (n_110_7), .A (n_106_5), .B (n_101_1), .C1 (n_105_3), .C2 (n_111_6) );
AOI211_X1 g_112_8 (.ZN (n_112_8), .A (n_108_6), .B (n_102_3), .C1 (n_103_2), .C2 (n_109_5) );
AOI211_X1 g_114_9 (.ZN (n_114_9), .A (n_110_7), .B (n_104_4), .C1 (n_101_1), .C2 (n_107_4) );
AOI211_X1 g_112_10 (.ZN (n_112_10), .A (n_112_8), .B (n_106_5), .C1 (n_102_3), .C2 (n_105_3) );
AOI211_X1 g_111_8 (.ZN (n_111_8), .A (n_114_9), .B (n_108_6), .C1 (n_104_4), .C2 (n_103_2) );
AOI211_X1 g_110_6 (.ZN (n_110_6), .A (n_112_10), .B (n_110_7), .C1 (n_106_5), .C2 (n_101_1) );
AOI211_X1 g_108_5 (.ZN (n_108_5), .A (n_111_8), .B (n_112_8), .C1 (n_108_6), .C2 (n_102_3) );
AOI211_X1 g_106_4 (.ZN (n_106_4), .A (n_110_6), .B (n_114_9), .C1 (n_110_7), .C2 (n_104_4) );
AOI211_X1 g_104_3 (.ZN (n_104_3), .A (n_108_5), .B (n_112_10), .C1 (n_112_8), .C2 (n_106_5) );
AOI211_X1 g_102_2 (.ZN (n_102_2), .A (n_106_4), .B (n_111_8), .C1 (n_114_9), .C2 (n_108_6) );
AOI211_X1 g_100_1 (.ZN (n_100_1), .A (n_104_3), .B (n_110_6), .C1 (n_112_10), .C2 (n_110_7) );
AOI211_X1 g_99_3 (.ZN (n_99_3), .A (n_102_2), .B (n_108_5), .C1 (n_111_8), .C2 (n_112_8) );
AOI211_X1 g_101_4 (.ZN (n_101_4), .A (n_100_1), .B (n_106_4), .C1 (n_110_6), .C2 (n_114_9) );
AOI211_X1 g_103_5 (.ZN (n_103_5), .A (n_99_3), .B (n_104_3), .C1 (n_108_5), .C2 (n_112_10) );
AOI211_X1 g_105_6 (.ZN (n_105_6), .A (n_101_4), .B (n_102_2), .C1 (n_106_4), .C2 (n_111_8) );
AOI211_X1 g_107_7 (.ZN (n_107_7), .A (n_103_5), .B (n_100_1), .C1 (n_104_3), .C2 (n_110_6) );
AOI211_X1 g_109_8 (.ZN (n_109_8), .A (n_105_6), .B (n_99_3), .C1 (n_102_2), .C2 (n_108_5) );
AOI211_X1 g_111_9 (.ZN (n_111_9), .A (n_107_7), .B (n_101_4), .C1 (n_100_1), .C2 (n_106_4) );
AOI211_X1 g_112_7 (.ZN (n_112_7), .A (n_109_8), .B (n_103_5), .C1 (n_99_3), .C2 (n_104_3) );
AOI211_X1 g_113_9 (.ZN (n_113_9), .A (n_111_9), .B (n_105_6), .C1 (n_101_4), .C2 (n_102_2) );
AOI211_X1 g_114_11 (.ZN (n_114_11), .A (n_112_7), .B (n_107_7), .C1 (n_103_5), .C2 (n_100_1) );
AOI211_X1 g_116_12 (.ZN (n_116_12), .A (n_113_9), .B (n_109_8), .C1 (n_105_6), .C2 (n_99_3) );
AOI211_X1 g_115_10 (.ZN (n_115_10), .A (n_114_11), .B (n_111_9), .C1 (n_107_7), .C2 (n_101_4) );
AOI211_X1 g_114_8 (.ZN (n_114_8), .A (n_116_12), .B (n_112_7), .C1 (n_109_8), .C2 (n_103_5) );
AOI211_X1 g_113_10 (.ZN (n_113_10), .A (n_115_10), .B (n_113_9), .C1 (n_111_9), .C2 (n_105_6) );
AOI211_X1 g_115_11 (.ZN (n_115_11), .A (n_114_8), .B (n_114_11), .C1 (n_112_7), .C2 (n_107_7) );
AOI211_X1 g_116_9 (.ZN (n_116_9), .A (n_113_10), .B (n_116_12), .C1 (n_113_9), .C2 (n_109_8) );
AOI211_X1 g_118_10 (.ZN (n_118_10), .A (n_115_11), .B (n_115_10), .C1 (n_114_11), .C2 (n_111_9) );
AOI211_X1 g_117_12 (.ZN (n_117_12), .A (n_116_9), .B (n_114_8), .C1 (n_116_12), .C2 (n_112_7) );
AOI211_X1 g_115_13 (.ZN (n_115_13), .A (n_118_10), .B (n_113_10), .C1 (n_115_10), .C2 (n_113_9) );
AOI211_X1 g_116_11 (.ZN (n_116_11), .A (n_117_12), .B (n_115_11), .C1 (n_114_8), .C2 (n_114_11) );
AOI211_X1 g_114_10 (.ZN (n_114_10), .A (n_115_13), .B (n_116_9), .C1 (n_113_10), .C2 (n_116_12) );
AOI211_X1 g_112_9 (.ZN (n_112_9), .A (n_116_11), .B (n_118_10), .C1 (n_115_11), .C2 (n_115_10) );
AOI211_X1 g_110_8 (.ZN (n_110_8), .A (n_114_10), .B (n_117_12), .C1 (n_116_9), .C2 (n_114_8) );
AOI211_X1 g_108_7 (.ZN (n_108_7), .A (n_112_9), .B (n_115_13), .C1 (n_118_10), .C2 (n_113_10) );
AOI211_X1 g_106_6 (.ZN (n_106_6), .A (n_110_8), .B (n_116_11), .C1 (n_117_12), .C2 (n_115_11) );
AOI211_X1 g_104_5 (.ZN (n_104_5), .A (n_108_7), .B (n_114_10), .C1 (n_115_13), .C2 (n_116_9) );
AOI211_X1 g_102_4 (.ZN (n_102_4), .A (n_106_6), .B (n_112_9), .C1 (n_116_11), .C2 (n_118_10) );
AOI211_X1 g_100_3 (.ZN (n_100_3), .A (n_104_5), .B (n_110_8), .C1 (n_114_10), .C2 (n_117_12) );
AOI211_X1 g_98_2 (.ZN (n_98_2), .A (n_102_4), .B (n_108_7), .C1 (n_112_9), .C2 (n_115_13) );
AOI211_X1 g_96_1 (.ZN (n_96_1), .A (n_100_3), .B (n_106_6), .C1 (n_110_8), .C2 (n_116_11) );
AOI211_X1 g_95_3 (.ZN (n_95_3), .A (n_98_2), .B (n_104_5), .C1 (n_108_7), .C2 (n_114_10) );
AOI211_X1 g_97_4 (.ZN (n_97_4), .A (n_96_1), .B (n_102_4), .C1 (n_106_6), .C2 (n_112_9) );
AOI211_X1 g_99_5 (.ZN (n_99_5), .A (n_95_3), .B (n_100_3), .C1 (n_104_5), .C2 (n_110_8) );
AOI211_X1 g_98_3 (.ZN (n_98_3), .A (n_97_4), .B (n_98_2), .C1 (n_102_4), .C2 (n_108_7) );
AOI211_X1 g_97_1 (.ZN (n_97_1), .A (n_99_5), .B (n_96_1), .C1 (n_100_3), .C2 (n_106_6) );
AOI211_X1 g_99_2 (.ZN (n_99_2), .A (n_98_3), .B (n_95_3), .C1 (n_98_2), .C2 (n_104_5) );
AOI211_X1 g_100_4 (.ZN (n_100_4), .A (n_97_1), .B (n_97_4), .C1 (n_96_1), .C2 (n_102_4) );
AOI211_X1 g_101_6 (.ZN (n_101_6), .A (n_99_2), .B (n_99_5), .C1 (n_95_3), .C2 (n_100_3) );
AOI211_X1 g_103_7 (.ZN (n_103_7), .A (n_100_4), .B (n_98_3), .C1 (n_97_4), .C2 (n_98_2) );
AOI211_X1 g_102_5 (.ZN (n_102_5), .A (n_101_6), .B (n_97_1), .C1 (n_99_5), .C2 (n_96_1) );
AOI211_X1 g_101_3 (.ZN (n_101_3), .A (n_103_7), .B (n_99_2), .C1 (n_98_3), .C2 (n_95_3) );
AOI211_X1 g_103_4 (.ZN (n_103_4), .A (n_102_5), .B (n_100_4), .C1 (n_97_1), .C2 (n_97_4) );
AOI211_X1 g_104_6 (.ZN (n_104_6), .A (n_101_3), .B (n_101_6), .C1 (n_99_2), .C2 (n_99_5) );
AOI211_X1 g_105_8 (.ZN (n_105_8), .A (n_103_4), .B (n_103_7), .C1 (n_100_4), .C2 (n_98_3) );
AOI211_X1 g_107_9 (.ZN (n_107_9), .A (n_104_6), .B (n_102_5), .C1 (n_101_6), .C2 (n_97_1) );
AOI211_X1 g_106_7 (.ZN (n_106_7), .A (n_105_8), .B (n_101_3), .C1 (n_103_7), .C2 (n_99_2) );
AOI211_X1 g_105_5 (.ZN (n_105_5), .A (n_107_9), .B (n_103_4), .C1 (n_102_5), .C2 (n_100_4) );
AOI211_X1 g_107_6 (.ZN (n_107_6), .A (n_106_7), .B (n_104_6), .C1 (n_101_3), .C2 (n_101_6) );
AOI211_X1 g_109_7 (.ZN (n_109_7), .A (n_105_5), .B (n_105_8), .C1 (n_103_4), .C2 (n_103_7) );
AOI211_X1 g_110_9 (.ZN (n_110_9), .A (n_107_6), .B (n_107_9), .C1 (n_104_6), .C2 (n_102_5) );
AOI211_X1 g_108_8 (.ZN (n_108_8), .A (n_109_7), .B (n_106_7), .C1 (n_105_8), .C2 (n_101_3) );
AOI211_X1 g_109_10 (.ZN (n_109_10), .A (n_110_9), .B (n_105_5), .C1 (n_107_9), .C2 (n_103_4) );
AOI211_X1 g_111_11 (.ZN (n_111_11), .A (n_108_8), .B (n_107_6), .C1 (n_106_7), .C2 (n_104_6) );
AOI211_X1 g_113_12 (.ZN (n_113_12), .A (n_109_10), .B (n_109_7), .C1 (n_105_5), .C2 (n_105_8) );
AOI211_X1 g_111_13 (.ZN (n_111_13), .A (n_111_11), .B (n_110_9), .C1 (n_107_6), .C2 (n_107_9) );
AOI211_X1 g_112_11 (.ZN (n_112_11), .A (n_113_12), .B (n_108_8), .C1 (n_109_7), .C2 (n_106_7) );
AOI211_X1 g_110_10 (.ZN (n_110_10), .A (n_111_13), .B (n_109_10), .C1 (n_110_9), .C2 (n_105_5) );
AOI211_X1 g_108_9 (.ZN (n_108_9), .A (n_112_11), .B (n_111_11), .C1 (n_108_8), .C2 (n_107_6) );
AOI211_X1 g_106_8 (.ZN (n_106_8), .A (n_110_10), .B (n_113_12), .C1 (n_109_10), .C2 (n_109_7) );
AOI211_X1 g_104_7 (.ZN (n_104_7), .A (n_108_9), .B (n_111_13), .C1 (n_111_11), .C2 (n_110_9) );
AOI211_X1 g_102_6 (.ZN (n_102_6), .A (n_106_8), .B (n_112_11), .C1 (n_113_12), .C2 (n_108_8) );
AOI211_X1 g_100_5 (.ZN (n_100_5), .A (n_104_7), .B (n_110_10), .C1 (n_111_13), .C2 (n_109_10) );
AOI211_X1 g_98_4 (.ZN (n_98_4), .A (n_102_6), .B (n_108_9), .C1 (n_112_11), .C2 (n_111_11) );
AOI211_X1 g_96_3 (.ZN (n_96_3), .A (n_100_5), .B (n_106_8), .C1 (n_110_10), .C2 (n_113_12) );
AOI211_X1 g_94_2 (.ZN (n_94_2), .A (n_98_4), .B (n_104_7), .C1 (n_108_9), .C2 (n_111_13) );
AOI211_X1 g_92_1 (.ZN (n_92_1), .A (n_96_3), .B (n_102_6), .C1 (n_106_8), .C2 (n_112_11) );
AOI211_X1 g_91_3 (.ZN (n_91_3), .A (n_94_2), .B (n_100_5), .C1 (n_104_7), .C2 (n_110_10) );
AOI211_X1 g_93_4 (.ZN (n_93_4), .A (n_92_1), .B (n_98_4), .C1 (n_102_6), .C2 (n_108_9) );
AOI211_X1 g_95_5 (.ZN (n_95_5), .A (n_91_3), .B (n_96_3), .C1 (n_100_5), .C2 (n_106_8) );
AOI211_X1 g_94_3 (.ZN (n_94_3), .A (n_93_4), .B (n_94_2), .C1 (n_98_4), .C2 (n_104_7) );
AOI211_X1 g_93_1 (.ZN (n_93_1), .A (n_95_5), .B (n_92_1), .C1 (n_96_3), .C2 (n_102_6) );
AOI211_X1 g_95_2 (.ZN (n_95_2), .A (n_94_3), .B (n_91_3), .C1 (n_94_2), .C2 (n_100_5) );
AOI211_X1 g_96_4 (.ZN (n_96_4), .A (n_93_1), .B (n_93_4), .C1 (n_92_1), .C2 (n_98_4) );
AOI211_X1 g_97_6 (.ZN (n_97_6), .A (n_95_2), .B (n_95_5), .C1 (n_91_3), .C2 (n_96_3) );
AOI211_X1 g_99_7 (.ZN (n_99_7), .A (n_96_4), .B (n_94_3), .C1 (n_93_4), .C2 (n_94_2) );
AOI211_X1 g_98_5 (.ZN (n_98_5), .A (n_97_6), .B (n_93_1), .C1 (n_95_5), .C2 (n_92_1) );
AOI211_X1 g_97_3 (.ZN (n_97_3), .A (n_99_7), .B (n_95_2), .C1 (n_94_3), .C2 (n_91_3) );
AOI211_X1 g_99_4 (.ZN (n_99_4), .A (n_98_5), .B (n_96_4), .C1 (n_93_1), .C2 (n_93_4) );
AOI211_X1 g_100_6 (.ZN (n_100_6), .A (n_97_3), .B (n_97_6), .C1 (n_95_2), .C2 (n_95_5) );
AOI211_X1 g_101_8 (.ZN (n_101_8), .A (n_99_4), .B (n_99_7), .C1 (n_96_4), .C2 (n_94_3) );
AOI211_X1 g_103_9 (.ZN (n_103_9), .A (n_100_6), .B (n_98_5), .C1 (n_97_6), .C2 (n_93_1) );
AOI211_X1 g_102_7 (.ZN (n_102_7), .A (n_101_8), .B (n_97_3), .C1 (n_99_7), .C2 (n_95_2) );
AOI211_X1 g_101_5 (.ZN (n_101_5), .A (n_103_9), .B (n_99_4), .C1 (n_98_5), .C2 (n_96_4) );
AOI211_X1 g_103_6 (.ZN (n_103_6), .A (n_102_7), .B (n_100_6), .C1 (n_97_3), .C2 (n_97_6) );
AOI211_X1 g_104_8 (.ZN (n_104_8), .A (n_101_5), .B (n_101_8), .C1 (n_99_4), .C2 (n_99_7) );
AOI211_X1 g_105_10 (.ZN (n_105_10), .A (n_103_6), .B (n_103_9), .C1 (n_100_6), .C2 (n_98_5) );
AOI211_X1 g_107_11 (.ZN (n_107_11), .A (n_104_8), .B (n_102_7), .C1 (n_101_8), .C2 (n_97_3) );
AOI211_X1 g_106_9 (.ZN (n_106_9), .A (n_105_10), .B (n_101_5), .C1 (n_103_9), .C2 (n_99_4) );
AOI211_X1 g_105_7 (.ZN (n_105_7), .A (n_107_11), .B (n_103_6), .C1 (n_102_7), .C2 (n_100_6) );
AOI211_X1 g_107_8 (.ZN (n_107_8), .A (n_106_9), .B (n_104_8), .C1 (n_101_5), .C2 (n_101_8) );
AOI211_X1 g_108_10 (.ZN (n_108_10), .A (n_105_7), .B (n_105_10), .C1 (n_103_6), .C2 (n_103_9) );
AOI211_X1 g_109_12 (.ZN (n_109_12), .A (n_107_8), .B (n_107_11), .C1 (n_104_8), .C2 (n_102_7) );
AOI211_X1 g_107_13 (.ZN (n_107_13), .A (n_108_10), .B (n_106_9), .C1 (n_105_10), .C2 (n_101_5) );
AOI211_X1 g_108_11 (.ZN (n_108_11), .A (n_109_12), .B (n_105_7), .C1 (n_107_11), .C2 (n_103_6) );
AOI211_X1 g_109_9 (.ZN (n_109_9), .A (n_107_13), .B (n_107_8), .C1 (n_106_9), .C2 (n_104_8) );
AOI211_X1 g_110_11 (.ZN (n_110_11), .A (n_108_11), .B (n_108_10), .C1 (n_105_7), .C2 (n_105_10) );
AOI211_X1 g_112_12 (.ZN (n_112_12), .A (n_109_9), .B (n_109_12), .C1 (n_107_8), .C2 (n_107_11) );
AOI211_X1 g_111_10 (.ZN (n_111_10), .A (n_110_11), .B (n_107_13), .C1 (n_108_10), .C2 (n_106_9) );
AOI211_X1 g_110_12 (.ZN (n_110_12), .A (n_112_12), .B (n_108_11), .C1 (n_109_12), .C2 (n_105_7) );
AOI211_X1 g_109_14 (.ZN (n_109_14), .A (n_111_10), .B (n_109_9), .C1 (n_107_13), .C2 (n_107_8) );
AOI211_X1 g_108_12 (.ZN (n_108_12), .A (n_110_12), .B (n_110_11), .C1 (n_108_11), .C2 (n_108_10) );
AOI211_X1 g_107_10 (.ZN (n_107_10), .A (n_109_14), .B (n_112_12), .C1 (n_109_9), .C2 (n_109_12) );
AOI211_X1 g_105_9 (.ZN (n_105_9), .A (n_108_12), .B (n_111_10), .C1 (n_110_11), .C2 (n_107_13) );
AOI211_X1 g_106_11 (.ZN (n_106_11), .A (n_107_10), .B (n_110_12), .C1 (n_112_12), .C2 (n_108_11) );
AOI211_X1 g_104_10 (.ZN (n_104_10), .A (n_105_9), .B (n_109_14), .C1 (n_111_10), .C2 (n_109_9) );
AOI211_X1 g_103_8 (.ZN (n_103_8), .A (n_106_11), .B (n_108_12), .C1 (n_110_12), .C2 (n_110_11) );
AOI211_X1 g_101_7 (.ZN (n_101_7), .A (n_104_10), .B (n_107_10), .C1 (n_109_14), .C2 (n_112_12) );
AOI211_X1 g_99_6 (.ZN (n_99_6), .A (n_103_8), .B (n_105_9), .C1 (n_108_12), .C2 (n_111_10) );
AOI211_X1 g_97_5 (.ZN (n_97_5), .A (n_101_7), .B (n_106_11), .C1 (n_107_10), .C2 (n_110_12) );
AOI211_X1 g_95_4 (.ZN (n_95_4), .A (n_99_6), .B (n_104_10), .C1 (n_105_9), .C2 (n_109_14) );
AOI211_X1 g_93_3 (.ZN (n_93_3), .A (n_97_5), .B (n_103_8), .C1 (n_106_11), .C2 (n_108_12) );
AOI211_X1 g_91_2 (.ZN (n_91_2), .A (n_95_4), .B (n_101_7), .C1 (n_104_10), .C2 (n_107_10) );
AOI211_X1 g_89_1 (.ZN (n_89_1), .A (n_93_3), .B (n_99_6), .C1 (n_103_8), .C2 (n_105_9) );
AOI211_X1 g_90_3 (.ZN (n_90_3), .A (n_91_2), .B (n_97_5), .C1 (n_101_7), .C2 (n_106_11) );
AOI211_X1 g_92_4 (.ZN (n_92_4), .A (n_89_1), .B (n_95_4), .C1 (n_99_6), .C2 (n_104_10) );
AOI211_X1 g_94_5 (.ZN (n_94_5), .A (n_90_3), .B (n_93_3), .C1 (n_97_5), .C2 (n_103_8) );
AOI211_X1 g_96_6 (.ZN (n_96_6), .A (n_92_4), .B (n_91_2), .C1 (n_95_4), .C2 (n_101_7) );
AOI211_X1 g_98_7 (.ZN (n_98_7), .A (n_94_5), .B (n_89_1), .C1 (n_93_3), .C2 (n_99_6) );
AOI211_X1 g_100_8 (.ZN (n_100_8), .A (n_96_6), .B (n_90_3), .C1 (n_91_2), .C2 (n_97_5) );
AOI211_X1 g_102_9 (.ZN (n_102_9), .A (n_98_7), .B (n_92_4), .C1 (n_89_1), .C2 (n_95_4) );
AOI211_X1 g_100_10 (.ZN (n_100_10), .A (n_100_8), .B (n_94_5), .C1 (n_90_3), .C2 (n_93_3) );
AOI211_X1 g_99_8 (.ZN (n_99_8), .A (n_102_9), .B (n_96_6), .C1 (n_92_4), .C2 (n_91_2) );
AOI211_X1 g_98_6 (.ZN (n_98_6), .A (n_100_10), .B (n_98_7), .C1 (n_94_5), .C2 (n_89_1) );
AOI211_X1 g_96_5 (.ZN (n_96_5), .A (n_99_8), .B (n_100_8), .C1 (n_96_6), .C2 (n_90_3) );
AOI211_X1 g_94_4 (.ZN (n_94_4), .A (n_98_6), .B (n_102_9), .C1 (n_98_7), .C2 (n_92_4) );
AOI211_X1 g_92_3 (.ZN (n_92_3), .A (n_96_5), .B (n_100_10), .C1 (n_100_8), .C2 (n_94_5) );
AOI211_X1 g_90_2 (.ZN (n_90_2), .A (n_94_4), .B (n_99_8), .C1 (n_102_9), .C2 (n_96_6) );
AOI211_X1 g_88_1 (.ZN (n_88_1), .A (n_92_3), .B (n_98_6), .C1 (n_100_10), .C2 (n_98_7) );
AOI211_X1 g_87_3 (.ZN (n_87_3), .A (n_90_2), .B (n_96_5), .C1 (n_99_8), .C2 (n_100_8) );
AOI211_X1 g_89_4 (.ZN (n_89_4), .A (n_88_1), .B (n_94_4), .C1 (n_98_6), .C2 (n_102_9) );
AOI211_X1 g_91_5 (.ZN (n_91_5), .A (n_87_3), .B (n_92_3), .C1 (n_96_5), .C2 (n_100_10) );
AOI211_X1 g_93_6 (.ZN (n_93_6), .A (n_89_4), .B (n_90_2), .C1 (n_94_4), .C2 (n_99_8) );
AOI211_X1 g_95_7 (.ZN (n_95_7), .A (n_91_5), .B (n_88_1), .C1 (n_92_3), .C2 (n_98_6) );
AOI211_X1 g_97_8 (.ZN (n_97_8), .A (n_93_6), .B (n_87_3), .C1 (n_90_2), .C2 (n_96_5) );
AOI211_X1 g_99_9 (.ZN (n_99_9), .A (n_95_7), .B (n_89_4), .C1 (n_88_1), .C2 (n_94_4) );
AOI211_X1 g_100_7 (.ZN (n_100_7), .A (n_97_8), .B (n_91_5), .C1 (n_87_3), .C2 (n_92_3) );
AOI211_X1 g_101_9 (.ZN (n_101_9), .A (n_99_9), .B (n_93_6), .C1 (n_89_4), .C2 (n_90_2) );
AOI211_X1 g_102_11 (.ZN (n_102_11), .A (n_100_7), .B (n_95_7), .C1 (n_91_5), .C2 (n_88_1) );
AOI211_X1 g_104_12 (.ZN (n_104_12), .A (n_101_9), .B (n_97_8), .C1 (n_93_6), .C2 (n_87_3) );
AOI211_X1 g_103_10 (.ZN (n_103_10), .A (n_102_11), .B (n_99_9), .C1 (n_95_7), .C2 (n_89_4) );
AOI211_X1 g_102_8 (.ZN (n_102_8), .A (n_104_12), .B (n_100_7), .C1 (n_97_8), .C2 (n_91_5) );
AOI211_X1 g_101_10 (.ZN (n_101_10), .A (n_103_10), .B (n_101_9), .C1 (n_99_9), .C2 (n_93_6) );
AOI211_X1 g_103_11 (.ZN (n_103_11), .A (n_102_8), .B (n_102_11), .C1 (n_100_7), .C2 (n_95_7) );
AOI211_X1 g_104_9 (.ZN (n_104_9), .A (n_101_10), .B (n_104_12), .C1 (n_101_9), .C2 (n_97_8) );
AOI211_X1 g_106_10 (.ZN (n_106_10), .A (n_103_11), .B (n_103_10), .C1 (n_102_11), .C2 (n_99_9) );
AOI211_X1 g_105_12 (.ZN (n_105_12), .A (n_104_9), .B (n_102_8), .C1 (n_104_12), .C2 (n_100_7) );
AOI211_X1 g_103_13 (.ZN (n_103_13), .A (n_106_10), .B (n_101_10), .C1 (n_103_10), .C2 (n_101_9) );
AOI211_X1 g_104_11 (.ZN (n_104_11), .A (n_105_12), .B (n_103_11), .C1 (n_102_8), .C2 (n_102_11) );
AOI211_X1 g_102_10 (.ZN (n_102_10), .A (n_103_13), .B (n_104_9), .C1 (n_101_10), .C2 (n_104_12) );
AOI211_X1 g_100_9 (.ZN (n_100_9), .A (n_104_11), .B (n_106_10), .C1 (n_103_11), .C2 (n_103_10) );
AOI211_X1 g_98_8 (.ZN (n_98_8), .A (n_102_10), .B (n_105_12), .C1 (n_104_9), .C2 (n_102_8) );
AOI211_X1 g_96_7 (.ZN (n_96_7), .A (n_100_9), .B (n_103_13), .C1 (n_106_10), .C2 (n_101_10) );
AOI211_X1 g_94_6 (.ZN (n_94_6), .A (n_98_8), .B (n_104_11), .C1 (n_105_12), .C2 (n_103_11) );
AOI211_X1 g_92_5 (.ZN (n_92_5), .A (n_96_7), .B (n_102_10), .C1 (n_103_13), .C2 (n_104_9) );
AOI211_X1 g_90_4 (.ZN (n_90_4), .A (n_94_6), .B (n_100_9), .C1 (n_104_11), .C2 (n_106_10) );
AOI211_X1 g_88_3 (.ZN (n_88_3), .A (n_92_5), .B (n_98_8), .C1 (n_102_10), .C2 (n_105_12) );
AOI211_X1 g_86_2 (.ZN (n_86_2), .A (n_90_4), .B (n_96_7), .C1 (n_100_9), .C2 (n_103_13) );
AOI211_X1 g_84_1 (.ZN (n_84_1), .A (n_88_3), .B (n_94_6), .C1 (n_98_8), .C2 (n_104_11) );
AOI211_X1 g_83_3 (.ZN (n_83_3), .A (n_86_2), .B (n_92_5), .C1 (n_96_7), .C2 (n_102_10) );
AOI211_X1 g_85_4 (.ZN (n_85_4), .A (n_84_1), .B (n_90_4), .C1 (n_94_6), .C2 (n_100_9) );
AOI211_X1 g_87_5 (.ZN (n_87_5), .A (n_83_3), .B (n_88_3), .C1 (n_92_5), .C2 (n_98_8) );
AOI211_X1 g_86_3 (.ZN (n_86_3), .A (n_85_4), .B (n_86_2), .C1 (n_90_4), .C2 (n_96_7) );
AOI211_X1 g_85_1 (.ZN (n_85_1), .A (n_87_5), .B (n_84_1), .C1 (n_88_3), .C2 (n_94_6) );
AOI211_X1 g_87_2 (.ZN (n_87_2), .A (n_86_3), .B (n_83_3), .C1 (n_86_2), .C2 (n_92_5) );
AOI211_X1 g_88_4 (.ZN (n_88_4), .A (n_85_1), .B (n_85_4), .C1 (n_84_1), .C2 (n_90_4) );
AOI211_X1 g_89_6 (.ZN (n_89_6), .A (n_87_2), .B (n_87_5), .C1 (n_83_3), .C2 (n_88_3) );
AOI211_X1 g_91_7 (.ZN (n_91_7), .A (n_88_4), .B (n_86_3), .C1 (n_85_4), .C2 (n_86_2) );
AOI211_X1 g_90_5 (.ZN (n_90_5), .A (n_89_6), .B (n_85_1), .C1 (n_87_5), .C2 (n_84_1) );
AOI211_X1 g_89_3 (.ZN (n_89_3), .A (n_91_7), .B (n_87_2), .C1 (n_86_3), .C2 (n_83_3) );
AOI211_X1 g_91_4 (.ZN (n_91_4), .A (n_90_5), .B (n_88_4), .C1 (n_85_1), .C2 (n_85_4) );
AOI211_X1 g_92_6 (.ZN (n_92_6), .A (n_89_3), .B (n_89_6), .C1 (n_87_2), .C2 (n_87_5) );
AOI211_X1 g_93_8 (.ZN (n_93_8), .A (n_91_4), .B (n_91_7), .C1 (n_88_4), .C2 (n_86_3) );
AOI211_X1 g_95_9 (.ZN (n_95_9), .A (n_92_6), .B (n_90_5), .C1 (n_89_6), .C2 (n_85_1) );
AOI211_X1 g_94_7 (.ZN (n_94_7), .A (n_93_8), .B (n_89_3), .C1 (n_91_7), .C2 (n_87_2) );
AOI211_X1 g_93_5 (.ZN (n_93_5), .A (n_95_9), .B (n_91_4), .C1 (n_90_5), .C2 (n_88_4) );
AOI211_X1 g_95_6 (.ZN (n_95_6), .A (n_94_7), .B (n_92_6), .C1 (n_89_3), .C2 (n_89_6) );
AOI211_X1 g_97_7 (.ZN (n_97_7), .A (n_93_5), .B (n_93_8), .C1 (n_91_4), .C2 (n_91_7) );
AOI211_X1 g_98_9 (.ZN (n_98_9), .A (n_95_6), .B (n_95_9), .C1 (n_92_6), .C2 (n_90_5) );
AOI211_X1 g_96_8 (.ZN (n_96_8), .A (n_97_7), .B (n_94_7), .C1 (n_93_8), .C2 (n_89_3) );
AOI211_X1 g_97_10 (.ZN (n_97_10), .A (n_98_9), .B (n_93_5), .C1 (n_95_9), .C2 (n_91_4) );
AOI211_X1 g_99_11 (.ZN (n_99_11), .A (n_96_8), .B (n_95_6), .C1 (n_94_7), .C2 (n_92_6) );
AOI211_X1 g_101_12 (.ZN (n_101_12), .A (n_97_10), .B (n_97_7), .C1 (n_93_5), .C2 (n_93_8) );
AOI211_X1 g_99_13 (.ZN (n_99_13), .A (n_99_11), .B (n_98_9), .C1 (n_95_6), .C2 (n_95_9) );
AOI211_X1 g_100_11 (.ZN (n_100_11), .A (n_101_12), .B (n_96_8), .C1 (n_97_7), .C2 (n_94_7) );
AOI211_X1 g_98_10 (.ZN (n_98_10), .A (n_99_13), .B (n_97_10), .C1 (n_98_9), .C2 (n_93_5) );
AOI211_X1 g_96_9 (.ZN (n_96_9), .A (n_100_11), .B (n_99_11), .C1 (n_96_8), .C2 (n_95_6) );
AOI211_X1 g_94_8 (.ZN (n_94_8), .A (n_98_10), .B (n_101_12), .C1 (n_97_10), .C2 (n_97_7) );
AOI211_X1 g_92_7 (.ZN (n_92_7), .A (n_96_9), .B (n_99_13), .C1 (n_99_11), .C2 (n_98_9) );
AOI211_X1 g_90_6 (.ZN (n_90_6), .A (n_94_8), .B (n_100_11), .C1 (n_101_12), .C2 (n_96_8) );
AOI211_X1 g_88_5 (.ZN (n_88_5), .A (n_92_7), .B (n_98_10), .C1 (n_99_13), .C2 (n_97_10) );
AOI211_X1 g_86_4 (.ZN (n_86_4), .A (n_90_6), .B (n_96_9), .C1 (n_100_11), .C2 (n_99_11) );
AOI211_X1 g_84_3 (.ZN (n_84_3), .A (n_88_5), .B (n_94_8), .C1 (n_98_10), .C2 (n_101_12) );
AOI211_X1 g_82_2 (.ZN (n_82_2), .A (n_86_4), .B (n_92_7), .C1 (n_96_9), .C2 (n_99_13) );
AOI211_X1 g_80_1 (.ZN (n_80_1), .A (n_84_3), .B (n_90_6), .C1 (n_94_8), .C2 (n_100_11) );
AOI211_X1 g_79_3 (.ZN (n_79_3), .A (n_82_2), .B (n_88_5), .C1 (n_92_7), .C2 (n_98_10) );
AOI211_X1 g_81_4 (.ZN (n_81_4), .A (n_80_1), .B (n_86_4), .C1 (n_90_6), .C2 (n_96_9) );
AOI211_X1 g_83_5 (.ZN (n_83_5), .A (n_79_3), .B (n_84_3), .C1 (n_88_5), .C2 (n_94_8) );
AOI211_X1 g_82_3 (.ZN (n_82_3), .A (n_81_4), .B (n_82_2), .C1 (n_86_4), .C2 (n_92_7) );
AOI211_X1 g_81_1 (.ZN (n_81_1), .A (n_83_5), .B (n_80_1), .C1 (n_84_3), .C2 (n_90_6) );
AOI211_X1 g_83_2 (.ZN (n_83_2), .A (n_82_3), .B (n_79_3), .C1 (n_82_2), .C2 (n_88_5) );
AOI211_X1 g_84_4 (.ZN (n_84_4), .A (n_81_1), .B (n_81_4), .C1 (n_80_1), .C2 (n_86_4) );
AOI211_X1 g_85_6 (.ZN (n_85_6), .A (n_83_2), .B (n_83_5), .C1 (n_79_3), .C2 (n_84_3) );
AOI211_X1 g_87_7 (.ZN (n_87_7), .A (n_84_4), .B (n_82_3), .C1 (n_81_4), .C2 (n_82_2) );
AOI211_X1 g_86_5 (.ZN (n_86_5), .A (n_85_6), .B (n_81_1), .C1 (n_83_5), .C2 (n_80_1) );
AOI211_X1 g_85_3 (.ZN (n_85_3), .A (n_87_7), .B (n_83_2), .C1 (n_82_3), .C2 (n_79_3) );
AOI211_X1 g_87_4 (.ZN (n_87_4), .A (n_86_5), .B (n_84_4), .C1 (n_81_1), .C2 (n_81_4) );
AOI211_X1 g_88_6 (.ZN (n_88_6), .A (n_85_3), .B (n_85_6), .C1 (n_83_2), .C2 (n_83_5) );
AOI211_X1 g_89_8 (.ZN (n_89_8), .A (n_87_4), .B (n_87_7), .C1 (n_84_4), .C2 (n_82_3) );
AOI211_X1 g_91_9 (.ZN (n_91_9), .A (n_88_6), .B (n_86_5), .C1 (n_85_6), .C2 (n_81_1) );
AOI211_X1 g_90_7 (.ZN (n_90_7), .A (n_89_8), .B (n_85_3), .C1 (n_87_7), .C2 (n_83_2) );
AOI211_X1 g_89_5 (.ZN (n_89_5), .A (n_91_9), .B (n_87_4), .C1 (n_86_5), .C2 (n_84_4) );
AOI211_X1 g_91_6 (.ZN (n_91_6), .A (n_90_7), .B (n_88_6), .C1 (n_85_3), .C2 (n_85_6) );
AOI211_X1 g_92_8 (.ZN (n_92_8), .A (n_89_5), .B (n_89_8), .C1 (n_87_4), .C2 (n_87_7) );
AOI211_X1 g_93_10 (.ZN (n_93_10), .A (n_91_6), .B (n_91_9), .C1 (n_88_6), .C2 (n_86_5) );
AOI211_X1 g_95_11 (.ZN (n_95_11), .A (n_92_8), .B (n_90_7), .C1 (n_89_8), .C2 (n_85_3) );
AOI211_X1 g_94_9 (.ZN (n_94_9), .A (n_93_10), .B (n_89_5), .C1 (n_91_9), .C2 (n_87_4) );
AOI211_X1 g_93_7 (.ZN (n_93_7), .A (n_95_11), .B (n_91_6), .C1 (n_90_7), .C2 (n_88_6) );
AOI211_X1 g_95_8 (.ZN (n_95_8), .A (n_94_9), .B (n_92_8), .C1 (n_89_5), .C2 (n_89_8) );
AOI211_X1 g_96_10 (.ZN (n_96_10), .A (n_93_7), .B (n_93_10), .C1 (n_91_6), .C2 (n_91_9) );
AOI211_X1 g_97_12 (.ZN (n_97_12), .A (n_95_8), .B (n_95_11), .C1 (n_92_8), .C2 (n_90_7) );
AOI211_X1 g_95_13 (.ZN (n_95_13), .A (n_96_10), .B (n_94_9), .C1 (n_93_10), .C2 (n_89_5) );
AOI211_X1 g_96_11 (.ZN (n_96_11), .A (n_97_12), .B (n_93_7), .C1 (n_95_11), .C2 (n_91_6) );
AOI211_X1 g_97_9 (.ZN (n_97_9), .A (n_95_13), .B (n_95_8), .C1 (n_94_9), .C2 (n_92_8) );
AOI211_X1 g_98_11 (.ZN (n_98_11), .A (n_96_11), .B (n_96_10), .C1 (n_93_7), .C2 (n_93_10) );
AOI211_X1 g_100_12 (.ZN (n_100_12), .A (n_97_9), .B (n_97_12), .C1 (n_95_8), .C2 (n_95_11) );
AOI211_X1 g_99_10 (.ZN (n_99_10), .A (n_98_11), .B (n_95_13), .C1 (n_96_10), .C2 (n_94_9) );
AOI211_X1 g_98_12 (.ZN (n_98_12), .A (n_100_12), .B (n_96_11), .C1 (n_97_12), .C2 (n_93_7) );
AOI211_X1 g_97_14 (.ZN (n_97_14), .A (n_99_10), .B (n_97_9), .C1 (n_95_13), .C2 (n_95_8) );
AOI211_X1 g_96_12 (.ZN (n_96_12), .A (n_98_12), .B (n_98_11), .C1 (n_96_11), .C2 (n_96_10) );
AOI211_X1 g_95_10 (.ZN (n_95_10), .A (n_97_14), .B (n_100_12), .C1 (n_97_9), .C2 (n_97_12) );
AOI211_X1 g_93_9 (.ZN (n_93_9), .A (n_96_12), .B (n_99_10), .C1 (n_98_11), .C2 (n_95_13) );
AOI211_X1 g_94_11 (.ZN (n_94_11), .A (n_95_10), .B (n_98_12), .C1 (n_100_12), .C2 (n_96_11) );
AOI211_X1 g_92_10 (.ZN (n_92_10), .A (n_93_9), .B (n_97_14), .C1 (n_99_10), .C2 (n_97_9) );
AOI211_X1 g_91_8 (.ZN (n_91_8), .A (n_94_11), .B (n_96_12), .C1 (n_98_12), .C2 (n_98_11) );
AOI211_X1 g_89_7 (.ZN (n_89_7), .A (n_92_10), .B (n_95_10), .C1 (n_97_14), .C2 (n_100_12) );
AOI211_X1 g_87_6 (.ZN (n_87_6), .A (n_91_8), .B (n_93_9), .C1 (n_96_12), .C2 (n_99_10) );
AOI211_X1 g_85_5 (.ZN (n_85_5), .A (n_89_7), .B (n_94_11), .C1 (n_95_10), .C2 (n_98_12) );
AOI211_X1 g_83_4 (.ZN (n_83_4), .A (n_87_6), .B (n_92_10), .C1 (n_93_9), .C2 (n_97_14) );
AOI211_X1 g_81_3 (.ZN (n_81_3), .A (n_85_5), .B (n_91_8), .C1 (n_94_11), .C2 (n_96_12) );
AOI211_X1 g_79_2 (.ZN (n_79_2), .A (n_83_4), .B (n_89_7), .C1 (n_92_10), .C2 (n_95_10) );
AOI211_X1 g_77_1 (.ZN (n_77_1), .A (n_81_3), .B (n_87_6), .C1 (n_91_8), .C2 (n_93_9) );
AOI211_X1 g_78_3 (.ZN (n_78_3), .A (n_79_2), .B (n_85_5), .C1 (n_89_7), .C2 (n_94_11) );
AOI211_X1 g_80_4 (.ZN (n_80_4), .A (n_77_1), .B (n_83_4), .C1 (n_87_6), .C2 (n_92_10) );
AOI211_X1 g_82_5 (.ZN (n_82_5), .A (n_78_3), .B (n_81_3), .C1 (n_85_5), .C2 (n_91_8) );
AOI211_X1 g_84_6 (.ZN (n_84_6), .A (n_80_4), .B (n_79_2), .C1 (n_83_4), .C2 (n_89_7) );
AOI211_X1 g_86_7 (.ZN (n_86_7), .A (n_82_5), .B (n_77_1), .C1 (n_81_3), .C2 (n_87_6) );
AOI211_X1 g_88_8 (.ZN (n_88_8), .A (n_84_6), .B (n_78_3), .C1 (n_79_2), .C2 (n_85_5) );
AOI211_X1 g_90_9 (.ZN (n_90_9), .A (n_86_7), .B (n_80_4), .C1 (n_77_1), .C2 (n_83_4) );
AOI211_X1 g_88_10 (.ZN (n_88_10), .A (n_88_8), .B (n_82_5), .C1 (n_78_3), .C2 (n_81_3) );
AOI211_X1 g_87_8 (.ZN (n_87_8), .A (n_90_9), .B (n_84_6), .C1 (n_80_4), .C2 (n_79_2) );
AOI211_X1 g_86_6 (.ZN (n_86_6), .A (n_88_10), .B (n_86_7), .C1 (n_82_5), .C2 (n_77_1) );
AOI211_X1 g_84_5 (.ZN (n_84_5), .A (n_87_8), .B (n_88_8), .C1 (n_84_6), .C2 (n_78_3) );
AOI211_X1 g_82_4 (.ZN (n_82_4), .A (n_86_6), .B (n_90_9), .C1 (n_86_7), .C2 (n_80_4) );
AOI211_X1 g_80_3 (.ZN (n_80_3), .A (n_84_5), .B (n_88_10), .C1 (n_88_8), .C2 (n_82_5) );
AOI211_X1 g_78_2 (.ZN (n_78_2), .A (n_82_4), .B (n_87_8), .C1 (n_90_9), .C2 (n_84_6) );
AOI211_X1 g_76_1 (.ZN (n_76_1), .A (n_80_3), .B (n_86_6), .C1 (n_88_10), .C2 (n_86_7) );
AOI211_X1 g_75_3 (.ZN (n_75_3), .A (n_78_2), .B (n_84_5), .C1 (n_87_8), .C2 (n_88_8) );
AOI211_X1 g_77_4 (.ZN (n_77_4), .A (n_76_1), .B (n_82_4), .C1 (n_86_6), .C2 (n_90_9) );
AOI211_X1 g_79_5 (.ZN (n_79_5), .A (n_75_3), .B (n_80_3), .C1 (n_84_5), .C2 (n_88_10) );
AOI211_X1 g_81_6 (.ZN (n_81_6), .A (n_77_4), .B (n_78_2), .C1 (n_82_4), .C2 (n_87_8) );
AOI211_X1 g_83_7 (.ZN (n_83_7), .A (n_79_5), .B (n_76_1), .C1 (n_80_3), .C2 (n_86_6) );
AOI211_X1 g_85_8 (.ZN (n_85_8), .A (n_81_6), .B (n_75_3), .C1 (n_78_2), .C2 (n_84_5) );
AOI211_X1 g_87_9 (.ZN (n_87_9), .A (n_83_7), .B (n_77_4), .C1 (n_76_1), .C2 (n_82_4) );
AOI211_X1 g_88_7 (.ZN (n_88_7), .A (n_85_8), .B (n_79_5), .C1 (n_75_3), .C2 (n_80_3) );
AOI211_X1 g_89_9 (.ZN (n_89_9), .A (n_87_9), .B (n_81_6), .C1 (n_77_4), .C2 (n_78_2) );
AOI211_X1 g_90_11 (.ZN (n_90_11), .A (n_88_7), .B (n_83_7), .C1 (n_79_5), .C2 (n_76_1) );
AOI211_X1 g_92_12 (.ZN (n_92_12), .A (n_89_9), .B (n_85_8), .C1 (n_81_6), .C2 (n_75_3) );
AOI211_X1 g_91_10 (.ZN (n_91_10), .A (n_90_11), .B (n_87_9), .C1 (n_83_7), .C2 (n_77_4) );
AOI211_X1 g_90_8 (.ZN (n_90_8), .A (n_92_12), .B (n_88_7), .C1 (n_85_8), .C2 (n_79_5) );
AOI211_X1 g_89_10 (.ZN (n_89_10), .A (n_91_10), .B (n_89_9), .C1 (n_87_9), .C2 (n_81_6) );
AOI211_X1 g_91_11 (.ZN (n_91_11), .A (n_90_8), .B (n_90_11), .C1 (n_88_7), .C2 (n_83_7) );
AOI211_X1 g_92_9 (.ZN (n_92_9), .A (n_89_10), .B (n_92_12), .C1 (n_89_9), .C2 (n_85_8) );
AOI211_X1 g_94_10 (.ZN (n_94_10), .A (n_91_11), .B (n_91_10), .C1 (n_90_11), .C2 (n_87_9) );
AOI211_X1 g_93_12 (.ZN (n_93_12), .A (n_92_9), .B (n_90_8), .C1 (n_92_12), .C2 (n_88_7) );
AOI211_X1 g_91_13 (.ZN (n_91_13), .A (n_94_10), .B (n_89_10), .C1 (n_91_10), .C2 (n_89_9) );
AOI211_X1 g_92_11 (.ZN (n_92_11), .A (n_93_12), .B (n_91_11), .C1 (n_90_8), .C2 (n_90_11) );
AOI211_X1 g_90_10 (.ZN (n_90_10), .A (n_91_13), .B (n_92_9), .C1 (n_89_10), .C2 (n_92_12) );
AOI211_X1 g_88_9 (.ZN (n_88_9), .A (n_92_11), .B (n_94_10), .C1 (n_91_11), .C2 (n_91_10) );
AOI211_X1 g_86_8 (.ZN (n_86_8), .A (n_90_10), .B (n_93_12), .C1 (n_92_9), .C2 (n_90_8) );
AOI211_X1 g_84_7 (.ZN (n_84_7), .A (n_88_9), .B (n_91_13), .C1 (n_94_10), .C2 (n_89_10) );
AOI211_X1 g_82_6 (.ZN (n_82_6), .A (n_86_8), .B (n_92_11), .C1 (n_93_12), .C2 (n_91_11) );
AOI211_X1 g_80_5 (.ZN (n_80_5), .A (n_84_7), .B (n_90_10), .C1 (n_91_13), .C2 (n_92_9) );
AOI211_X1 g_78_4 (.ZN (n_78_4), .A (n_82_6), .B (n_88_9), .C1 (n_92_11), .C2 (n_94_10) );
AOI211_X1 g_76_3 (.ZN (n_76_3), .A (n_80_5), .B (n_86_8), .C1 (n_90_10), .C2 (n_93_12) );
AOI211_X1 g_74_2 (.ZN (n_74_2), .A (n_78_4), .B (n_84_7), .C1 (n_88_9), .C2 (n_91_13) );
AOI211_X1 g_72_1 (.ZN (n_72_1), .A (n_76_3), .B (n_82_6), .C1 (n_86_8), .C2 (n_92_11) );
AOI211_X1 g_71_3 (.ZN (n_71_3), .A (n_74_2), .B (n_80_5), .C1 (n_84_7), .C2 (n_90_10) );
AOI211_X1 g_73_4 (.ZN (n_73_4), .A (n_72_1), .B (n_78_4), .C1 (n_82_6), .C2 (n_88_9) );
AOI211_X1 g_75_5 (.ZN (n_75_5), .A (n_71_3), .B (n_76_3), .C1 (n_80_5), .C2 (n_86_8) );
AOI211_X1 g_74_3 (.ZN (n_74_3), .A (n_73_4), .B (n_74_2), .C1 (n_78_4), .C2 (n_84_7) );
AOI211_X1 g_73_1 (.ZN (n_73_1), .A (n_75_5), .B (n_72_1), .C1 (n_76_3), .C2 (n_82_6) );
AOI211_X1 g_75_2 (.ZN (n_75_2), .A (n_74_3), .B (n_71_3), .C1 (n_74_2), .C2 (n_80_5) );
AOI211_X1 g_76_4 (.ZN (n_76_4), .A (n_73_1), .B (n_73_4), .C1 (n_72_1), .C2 (n_78_4) );
AOI211_X1 g_77_6 (.ZN (n_77_6), .A (n_75_2), .B (n_75_5), .C1 (n_71_3), .C2 (n_76_3) );
AOI211_X1 g_79_7 (.ZN (n_79_7), .A (n_76_4), .B (n_74_3), .C1 (n_73_4), .C2 (n_74_2) );
AOI211_X1 g_78_5 (.ZN (n_78_5), .A (n_77_6), .B (n_73_1), .C1 (n_75_5), .C2 (n_72_1) );
AOI211_X1 g_77_3 (.ZN (n_77_3), .A (n_79_7), .B (n_75_2), .C1 (n_74_3), .C2 (n_71_3) );
AOI211_X1 g_79_4 (.ZN (n_79_4), .A (n_78_5), .B (n_76_4), .C1 (n_73_1), .C2 (n_73_4) );
AOI211_X1 g_80_6 (.ZN (n_80_6), .A (n_77_3), .B (n_77_6), .C1 (n_75_2), .C2 (n_75_5) );
AOI211_X1 g_81_8 (.ZN (n_81_8), .A (n_79_4), .B (n_79_7), .C1 (n_76_4), .C2 (n_74_3) );
AOI211_X1 g_83_9 (.ZN (n_83_9), .A (n_80_6), .B (n_78_5), .C1 (n_77_6), .C2 (n_73_1) );
AOI211_X1 g_82_7 (.ZN (n_82_7), .A (n_81_8), .B (n_77_3), .C1 (n_79_7), .C2 (n_75_2) );
AOI211_X1 g_81_5 (.ZN (n_81_5), .A (n_83_9), .B (n_79_4), .C1 (n_78_5), .C2 (n_76_4) );
AOI211_X1 g_83_6 (.ZN (n_83_6), .A (n_82_7), .B (n_80_6), .C1 (n_77_3), .C2 (n_77_6) );
AOI211_X1 g_85_7 (.ZN (n_85_7), .A (n_81_5), .B (n_81_8), .C1 (n_79_4), .C2 (n_79_7) );
AOI211_X1 g_86_9 (.ZN (n_86_9), .A (n_83_6), .B (n_83_9), .C1 (n_80_6), .C2 (n_78_5) );
AOI211_X1 g_84_8 (.ZN (n_84_8), .A (n_85_7), .B (n_82_7), .C1 (n_81_8), .C2 (n_77_3) );
AOI211_X1 g_85_10 (.ZN (n_85_10), .A (n_86_9), .B (n_81_5), .C1 (n_83_9), .C2 (n_79_4) );
AOI211_X1 g_87_11 (.ZN (n_87_11), .A (n_84_8), .B (n_83_6), .C1 (n_82_7), .C2 (n_80_6) );
AOI211_X1 g_89_12 (.ZN (n_89_12), .A (n_85_10), .B (n_85_7), .C1 (n_81_5), .C2 (n_81_8) );
AOI211_X1 g_87_13 (.ZN (n_87_13), .A (n_87_11), .B (n_86_9), .C1 (n_83_6), .C2 (n_83_9) );
AOI211_X1 g_88_11 (.ZN (n_88_11), .A (n_89_12), .B (n_84_8), .C1 (n_85_7), .C2 (n_82_7) );
AOI211_X1 g_86_10 (.ZN (n_86_10), .A (n_87_13), .B (n_85_10), .C1 (n_86_9), .C2 (n_81_5) );
AOI211_X1 g_84_9 (.ZN (n_84_9), .A (n_88_11), .B (n_87_11), .C1 (n_84_8), .C2 (n_83_6) );
AOI211_X1 g_82_8 (.ZN (n_82_8), .A (n_86_10), .B (n_89_12), .C1 (n_85_10), .C2 (n_85_7) );
AOI211_X1 g_80_7 (.ZN (n_80_7), .A (n_84_9), .B (n_87_13), .C1 (n_87_11), .C2 (n_86_9) );
AOI211_X1 g_78_6 (.ZN (n_78_6), .A (n_82_8), .B (n_88_11), .C1 (n_89_12), .C2 (n_84_8) );
AOI211_X1 g_76_5 (.ZN (n_76_5), .A (n_80_7), .B (n_86_10), .C1 (n_87_13), .C2 (n_85_10) );
AOI211_X1 g_74_4 (.ZN (n_74_4), .A (n_78_6), .B (n_84_9), .C1 (n_88_11), .C2 (n_87_11) );
AOI211_X1 g_72_3 (.ZN (n_72_3), .A (n_76_5), .B (n_82_8), .C1 (n_86_10), .C2 (n_89_12) );
AOI211_X1 g_70_2 (.ZN (n_70_2), .A (n_74_4), .B (n_80_7), .C1 (n_84_9), .C2 (n_87_13) );
AOI211_X1 g_68_1 (.ZN (n_68_1), .A (n_72_3), .B (n_78_6), .C1 (n_82_8), .C2 (n_88_11) );
AOI211_X1 g_67_3 (.ZN (n_67_3), .A (n_70_2), .B (n_76_5), .C1 (n_80_7), .C2 (n_86_10) );
AOI211_X1 g_69_4 (.ZN (n_69_4), .A (n_68_1), .B (n_74_4), .C1 (n_78_6), .C2 (n_84_9) );
AOI211_X1 g_71_5 (.ZN (n_71_5), .A (n_67_3), .B (n_72_3), .C1 (n_76_5), .C2 (n_82_8) );
AOI211_X1 g_70_3 (.ZN (n_70_3), .A (n_69_4), .B (n_70_2), .C1 (n_74_4), .C2 (n_80_7) );
AOI211_X1 g_69_1 (.ZN (n_69_1), .A (n_71_5), .B (n_68_1), .C1 (n_72_3), .C2 (n_78_6) );
AOI211_X1 g_71_2 (.ZN (n_71_2), .A (n_70_3), .B (n_67_3), .C1 (n_70_2), .C2 (n_76_5) );
AOI211_X1 g_72_4 (.ZN (n_72_4), .A (n_69_1), .B (n_69_4), .C1 (n_68_1), .C2 (n_74_4) );
AOI211_X1 g_73_6 (.ZN (n_73_6), .A (n_71_2), .B (n_71_5), .C1 (n_67_3), .C2 (n_72_3) );
AOI211_X1 g_75_7 (.ZN (n_75_7), .A (n_72_4), .B (n_70_3), .C1 (n_69_4), .C2 (n_70_2) );
AOI211_X1 g_74_5 (.ZN (n_74_5), .A (n_73_6), .B (n_69_1), .C1 (n_71_5), .C2 (n_68_1) );
AOI211_X1 g_73_3 (.ZN (n_73_3), .A (n_75_7), .B (n_71_2), .C1 (n_70_3), .C2 (n_67_3) );
AOI211_X1 g_75_4 (.ZN (n_75_4), .A (n_74_5), .B (n_72_4), .C1 (n_69_1), .C2 (n_69_4) );
AOI211_X1 g_76_6 (.ZN (n_76_6), .A (n_73_3), .B (n_73_6), .C1 (n_71_2), .C2 (n_71_5) );
AOI211_X1 g_77_8 (.ZN (n_77_8), .A (n_75_4), .B (n_75_7), .C1 (n_72_4), .C2 (n_70_3) );
AOI211_X1 g_79_9 (.ZN (n_79_9), .A (n_76_6), .B (n_74_5), .C1 (n_73_6), .C2 (n_69_1) );
AOI211_X1 g_78_7 (.ZN (n_78_7), .A (n_77_8), .B (n_73_3), .C1 (n_75_7), .C2 (n_71_2) );
AOI211_X1 g_77_5 (.ZN (n_77_5), .A (n_79_9), .B (n_75_4), .C1 (n_74_5), .C2 (n_72_4) );
AOI211_X1 g_79_6 (.ZN (n_79_6), .A (n_78_7), .B (n_76_6), .C1 (n_73_3), .C2 (n_73_6) );
AOI211_X1 g_80_8 (.ZN (n_80_8), .A (n_77_5), .B (n_77_8), .C1 (n_75_4), .C2 (n_75_7) );
AOI211_X1 g_81_10 (.ZN (n_81_10), .A (n_79_6), .B (n_79_9), .C1 (n_76_6), .C2 (n_74_5) );
AOI211_X1 g_83_11 (.ZN (n_83_11), .A (n_80_8), .B (n_78_7), .C1 (n_77_8), .C2 (n_73_3) );
AOI211_X1 g_82_9 (.ZN (n_82_9), .A (n_81_10), .B (n_77_5), .C1 (n_79_9), .C2 (n_75_4) );
AOI211_X1 g_81_7 (.ZN (n_81_7), .A (n_83_11), .B (n_79_6), .C1 (n_78_7), .C2 (n_76_6) );
AOI211_X1 g_83_8 (.ZN (n_83_8), .A (n_82_9), .B (n_80_8), .C1 (n_77_5), .C2 (n_77_8) );
AOI211_X1 g_84_10 (.ZN (n_84_10), .A (n_81_7), .B (n_81_10), .C1 (n_79_6), .C2 (n_79_9) );
AOI211_X1 g_85_12 (.ZN (n_85_12), .A (n_83_8), .B (n_83_11), .C1 (n_80_8), .C2 (n_78_7) );
AOI211_X1 g_83_13 (.ZN (n_83_13), .A (n_84_10), .B (n_82_9), .C1 (n_81_10), .C2 (n_77_5) );
AOI211_X1 g_84_11 (.ZN (n_84_11), .A (n_85_12), .B (n_81_7), .C1 (n_83_11), .C2 (n_79_6) );
AOI211_X1 g_85_9 (.ZN (n_85_9), .A (n_83_13), .B (n_83_8), .C1 (n_82_9), .C2 (n_80_8) );
AOI211_X1 g_86_11 (.ZN (n_86_11), .A (n_84_11), .B (n_84_10), .C1 (n_81_7), .C2 (n_81_10) );
AOI211_X1 g_88_12 (.ZN (n_88_12), .A (n_85_9), .B (n_85_12), .C1 (n_83_8), .C2 (n_83_11) );
AOI211_X1 g_87_10 (.ZN (n_87_10), .A (n_86_11), .B (n_83_13), .C1 (n_84_10), .C2 (n_82_9) );
AOI211_X1 g_86_12 (.ZN (n_86_12), .A (n_88_12), .B (n_84_11), .C1 (n_85_12), .C2 (n_81_7) );
AOI211_X1 g_85_14 (.ZN (n_85_14), .A (n_87_10), .B (n_85_9), .C1 (n_83_13), .C2 (n_83_8) );
AOI211_X1 g_84_12 (.ZN (n_84_12), .A (n_86_12), .B (n_86_11), .C1 (n_84_11), .C2 (n_84_10) );
AOI211_X1 g_83_10 (.ZN (n_83_10), .A (n_85_14), .B (n_88_12), .C1 (n_85_9), .C2 (n_85_12) );
AOI211_X1 g_81_9 (.ZN (n_81_9), .A (n_84_12), .B (n_87_10), .C1 (n_86_11), .C2 (n_83_13) );
AOI211_X1 g_82_11 (.ZN (n_82_11), .A (n_83_10), .B (n_86_12), .C1 (n_88_12), .C2 (n_84_11) );
AOI211_X1 g_80_10 (.ZN (n_80_10), .A (n_81_9), .B (n_85_14), .C1 (n_87_10), .C2 (n_85_9) );
AOI211_X1 g_79_8 (.ZN (n_79_8), .A (n_82_11), .B (n_84_12), .C1 (n_86_12), .C2 (n_86_11) );
AOI211_X1 g_77_7 (.ZN (n_77_7), .A (n_80_10), .B (n_83_10), .C1 (n_85_14), .C2 (n_88_12) );
AOI211_X1 g_75_6 (.ZN (n_75_6), .A (n_79_8), .B (n_81_9), .C1 (n_84_12), .C2 (n_87_10) );
AOI211_X1 g_73_5 (.ZN (n_73_5), .A (n_77_7), .B (n_82_11), .C1 (n_83_10), .C2 (n_86_12) );
AOI211_X1 g_71_4 (.ZN (n_71_4), .A (n_75_6), .B (n_80_10), .C1 (n_81_9), .C2 (n_85_14) );
AOI211_X1 g_69_3 (.ZN (n_69_3), .A (n_73_5), .B (n_79_8), .C1 (n_82_11), .C2 (n_84_12) );
AOI211_X1 g_67_2 (.ZN (n_67_2), .A (n_71_4), .B (n_77_7), .C1 (n_80_10), .C2 (n_83_10) );
AOI211_X1 g_65_1 (.ZN (n_65_1), .A (n_69_3), .B (n_75_6), .C1 (n_79_8), .C2 (n_81_9) );
AOI211_X1 g_66_3 (.ZN (n_66_3), .A (n_67_2), .B (n_73_5), .C1 (n_77_7), .C2 (n_82_11) );
AOI211_X1 g_68_4 (.ZN (n_68_4), .A (n_65_1), .B (n_71_4), .C1 (n_75_6), .C2 (n_80_10) );
AOI211_X1 g_70_5 (.ZN (n_70_5), .A (n_66_3), .B (n_69_3), .C1 (n_73_5), .C2 (n_79_8) );
AOI211_X1 g_72_6 (.ZN (n_72_6), .A (n_68_4), .B (n_67_2), .C1 (n_71_4), .C2 (n_77_7) );
AOI211_X1 g_74_7 (.ZN (n_74_7), .A (n_70_5), .B (n_65_1), .C1 (n_69_3), .C2 (n_75_6) );
AOI211_X1 g_76_8 (.ZN (n_76_8), .A (n_72_6), .B (n_66_3), .C1 (n_67_2), .C2 (n_73_5) );
AOI211_X1 g_78_9 (.ZN (n_78_9), .A (n_74_7), .B (n_68_4), .C1 (n_65_1), .C2 (n_71_4) );
AOI211_X1 g_76_10 (.ZN (n_76_10), .A (n_76_8), .B (n_70_5), .C1 (n_66_3), .C2 (n_69_3) );
AOI211_X1 g_75_8 (.ZN (n_75_8), .A (n_78_9), .B (n_72_6), .C1 (n_68_4), .C2 (n_67_2) );
AOI211_X1 g_74_6 (.ZN (n_74_6), .A (n_76_10), .B (n_74_7), .C1 (n_70_5), .C2 (n_65_1) );
AOI211_X1 g_72_5 (.ZN (n_72_5), .A (n_75_8), .B (n_76_8), .C1 (n_72_6), .C2 (n_66_3) );
AOI211_X1 g_70_4 (.ZN (n_70_4), .A (n_74_6), .B (n_78_9), .C1 (n_74_7), .C2 (n_68_4) );
AOI211_X1 g_68_3 (.ZN (n_68_3), .A (n_72_5), .B (n_76_10), .C1 (n_76_8), .C2 (n_70_5) );
AOI211_X1 g_66_2 (.ZN (n_66_2), .A (n_70_4), .B (n_75_8), .C1 (n_78_9), .C2 (n_72_6) );
AOI211_X1 g_64_1 (.ZN (n_64_1), .A (n_68_3), .B (n_74_6), .C1 (n_76_10), .C2 (n_74_7) );
AOI211_X1 g_63_3 (.ZN (n_63_3), .A (n_66_2), .B (n_72_5), .C1 (n_75_8), .C2 (n_76_8) );
AOI211_X1 g_65_4 (.ZN (n_65_4), .A (n_64_1), .B (n_70_4), .C1 (n_74_6), .C2 (n_78_9) );
AOI211_X1 g_67_5 (.ZN (n_67_5), .A (n_63_3), .B (n_68_3), .C1 (n_72_5), .C2 (n_76_10) );
AOI211_X1 g_69_6 (.ZN (n_69_6), .A (n_65_4), .B (n_66_2), .C1 (n_70_4), .C2 (n_75_8) );
AOI211_X1 g_71_7 (.ZN (n_71_7), .A (n_67_5), .B (n_64_1), .C1 (n_68_3), .C2 (n_74_6) );
AOI211_X1 g_73_8 (.ZN (n_73_8), .A (n_69_6), .B (n_63_3), .C1 (n_66_2), .C2 (n_72_5) );
AOI211_X1 g_75_9 (.ZN (n_75_9), .A (n_71_7), .B (n_65_4), .C1 (n_64_1), .C2 (n_70_4) );
AOI211_X1 g_76_7 (.ZN (n_76_7), .A (n_73_8), .B (n_67_5), .C1 (n_63_3), .C2 (n_68_3) );
AOI211_X1 g_77_9 (.ZN (n_77_9), .A (n_75_9), .B (n_69_6), .C1 (n_65_4), .C2 (n_66_2) );
AOI211_X1 g_78_11 (.ZN (n_78_11), .A (n_76_7), .B (n_71_7), .C1 (n_67_5), .C2 (n_64_1) );
AOI211_X1 g_80_12 (.ZN (n_80_12), .A (n_77_9), .B (n_73_8), .C1 (n_69_6), .C2 (n_63_3) );
AOI211_X1 g_79_10 (.ZN (n_79_10), .A (n_78_11), .B (n_75_9), .C1 (n_71_7), .C2 (n_65_4) );
AOI211_X1 g_78_8 (.ZN (n_78_8), .A (n_80_12), .B (n_76_7), .C1 (n_73_8), .C2 (n_67_5) );
AOI211_X1 g_77_10 (.ZN (n_77_10), .A (n_79_10), .B (n_77_9), .C1 (n_75_9), .C2 (n_69_6) );
AOI211_X1 g_79_11 (.ZN (n_79_11), .A (n_78_8), .B (n_78_11), .C1 (n_76_7), .C2 (n_71_7) );
AOI211_X1 g_80_9 (.ZN (n_80_9), .A (n_77_10), .B (n_80_12), .C1 (n_77_9), .C2 (n_73_8) );
AOI211_X1 g_82_10 (.ZN (n_82_10), .A (n_79_11), .B (n_79_10), .C1 (n_78_11), .C2 (n_75_9) );
AOI211_X1 g_81_12 (.ZN (n_81_12), .A (n_80_9), .B (n_78_8), .C1 (n_80_12), .C2 (n_76_7) );
AOI211_X1 g_79_13 (.ZN (n_79_13), .A (n_82_10), .B (n_77_10), .C1 (n_79_10), .C2 (n_77_9) );
AOI211_X1 g_80_11 (.ZN (n_80_11), .A (n_81_12), .B (n_79_11), .C1 (n_78_8), .C2 (n_78_11) );
AOI211_X1 g_78_10 (.ZN (n_78_10), .A (n_79_13), .B (n_80_9), .C1 (n_77_10), .C2 (n_80_12) );
AOI211_X1 g_76_9 (.ZN (n_76_9), .A (n_80_11), .B (n_82_10), .C1 (n_79_11), .C2 (n_79_10) );
AOI211_X1 g_74_8 (.ZN (n_74_8), .A (n_78_10), .B (n_81_12), .C1 (n_80_9), .C2 (n_78_8) );
AOI211_X1 g_72_7 (.ZN (n_72_7), .A (n_76_9), .B (n_79_13), .C1 (n_82_10), .C2 (n_77_10) );
AOI211_X1 g_70_6 (.ZN (n_70_6), .A (n_74_8), .B (n_80_11), .C1 (n_81_12), .C2 (n_79_11) );
AOI211_X1 g_68_5 (.ZN (n_68_5), .A (n_72_7), .B (n_78_10), .C1 (n_79_13), .C2 (n_80_9) );
AOI211_X1 g_66_4 (.ZN (n_66_4), .A (n_70_6), .B (n_76_9), .C1 (n_80_11), .C2 (n_82_10) );
AOI211_X1 g_64_3 (.ZN (n_64_3), .A (n_68_5), .B (n_74_8), .C1 (n_78_10), .C2 (n_81_12) );
AOI211_X1 g_62_2 (.ZN (n_62_2), .A (n_66_4), .B (n_72_7), .C1 (n_76_9), .C2 (n_79_13) );
AOI211_X1 g_60_1 (.ZN (n_60_1), .A (n_64_3), .B (n_70_6), .C1 (n_74_8), .C2 (n_80_11) );
AOI211_X1 g_59_3 (.ZN (n_59_3), .A (n_62_2), .B (n_68_5), .C1 (n_72_7), .C2 (n_78_10) );
AOI211_X1 g_61_4 (.ZN (n_61_4), .A (n_60_1), .B (n_66_4), .C1 (n_70_6), .C2 (n_76_9) );
AOI211_X1 g_63_5 (.ZN (n_63_5), .A (n_59_3), .B (n_64_3), .C1 (n_68_5), .C2 (n_74_8) );
AOI211_X1 g_62_3 (.ZN (n_62_3), .A (n_61_4), .B (n_62_2), .C1 (n_66_4), .C2 (n_72_7) );
AOI211_X1 g_61_1 (.ZN (n_61_1), .A (n_63_5), .B (n_60_1), .C1 (n_64_3), .C2 (n_70_6) );
AOI211_X1 g_63_2 (.ZN (n_63_2), .A (n_62_3), .B (n_59_3), .C1 (n_62_2), .C2 (n_68_5) );
AOI211_X1 g_64_4 (.ZN (n_64_4), .A (n_61_1), .B (n_61_4), .C1 (n_60_1), .C2 (n_66_4) );
AOI211_X1 g_65_6 (.ZN (n_65_6), .A (n_63_2), .B (n_63_5), .C1 (n_59_3), .C2 (n_64_3) );
AOI211_X1 g_67_7 (.ZN (n_67_7), .A (n_64_4), .B (n_62_3), .C1 (n_61_4), .C2 (n_62_2) );
AOI211_X1 g_66_5 (.ZN (n_66_5), .A (n_65_6), .B (n_61_1), .C1 (n_63_5), .C2 (n_60_1) );
AOI211_X1 g_65_3 (.ZN (n_65_3), .A (n_67_7), .B (n_63_2), .C1 (n_62_3), .C2 (n_59_3) );
AOI211_X1 g_67_4 (.ZN (n_67_4), .A (n_66_5), .B (n_64_4), .C1 (n_61_1), .C2 (n_61_4) );
AOI211_X1 g_68_6 (.ZN (n_68_6), .A (n_65_3), .B (n_65_6), .C1 (n_63_2), .C2 (n_63_5) );
AOI211_X1 g_69_8 (.ZN (n_69_8), .A (n_67_4), .B (n_67_7), .C1 (n_64_4), .C2 (n_62_3) );
AOI211_X1 g_71_9 (.ZN (n_71_9), .A (n_68_6), .B (n_66_5), .C1 (n_65_6), .C2 (n_61_1) );
AOI211_X1 g_70_7 (.ZN (n_70_7), .A (n_69_8), .B (n_65_3), .C1 (n_67_7), .C2 (n_63_2) );
AOI211_X1 g_69_5 (.ZN (n_69_5), .A (n_71_9), .B (n_67_4), .C1 (n_66_5), .C2 (n_64_4) );
AOI211_X1 g_71_6 (.ZN (n_71_6), .A (n_70_7), .B (n_68_6), .C1 (n_65_3), .C2 (n_65_6) );
AOI211_X1 g_73_7 (.ZN (n_73_7), .A (n_69_5), .B (n_69_8), .C1 (n_67_4), .C2 (n_67_7) );
AOI211_X1 g_74_9 (.ZN (n_74_9), .A (n_71_6), .B (n_71_9), .C1 (n_68_6), .C2 (n_66_5) );
AOI211_X1 g_72_8 (.ZN (n_72_8), .A (n_73_7), .B (n_70_7), .C1 (n_69_8), .C2 (n_65_3) );
AOI211_X1 g_73_10 (.ZN (n_73_10), .A (n_74_9), .B (n_69_5), .C1 (n_71_9), .C2 (n_67_4) );
AOI211_X1 g_75_11 (.ZN (n_75_11), .A (n_72_8), .B (n_71_6), .C1 (n_70_7), .C2 (n_68_6) );
AOI211_X1 g_77_12 (.ZN (n_77_12), .A (n_73_10), .B (n_73_7), .C1 (n_69_5), .C2 (n_69_8) );
AOI211_X1 g_75_13 (.ZN (n_75_13), .A (n_75_11), .B (n_74_9), .C1 (n_71_6), .C2 (n_71_9) );
AOI211_X1 g_76_11 (.ZN (n_76_11), .A (n_77_12), .B (n_72_8), .C1 (n_73_7), .C2 (n_70_7) );
AOI211_X1 g_74_10 (.ZN (n_74_10), .A (n_75_13), .B (n_73_10), .C1 (n_74_9), .C2 (n_69_5) );
AOI211_X1 g_72_9 (.ZN (n_72_9), .A (n_76_11), .B (n_75_11), .C1 (n_72_8), .C2 (n_71_6) );
AOI211_X1 g_70_8 (.ZN (n_70_8), .A (n_74_10), .B (n_77_12), .C1 (n_73_10), .C2 (n_73_7) );
AOI211_X1 g_68_7 (.ZN (n_68_7), .A (n_72_9), .B (n_75_13), .C1 (n_75_11), .C2 (n_74_9) );
AOI211_X1 g_66_6 (.ZN (n_66_6), .A (n_70_8), .B (n_76_11), .C1 (n_77_12), .C2 (n_72_8) );
AOI211_X1 g_64_5 (.ZN (n_64_5), .A (n_68_7), .B (n_74_10), .C1 (n_75_13), .C2 (n_73_10) );
AOI211_X1 g_62_4 (.ZN (n_62_4), .A (n_66_6), .B (n_72_9), .C1 (n_76_11), .C2 (n_75_11) );
AOI211_X1 g_60_3 (.ZN (n_60_3), .A (n_64_5), .B (n_70_8), .C1 (n_74_10), .C2 (n_77_12) );
AOI211_X1 g_58_2 (.ZN (n_58_2), .A (n_62_4), .B (n_68_7), .C1 (n_72_9), .C2 (n_75_13) );
AOI211_X1 g_56_1 (.ZN (n_56_1), .A (n_60_3), .B (n_66_6), .C1 (n_70_8), .C2 (n_76_11) );
AOI211_X1 g_55_3 (.ZN (n_55_3), .A (n_58_2), .B (n_64_5), .C1 (n_68_7), .C2 (n_74_10) );
AOI211_X1 g_57_4 (.ZN (n_57_4), .A (n_56_1), .B (n_62_4), .C1 (n_66_6), .C2 (n_72_9) );
AOI211_X1 g_59_5 (.ZN (n_59_5), .A (n_55_3), .B (n_60_3), .C1 (n_64_5), .C2 (n_70_8) );
AOI211_X1 g_58_3 (.ZN (n_58_3), .A (n_57_4), .B (n_58_2), .C1 (n_62_4), .C2 (n_68_7) );
AOI211_X1 g_57_1 (.ZN (n_57_1), .A (n_59_5), .B (n_56_1), .C1 (n_60_3), .C2 (n_66_6) );
AOI211_X1 g_59_2 (.ZN (n_59_2), .A (n_58_3), .B (n_55_3), .C1 (n_58_2), .C2 (n_64_5) );
AOI211_X1 g_60_4 (.ZN (n_60_4), .A (n_57_1), .B (n_57_4), .C1 (n_56_1), .C2 (n_62_4) );
AOI211_X1 g_61_6 (.ZN (n_61_6), .A (n_59_2), .B (n_59_5), .C1 (n_55_3), .C2 (n_60_3) );
AOI211_X1 g_63_7 (.ZN (n_63_7), .A (n_60_4), .B (n_58_3), .C1 (n_57_4), .C2 (n_58_2) );
AOI211_X1 g_62_5 (.ZN (n_62_5), .A (n_61_6), .B (n_57_1), .C1 (n_59_5), .C2 (n_56_1) );
AOI211_X1 g_61_3 (.ZN (n_61_3), .A (n_63_7), .B (n_59_2), .C1 (n_58_3), .C2 (n_55_3) );
AOI211_X1 g_63_4 (.ZN (n_63_4), .A (n_62_5), .B (n_60_4), .C1 (n_57_1), .C2 (n_57_4) );
AOI211_X1 g_64_6 (.ZN (n_64_6), .A (n_61_3), .B (n_61_6), .C1 (n_59_2), .C2 (n_59_5) );
AOI211_X1 g_65_8 (.ZN (n_65_8), .A (n_63_4), .B (n_63_7), .C1 (n_60_4), .C2 (n_58_3) );
AOI211_X1 g_67_9 (.ZN (n_67_9), .A (n_64_6), .B (n_62_5), .C1 (n_61_6), .C2 (n_57_1) );
AOI211_X1 g_66_7 (.ZN (n_66_7), .A (n_65_8), .B (n_61_3), .C1 (n_63_7), .C2 (n_59_2) );
AOI211_X1 g_65_5 (.ZN (n_65_5), .A (n_67_9), .B (n_63_4), .C1 (n_62_5), .C2 (n_60_4) );
AOI211_X1 g_67_6 (.ZN (n_67_6), .A (n_66_7), .B (n_64_6), .C1 (n_61_3), .C2 (n_61_6) );
AOI211_X1 g_68_8 (.ZN (n_68_8), .A (n_65_5), .B (n_65_8), .C1 (n_63_4), .C2 (n_63_7) );
AOI211_X1 g_69_10 (.ZN (n_69_10), .A (n_67_6), .B (n_67_9), .C1 (n_64_6), .C2 (n_62_5) );
AOI211_X1 g_71_11 (.ZN (n_71_11), .A (n_68_8), .B (n_66_7), .C1 (n_65_8), .C2 (n_61_3) );
AOI211_X1 g_70_9 (.ZN (n_70_9), .A (n_69_10), .B (n_65_5), .C1 (n_67_9), .C2 (n_63_4) );
AOI211_X1 g_69_7 (.ZN (n_69_7), .A (n_71_11), .B (n_67_6), .C1 (n_66_7), .C2 (n_64_6) );
AOI211_X1 g_71_8 (.ZN (n_71_8), .A (n_70_9), .B (n_68_8), .C1 (n_65_5), .C2 (n_65_8) );
AOI211_X1 g_72_10 (.ZN (n_72_10), .A (n_69_7), .B (n_69_10), .C1 (n_67_6), .C2 (n_67_9) );
AOI211_X1 g_73_12 (.ZN (n_73_12), .A (n_71_8), .B (n_71_11), .C1 (n_68_8), .C2 (n_66_7) );
AOI211_X1 g_71_13 (.ZN (n_71_13), .A (n_72_10), .B (n_70_9), .C1 (n_69_10), .C2 (n_65_5) );
AOI211_X1 g_72_11 (.ZN (n_72_11), .A (n_73_12), .B (n_69_7), .C1 (n_71_11), .C2 (n_67_6) );
AOI211_X1 g_73_9 (.ZN (n_73_9), .A (n_71_13), .B (n_71_8), .C1 (n_70_9), .C2 (n_68_8) );
AOI211_X1 g_74_11 (.ZN (n_74_11), .A (n_72_11), .B (n_72_10), .C1 (n_69_7), .C2 (n_69_10) );
AOI211_X1 g_76_12 (.ZN (n_76_12), .A (n_73_9), .B (n_73_12), .C1 (n_71_8), .C2 (n_71_11) );
AOI211_X1 g_75_10 (.ZN (n_75_10), .A (n_74_11), .B (n_71_13), .C1 (n_72_10), .C2 (n_70_9) );
AOI211_X1 g_74_12 (.ZN (n_74_12), .A (n_76_12), .B (n_72_11), .C1 (n_73_12), .C2 (n_69_7) );
AOI211_X1 g_73_14 (.ZN (n_73_14), .A (n_75_10), .B (n_73_9), .C1 (n_71_13), .C2 (n_71_8) );
AOI211_X1 g_72_12 (.ZN (n_72_12), .A (n_74_12), .B (n_74_11), .C1 (n_72_11), .C2 (n_72_10) );
AOI211_X1 g_71_10 (.ZN (n_71_10), .A (n_73_14), .B (n_76_12), .C1 (n_73_9), .C2 (n_73_12) );
AOI211_X1 g_69_9 (.ZN (n_69_9), .A (n_72_12), .B (n_75_10), .C1 (n_74_11), .C2 (n_71_13) );
AOI211_X1 g_70_11 (.ZN (n_70_11), .A (n_71_10), .B (n_74_12), .C1 (n_76_12), .C2 (n_72_11) );
AOI211_X1 g_68_10 (.ZN (n_68_10), .A (n_69_9), .B (n_73_14), .C1 (n_75_10), .C2 (n_73_9) );
AOI211_X1 g_67_8 (.ZN (n_67_8), .A (n_70_11), .B (n_72_12), .C1 (n_74_12), .C2 (n_74_11) );
AOI211_X1 g_65_7 (.ZN (n_65_7), .A (n_68_10), .B (n_71_10), .C1 (n_73_14), .C2 (n_76_12) );
AOI211_X1 g_63_6 (.ZN (n_63_6), .A (n_67_8), .B (n_69_9), .C1 (n_72_12), .C2 (n_75_10) );
AOI211_X1 g_61_5 (.ZN (n_61_5), .A (n_65_7), .B (n_70_11), .C1 (n_71_10), .C2 (n_74_12) );
AOI211_X1 g_59_4 (.ZN (n_59_4), .A (n_63_6), .B (n_68_10), .C1 (n_69_9), .C2 (n_73_14) );
AOI211_X1 g_57_3 (.ZN (n_57_3), .A (n_61_5), .B (n_67_8), .C1 (n_70_11), .C2 (n_72_12) );
AOI211_X1 g_55_2 (.ZN (n_55_2), .A (n_59_4), .B (n_65_7), .C1 (n_68_10), .C2 (n_71_10) );
AOI211_X1 g_53_1 (.ZN (n_53_1), .A (n_57_3), .B (n_63_6), .C1 (n_67_8), .C2 (n_69_9) );
AOI211_X1 g_54_3 (.ZN (n_54_3), .A (n_55_2), .B (n_61_5), .C1 (n_65_7), .C2 (n_70_11) );
AOI211_X1 g_56_4 (.ZN (n_56_4), .A (n_53_1), .B (n_59_4), .C1 (n_63_6), .C2 (n_68_10) );
AOI211_X1 g_58_5 (.ZN (n_58_5), .A (n_54_3), .B (n_57_3), .C1 (n_61_5), .C2 (n_67_8) );
AOI211_X1 g_60_6 (.ZN (n_60_6), .A (n_56_4), .B (n_55_2), .C1 (n_59_4), .C2 (n_65_7) );
AOI211_X1 g_62_7 (.ZN (n_62_7), .A (n_58_5), .B (n_53_1), .C1 (n_57_3), .C2 (n_63_6) );
AOI211_X1 g_64_8 (.ZN (n_64_8), .A (n_60_6), .B (n_54_3), .C1 (n_55_2), .C2 (n_61_5) );
AOI211_X1 g_66_9 (.ZN (n_66_9), .A (n_62_7), .B (n_56_4), .C1 (n_53_1), .C2 (n_59_4) );
AOI211_X1 g_64_10 (.ZN (n_64_10), .A (n_64_8), .B (n_58_5), .C1 (n_54_3), .C2 (n_57_3) );
AOI211_X1 g_63_8 (.ZN (n_63_8), .A (n_66_9), .B (n_60_6), .C1 (n_56_4), .C2 (n_55_2) );
AOI211_X1 g_62_6 (.ZN (n_62_6), .A (n_64_10), .B (n_62_7), .C1 (n_58_5), .C2 (n_53_1) );
AOI211_X1 g_60_5 (.ZN (n_60_5), .A (n_63_8), .B (n_64_8), .C1 (n_60_6), .C2 (n_54_3) );
AOI211_X1 g_58_4 (.ZN (n_58_4), .A (n_62_6), .B (n_66_9), .C1 (n_62_7), .C2 (n_56_4) );
AOI211_X1 g_56_3 (.ZN (n_56_3), .A (n_60_5), .B (n_64_10), .C1 (n_64_8), .C2 (n_58_5) );
AOI211_X1 g_54_2 (.ZN (n_54_2), .A (n_58_4), .B (n_63_8), .C1 (n_66_9), .C2 (n_60_6) );
AOI211_X1 g_52_1 (.ZN (n_52_1), .A (n_56_3), .B (n_62_6), .C1 (n_64_10), .C2 (n_62_7) );
AOI211_X1 g_50_2 (.ZN (n_50_2), .A (n_54_2), .B (n_60_5), .C1 (n_63_8), .C2 (n_64_8) );
AOI211_X1 g_52_3 (.ZN (n_52_3), .A (n_52_1), .B (n_58_4), .C1 (n_62_6), .C2 (n_66_9) );
AOI211_X1 g_54_4 (.ZN (n_54_4), .A (n_50_2), .B (n_56_3), .C1 (n_60_5), .C2 (n_64_10) );
AOI211_X1 g_56_5 (.ZN (n_56_5), .A (n_52_3), .B (n_54_2), .C1 (n_58_4), .C2 (n_63_8) );
AOI211_X1 g_58_6 (.ZN (n_58_6), .A (n_54_4), .B (n_52_1), .C1 (n_56_3), .C2 (n_62_6) );
AOI211_X1 g_60_7 (.ZN (n_60_7), .A (n_56_5), .B (n_50_2), .C1 (n_54_2), .C2 (n_60_5) );
AOI211_X1 g_61_9 (.ZN (n_61_9), .A (n_58_6), .B (n_52_3), .C1 (n_52_1), .C2 (n_58_4) );
AOI211_X1 g_59_8 (.ZN (n_59_8), .A (n_60_7), .B (n_54_4), .C1 (n_50_2), .C2 (n_56_3) );
AOI211_X1 g_61_7 (.ZN (n_61_7), .A (n_61_9), .B (n_56_5), .C1 (n_52_3), .C2 (n_54_2) );
AOI211_X1 g_59_6 (.ZN (n_59_6), .A (n_59_8), .B (n_58_6), .C1 (n_54_4), .C2 (n_52_1) );
AOI211_X1 g_57_5 (.ZN (n_57_5), .A (n_61_7), .B (n_60_7), .C1 (n_56_5), .C2 (n_50_2) );
AOI211_X1 g_55_4 (.ZN (n_55_4), .A (n_59_6), .B (n_61_9), .C1 (n_58_6), .C2 (n_52_3) );
AOI211_X1 g_53_3 (.ZN (n_53_3), .A (n_57_5), .B (n_59_8), .C1 (n_60_7), .C2 (n_54_4) );
AOI211_X1 g_51_2 (.ZN (n_51_2), .A (n_55_4), .B (n_61_7), .C1 (n_61_9), .C2 (n_56_5) );
AOI211_X1 g_49_1 (.ZN (n_49_1), .A (n_53_3), .B (n_59_6), .C1 (n_59_8), .C2 (n_58_6) );
AOI211_X1 g_47_2 (.ZN (n_47_2), .A (n_51_2), .B (n_57_5), .C1 (n_61_7), .C2 (n_60_7) );
AOI211_X1 g_45_3 (.ZN (n_45_3), .A (n_49_1), .B (n_55_4), .C1 (n_59_6), .C2 (n_61_9) );
AOI211_X1 g_43_4 (.ZN (n_43_4), .A (n_47_2), .B (n_53_3), .C1 (n_57_5), .C2 (n_59_8) );
AOI211_X1 g_41_5 (.ZN (n_41_5), .A (n_45_3), .B (n_51_2), .C1 (n_55_4), .C2 (n_61_7) );
AOI211_X1 g_39_6 (.ZN (n_39_6), .A (n_43_4), .B (n_49_1), .C1 (n_53_3), .C2 (n_59_6) );
AOI211_X1 g_37_7 (.ZN (n_37_7), .A (n_41_5), .B (n_47_2), .C1 (n_51_2), .C2 (n_57_5) );
AOI211_X1 g_35_8 (.ZN (n_35_8), .A (n_39_6), .B (n_45_3), .C1 (n_49_1), .C2 (n_55_4) );
AOI211_X1 g_33_9 (.ZN (n_33_9), .A (n_37_7), .B (n_43_4), .C1 (n_47_2), .C2 (n_53_3) );
AOI211_X1 g_31_10 (.ZN (n_31_10), .A (n_35_8), .B (n_41_5), .C1 (n_45_3), .C2 (n_51_2) );
AOI211_X1 g_29_11 (.ZN (n_29_11), .A (n_33_9), .B (n_39_6), .C1 (n_43_4), .C2 (n_49_1) );
AOI211_X1 g_27_12 (.ZN (n_27_12), .A (n_31_10), .B (n_37_7), .C1 (n_41_5), .C2 (n_47_2) );
AOI211_X1 g_25_13 (.ZN (n_25_13), .A (n_29_11), .B (n_35_8), .C1 (n_39_6), .C2 (n_45_3) );
AOI211_X1 g_23_14 (.ZN (n_23_14), .A (n_27_12), .B (n_33_9), .C1 (n_37_7), .C2 (n_43_4) );
AOI211_X1 g_21_15 (.ZN (n_21_15), .A (n_25_13), .B (n_31_10), .C1 (n_35_8), .C2 (n_41_5) );
AOI211_X1 g_19_16 (.ZN (n_19_16), .A (n_23_14), .B (n_29_11), .C1 (n_33_9), .C2 (n_39_6) );
AOI211_X1 g_17_17 (.ZN (n_17_17), .A (n_21_15), .B (n_27_12), .C1 (n_31_10), .C2 (n_37_7) );
AOI211_X1 g_15_18 (.ZN (n_15_18), .A (n_19_16), .B (n_25_13), .C1 (n_29_11), .C2 (n_35_8) );
AOI211_X1 g_13_19 (.ZN (n_13_19), .A (n_17_17), .B (n_23_14), .C1 (n_27_12), .C2 (n_33_9) );
AOI211_X1 g_11_20 (.ZN (n_11_20), .A (n_15_18), .B (n_21_15), .C1 (n_25_13), .C2 (n_31_10) );
AOI211_X1 g_9_21 (.ZN (n_9_21), .A (n_13_19), .B (n_19_16), .C1 (n_23_14), .C2 (n_29_11) );
AOI211_X1 g_7_22 (.ZN (n_7_22), .A (n_11_20), .B (n_17_17), .C1 (n_21_15), .C2 (n_27_12) );
AOI211_X1 g_8_20 (.ZN (n_8_20), .A (n_9_21), .B (n_15_18), .C1 (n_19_16), .C2 (n_25_13) );
AOI211_X1 g_6_21 (.ZN (n_6_21), .A (n_7_22), .B (n_13_19), .C1 (n_17_17), .C2 (n_23_14) );
AOI211_X1 g_5_23 (.ZN (n_5_23), .A (n_8_20), .B (n_11_20), .C1 (n_15_18), .C2 (n_21_15) );
AOI211_X1 g_3_24 (.ZN (n_3_24), .A (n_6_21), .B (n_9_21), .C1 (n_13_19), .C2 (n_19_16) );
AOI211_X1 g_2_26 (.ZN (n_2_26), .A (n_5_23), .B (n_7_22), .C1 (n_11_20), .C2 (n_17_17) );
AOI211_X1 g_1_28 (.ZN (n_1_28), .A (n_3_24), .B (n_8_20), .C1 (n_9_21), .C2 (n_15_18) );
AOI211_X1 g_3_27 (.ZN (n_3_27), .A (n_2_26), .B (n_6_21), .C1 (n_7_22), .C2 (n_13_19) );
AOI211_X1 g_4_25 (.ZN (n_4_25), .A (n_1_28), .B (n_5_23), .C1 (n_8_20), .C2 (n_11_20) );
AOI211_X1 g_6_24 (.ZN (n_6_24), .A (n_3_27), .B (n_3_24), .C1 (n_6_21), .C2 (n_9_21) );
AOI211_X1 g_4_23 (.ZN (n_4_23), .A (n_4_25), .B (n_2_26), .C1 (n_5_23), .C2 (n_7_22) );
AOI211_X1 g_3_25 (.ZN (n_3_25), .A (n_6_24), .B (n_1_28), .C1 (n_3_24), .C2 (n_8_20) );
AOI211_X1 g_5_26 (.ZN (n_5_26), .A (n_4_23), .B (n_3_27), .C1 (n_2_26), .C2 (n_6_21) );
AOI211_X1 g_7_25 (.ZN (n_7_25), .A (n_3_25), .B (n_4_25), .C1 (n_1_28), .C2 (n_5_23) );
AOI211_X1 g_6_23 (.ZN (n_6_23), .A (n_5_26), .B (n_6_24), .C1 (n_3_27), .C2 (n_3_24) );
AOI211_X1 g_8_22 (.ZN (n_8_22), .A (n_7_25), .B (n_4_23), .C1 (n_4_25), .C2 (n_2_26) );
AOI211_X1 g_10_21 (.ZN (n_10_21), .A (n_6_23), .B (n_3_25), .C1 (n_6_24), .C2 (n_1_28) );
AOI211_X1 g_12_20 (.ZN (n_12_20), .A (n_8_22), .B (n_5_26), .C1 (n_4_23), .C2 (n_3_27) );
AOI211_X1 g_14_19 (.ZN (n_14_19), .A (n_10_21), .B (n_7_25), .C1 (n_3_25), .C2 (n_4_25) );
AOI211_X1 g_16_18 (.ZN (n_16_18), .A (n_12_20), .B (n_6_23), .C1 (n_5_26), .C2 (n_6_24) );
AOI211_X1 g_18_17 (.ZN (n_18_17), .A (n_14_19), .B (n_8_22), .C1 (n_7_25), .C2 (n_4_23) );
AOI211_X1 g_20_16 (.ZN (n_20_16), .A (n_16_18), .B (n_10_21), .C1 (n_6_23), .C2 (n_3_25) );
AOI211_X1 g_22_15 (.ZN (n_22_15), .A (n_18_17), .B (n_12_20), .C1 (n_8_22), .C2 (n_5_26) );
AOI211_X1 g_24_14 (.ZN (n_24_14), .A (n_20_16), .B (n_14_19), .C1 (n_10_21), .C2 (n_7_25) );
AOI211_X1 g_26_13 (.ZN (n_26_13), .A (n_22_15), .B (n_16_18), .C1 (n_12_20), .C2 (n_6_23) );
AOI211_X1 g_25_15 (.ZN (n_25_15), .A (n_24_14), .B (n_18_17), .C1 (n_14_19), .C2 (n_8_22) );
AOI211_X1 g_27_14 (.ZN (n_27_14), .A (n_26_13), .B (n_20_16), .C1 (n_16_18), .C2 (n_10_21) );
AOI211_X1 g_29_13 (.ZN (n_29_13), .A (n_25_15), .B (n_22_15), .C1 (n_18_17), .C2 (n_12_20) );
AOI211_X1 g_31_12 (.ZN (n_31_12), .A (n_27_14), .B (n_24_14), .C1 (n_20_16), .C2 (n_14_19) );
AOI211_X1 g_33_11 (.ZN (n_33_11), .A (n_29_13), .B (n_26_13), .C1 (n_22_15), .C2 (n_16_18) );
AOI211_X1 g_35_10 (.ZN (n_35_10), .A (n_31_12), .B (n_25_15), .C1 (n_24_14), .C2 (n_18_17) );
AOI211_X1 g_37_9 (.ZN (n_37_9), .A (n_33_11), .B (n_27_14), .C1 (n_26_13), .C2 (n_20_16) );
AOI211_X1 g_39_8 (.ZN (n_39_8), .A (n_35_10), .B (n_29_13), .C1 (n_25_15), .C2 (n_22_15) );
AOI211_X1 g_41_7 (.ZN (n_41_7), .A (n_37_9), .B (n_31_12), .C1 (n_27_14), .C2 (n_24_14) );
AOI211_X1 g_43_6 (.ZN (n_43_6), .A (n_39_8), .B (n_33_11), .C1 (n_29_13), .C2 (n_26_13) );
AOI211_X1 g_45_5 (.ZN (n_45_5), .A (n_41_7), .B (n_35_10), .C1 (n_31_12), .C2 (n_25_15) );
AOI211_X1 g_47_4 (.ZN (n_47_4), .A (n_43_6), .B (n_37_9), .C1 (n_33_11), .C2 (n_27_14) );
AOI211_X1 g_49_3 (.ZN (n_49_3), .A (n_45_5), .B (n_39_8), .C1 (n_35_10), .C2 (n_29_13) );
AOI211_X1 g_51_4 (.ZN (n_51_4), .A (n_47_4), .B (n_41_7), .C1 (n_37_9), .C2 (n_31_12) );
AOI211_X1 g_53_5 (.ZN (n_53_5), .A (n_49_3), .B (n_43_6), .C1 (n_39_8), .C2 (n_33_11) );
AOI211_X1 g_55_6 (.ZN (n_55_6), .A (n_51_4), .B (n_45_5), .C1 (n_41_7), .C2 (n_35_10) );
AOI211_X1 g_57_7 (.ZN (n_57_7), .A (n_53_5), .B (n_47_4), .C1 (n_43_6), .C2 (n_37_9) );
AOI211_X1 g_55_8 (.ZN (n_55_8), .A (n_55_6), .B (n_49_3), .C1 (n_45_5), .C2 (n_39_8) );
AOI211_X1 g_56_6 (.ZN (n_56_6), .A (n_57_7), .B (n_51_4), .C1 (n_47_4), .C2 (n_41_7) );
AOI211_X1 g_54_5 (.ZN (n_54_5), .A (n_55_8), .B (n_53_5), .C1 (n_49_3), .C2 (n_43_6) );
AOI211_X1 g_52_4 (.ZN (n_52_4), .A (n_56_6), .B (n_55_6), .C1 (n_51_4), .C2 (n_45_5) );
AOI211_X1 g_50_3 (.ZN (n_50_3), .A (n_54_5), .B (n_57_7), .C1 (n_53_5), .C2 (n_47_4) );
AOI211_X1 g_48_4 (.ZN (n_48_4), .A (n_52_4), .B (n_55_8), .C1 (n_55_6), .C2 (n_49_3) );
AOI211_X1 g_46_5 (.ZN (n_46_5), .A (n_50_3), .B (n_56_6), .C1 (n_57_7), .C2 (n_51_4) );
AOI211_X1 g_44_6 (.ZN (n_44_6), .A (n_48_4), .B (n_54_5), .C1 (n_55_8), .C2 (n_53_5) );
AOI211_X1 g_42_7 (.ZN (n_42_7), .A (n_46_5), .B (n_52_4), .C1 (n_56_6), .C2 (n_55_6) );
AOI211_X1 g_40_8 (.ZN (n_40_8), .A (n_44_6), .B (n_50_3), .C1 (n_54_5), .C2 (n_57_7) );
AOI211_X1 g_38_9 (.ZN (n_38_9), .A (n_42_7), .B (n_48_4), .C1 (n_52_4), .C2 (n_55_8) );
AOI211_X1 g_36_10 (.ZN (n_36_10), .A (n_40_8), .B (n_46_5), .C1 (n_50_3), .C2 (n_56_6) );
AOI211_X1 g_34_11 (.ZN (n_34_11), .A (n_38_9), .B (n_44_6), .C1 (n_48_4), .C2 (n_54_5) );
AOI211_X1 g_32_12 (.ZN (n_32_12), .A (n_36_10), .B (n_42_7), .C1 (n_46_5), .C2 (n_52_4) );
AOI211_X1 g_30_13 (.ZN (n_30_13), .A (n_34_11), .B (n_40_8), .C1 (n_44_6), .C2 (n_50_3) );
AOI211_X1 g_28_14 (.ZN (n_28_14), .A (n_32_12), .B (n_38_9), .C1 (n_42_7), .C2 (n_48_4) );
AOI211_X1 g_26_15 (.ZN (n_26_15), .A (n_30_13), .B (n_36_10), .C1 (n_40_8), .C2 (n_46_5) );
AOI211_X1 g_27_13 (.ZN (n_27_13), .A (n_28_14), .B (n_34_11), .C1 (n_38_9), .C2 (n_44_6) );
AOI211_X1 g_25_14 (.ZN (n_25_14), .A (n_26_15), .B (n_32_12), .C1 (n_36_10), .C2 (n_42_7) );
AOI211_X1 g_23_15 (.ZN (n_23_15), .A (n_27_13), .B (n_30_13), .C1 (n_34_11), .C2 (n_40_8) );
AOI211_X1 g_21_16 (.ZN (n_21_16), .A (n_25_14), .B (n_28_14), .C1 (n_32_12), .C2 (n_38_9) );
AOI211_X1 g_19_17 (.ZN (n_19_17), .A (n_23_15), .B (n_26_15), .C1 (n_30_13), .C2 (n_36_10) );
AOI211_X1 g_17_18 (.ZN (n_17_18), .A (n_21_16), .B (n_27_13), .C1 (n_28_14), .C2 (n_34_11) );
AOI211_X1 g_15_19 (.ZN (n_15_19), .A (n_19_17), .B (n_25_14), .C1 (n_26_15), .C2 (n_32_12) );
AOI211_X1 g_13_20 (.ZN (n_13_20), .A (n_17_18), .B (n_23_15), .C1 (n_27_13), .C2 (n_30_13) );
AOI211_X1 g_11_21 (.ZN (n_11_21), .A (n_15_19), .B (n_21_16), .C1 (n_25_14), .C2 (n_28_14) );
AOI211_X1 g_9_22 (.ZN (n_9_22), .A (n_13_20), .B (n_19_17), .C1 (n_23_15), .C2 (n_26_15) );
AOI211_X1 g_10_20 (.ZN (n_10_20), .A (n_11_21), .B (n_17_18), .C1 (n_21_16), .C2 (n_27_13) );
AOI211_X1 g_8_21 (.ZN (n_8_21), .A (n_9_22), .B (n_15_19), .C1 (n_19_17), .C2 (n_25_14) );
AOI211_X1 g_6_22 (.ZN (n_6_22), .A (n_10_20), .B (n_13_20), .C1 (n_17_18), .C2 (n_23_15) );
AOI211_X1 g_5_24 (.ZN (n_5_24), .A (n_8_21), .B (n_11_21), .C1 (n_15_19), .C2 (n_21_16) );
AOI211_X1 g_7_23 (.ZN (n_7_23), .A (n_6_22), .B (n_9_22), .C1 (n_13_20), .C2 (n_19_17) );
AOI211_X1 g_6_25 (.ZN (n_6_25), .A (n_5_24), .B (n_10_20), .C1 (n_11_21), .C2 (n_17_18) );
AOI211_X1 g_4_26 (.ZN (n_4_26), .A (n_7_23), .B (n_8_21), .C1 (n_9_22), .C2 (n_15_19) );
AOI211_X1 g_3_28 (.ZN (n_3_28), .A (n_6_25), .B (n_6_22), .C1 (n_10_20), .C2 (n_13_20) );
AOI211_X1 g_5_27 (.ZN (n_5_27), .A (n_4_26), .B (n_5_24), .C1 (n_8_21), .C2 (n_11_21) );
AOI211_X1 g_4_29 (.ZN (n_4_29), .A (n_3_28), .B (n_7_23), .C1 (n_6_22), .C2 (n_9_22) );
AOI211_X1 g_2_30 (.ZN (n_2_30), .A (n_5_27), .B (n_6_25), .C1 (n_5_24), .C2 (n_10_20) );
AOI211_X1 g_1_32 (.ZN (n_1_32), .A (n_4_29), .B (n_4_26), .C1 (n_7_23), .C2 (n_8_21) );
AOI211_X1 g_3_31 (.ZN (n_3_31), .A (n_2_30), .B (n_3_28), .C1 (n_6_25), .C2 (n_6_22) );
AOI211_X1 g_5_30 (.ZN (n_5_30), .A (n_1_32), .B (n_5_27), .C1 (n_4_26), .C2 (n_5_24) );
AOI211_X1 g_3_29 (.ZN (n_3_29), .A (n_3_31), .B (n_4_29), .C1 (n_3_28), .C2 (n_7_23) );
AOI211_X1 g_4_27 (.ZN (n_4_27), .A (n_5_30), .B (n_2_30), .C1 (n_5_27), .C2 (n_6_25) );
AOI211_X1 g_5_25 (.ZN (n_5_25), .A (n_3_29), .B (n_1_32), .C1 (n_4_29), .C2 (n_4_26) );
AOI211_X1 g_7_24 (.ZN (n_7_24), .A (n_4_27), .B (n_3_31), .C1 (n_2_30), .C2 (n_3_28) );
AOI211_X1 g_9_23 (.ZN (n_9_23), .A (n_5_25), .B (n_5_30), .C1 (n_1_32), .C2 (n_5_27) );
AOI211_X1 g_11_22 (.ZN (n_11_22), .A (n_7_24), .B (n_3_29), .C1 (n_3_31), .C2 (n_4_29) );
AOI211_X1 g_13_21 (.ZN (n_13_21), .A (n_9_23), .B (n_4_27), .C1 (n_5_30), .C2 (n_2_30) );
AOI211_X1 g_15_20 (.ZN (n_15_20), .A (n_11_22), .B (n_5_25), .C1 (n_3_29), .C2 (n_1_32) );
AOI211_X1 g_17_19 (.ZN (n_17_19), .A (n_13_21), .B (n_7_24), .C1 (n_4_27), .C2 (n_3_31) );
AOI211_X1 g_19_18 (.ZN (n_19_18), .A (n_15_20), .B (n_9_23), .C1 (n_5_25), .C2 (n_5_30) );
AOI211_X1 g_21_17 (.ZN (n_21_17), .A (n_17_19), .B (n_11_22), .C1 (n_7_24), .C2 (n_3_29) );
AOI211_X1 g_23_16 (.ZN (n_23_16), .A (n_19_18), .B (n_13_21), .C1 (n_9_23), .C2 (n_4_27) );
AOI211_X1 g_22_18 (.ZN (n_22_18), .A (n_21_17), .B (n_15_20), .C1 (n_11_22), .C2 (n_5_25) );
AOI211_X1 g_20_17 (.ZN (n_20_17), .A (n_23_16), .B (n_17_19), .C1 (n_13_21), .C2 (n_7_24) );
AOI211_X1 g_22_16 (.ZN (n_22_16), .A (n_22_18), .B (n_19_18), .C1 (n_15_20), .C2 (n_9_23) );
AOI211_X1 g_24_15 (.ZN (n_24_15), .A (n_20_17), .B (n_21_17), .C1 (n_17_19), .C2 (n_11_22) );
AOI211_X1 g_26_14 (.ZN (n_26_14), .A (n_22_16), .B (n_23_16), .C1 (n_19_18), .C2 (n_13_21) );
AOI211_X1 g_28_13 (.ZN (n_28_13), .A (n_24_15), .B (n_22_18), .C1 (n_21_17), .C2 (n_15_20) );
AOI211_X1 g_30_12 (.ZN (n_30_12), .A (n_26_14), .B (n_20_17), .C1 (n_23_16), .C2 (n_17_19) );
AOI211_X1 g_32_11 (.ZN (n_32_11), .A (n_28_13), .B (n_22_16), .C1 (n_22_18), .C2 (n_19_18) );
AOI211_X1 g_34_10 (.ZN (n_34_10), .A (n_30_12), .B (n_24_15), .C1 (n_20_17), .C2 (n_21_17) );
AOI211_X1 g_36_9 (.ZN (n_36_9), .A (n_32_11), .B (n_26_14), .C1 (n_22_16), .C2 (n_23_16) );
AOI211_X1 g_38_8 (.ZN (n_38_8), .A (n_34_10), .B (n_28_13), .C1 (n_24_15), .C2 (n_22_18) );
AOI211_X1 g_40_7 (.ZN (n_40_7), .A (n_36_9), .B (n_30_12), .C1 (n_26_14), .C2 (n_20_17) );
AOI211_X1 g_42_6 (.ZN (n_42_6), .A (n_38_8), .B (n_32_11), .C1 (n_28_13), .C2 (n_22_16) );
AOI211_X1 g_44_5 (.ZN (n_44_5), .A (n_40_7), .B (n_34_10), .C1 (n_30_12), .C2 (n_24_15) );
AOI211_X1 g_46_4 (.ZN (n_46_4), .A (n_42_6), .B (n_36_9), .C1 (n_32_11), .C2 (n_26_14) );
AOI211_X1 g_48_3 (.ZN (n_48_3), .A (n_44_5), .B (n_38_8), .C1 (n_34_10), .C2 (n_28_13) );
AOI211_X1 g_49_5 (.ZN (n_49_5), .A (n_46_4), .B (n_40_7), .C1 (n_36_9), .C2 (n_30_12) );
AOI211_X1 g_47_6 (.ZN (n_47_6), .A (n_48_3), .B (n_42_6), .C1 (n_38_8), .C2 (n_32_11) );
AOI211_X1 g_45_7 (.ZN (n_45_7), .A (n_49_5), .B (n_44_5), .C1 (n_40_7), .C2 (n_34_10) );
AOI211_X1 g_43_8 (.ZN (n_43_8), .A (n_47_6), .B (n_46_4), .C1 (n_42_6), .C2 (n_36_9) );
AOI211_X1 g_41_9 (.ZN (n_41_9), .A (n_45_7), .B (n_48_3), .C1 (n_44_5), .C2 (n_38_8) );
AOI211_X1 g_39_10 (.ZN (n_39_10), .A (n_43_8), .B (n_49_5), .C1 (n_46_4), .C2 (n_40_7) );
AOI211_X1 g_37_11 (.ZN (n_37_11), .A (n_41_9), .B (n_47_6), .C1 (n_48_3), .C2 (n_42_6) );
AOI211_X1 g_35_12 (.ZN (n_35_12), .A (n_39_10), .B (n_45_7), .C1 (n_49_5), .C2 (n_44_5) );
AOI211_X1 g_33_13 (.ZN (n_33_13), .A (n_37_11), .B (n_43_8), .C1 (n_47_6), .C2 (n_46_4) );
AOI211_X1 g_31_14 (.ZN (n_31_14), .A (n_35_12), .B (n_41_9), .C1 (n_45_7), .C2 (n_48_3) );
AOI211_X1 g_29_15 (.ZN (n_29_15), .A (n_33_13), .B (n_39_10), .C1 (n_43_8), .C2 (n_49_5) );
AOI211_X1 g_27_16 (.ZN (n_27_16), .A (n_31_14), .B (n_37_11), .C1 (n_41_9), .C2 (n_47_6) );
AOI211_X1 g_25_17 (.ZN (n_25_17), .A (n_29_15), .B (n_35_12), .C1 (n_39_10), .C2 (n_45_7) );
AOI211_X1 g_23_18 (.ZN (n_23_18), .A (n_27_16), .B (n_33_13), .C1 (n_37_11), .C2 (n_43_8) );
AOI211_X1 g_24_16 (.ZN (n_24_16), .A (n_25_17), .B (n_31_14), .C1 (n_35_12), .C2 (n_41_9) );
AOI211_X1 g_22_17 (.ZN (n_22_17), .A (n_23_18), .B (n_29_15), .C1 (n_33_13), .C2 (n_39_10) );
AOI211_X1 g_20_18 (.ZN (n_20_18), .A (n_24_16), .B (n_27_16), .C1 (n_31_14), .C2 (n_37_11) );
AOI211_X1 g_18_19 (.ZN (n_18_19), .A (n_22_17), .B (n_25_17), .C1 (n_29_15), .C2 (n_35_12) );
AOI211_X1 g_16_20 (.ZN (n_16_20), .A (n_20_18), .B (n_23_18), .C1 (n_27_16), .C2 (n_33_13) );
AOI211_X1 g_14_21 (.ZN (n_14_21), .A (n_18_19), .B (n_24_16), .C1 (n_25_17), .C2 (n_31_14) );
AOI211_X1 g_12_22 (.ZN (n_12_22), .A (n_16_20), .B (n_22_17), .C1 (n_23_18), .C2 (n_29_15) );
AOI211_X1 g_10_23 (.ZN (n_10_23), .A (n_14_21), .B (n_20_18), .C1 (n_24_16), .C2 (n_27_16) );
AOI211_X1 g_8_24 (.ZN (n_8_24), .A (n_12_22), .B (n_18_19), .C1 (n_22_17), .C2 (n_25_17) );
AOI211_X1 g_7_26 (.ZN (n_7_26), .A (n_10_23), .B (n_16_20), .C1 (n_20_18), .C2 (n_23_18) );
AOI211_X1 g_6_28 (.ZN (n_6_28), .A (n_8_24), .B (n_14_21), .C1 (n_18_19), .C2 (n_24_16) );
AOI211_X1 g_8_27 (.ZN (n_8_27), .A (n_7_26), .B (n_12_22), .C1 (n_16_20), .C2 (n_22_17) );
AOI211_X1 g_6_26 (.ZN (n_6_26), .A (n_6_28), .B (n_10_23), .C1 (n_14_21), .C2 (n_20_18) );
AOI211_X1 g_8_25 (.ZN (n_8_25), .A (n_8_27), .B (n_8_24), .C1 (n_12_22), .C2 (n_18_19) );
AOI211_X1 g_10_24 (.ZN (n_10_24), .A (n_6_26), .B (n_7_26), .C1 (n_10_23), .C2 (n_16_20) );
AOI211_X1 g_8_23 (.ZN (n_8_23), .A (n_8_25), .B (n_6_28), .C1 (n_8_24), .C2 (n_14_21) );
AOI211_X1 g_9_25 (.ZN (n_9_25), .A (n_10_24), .B (n_8_27), .C1 (n_7_26), .C2 (n_12_22) );
AOI211_X1 g_11_24 (.ZN (n_11_24), .A (n_8_23), .B (n_6_26), .C1 (n_6_28), .C2 (n_10_23) );
AOI211_X1 g_10_22 (.ZN (n_10_22), .A (n_9_25), .B (n_8_25), .C1 (n_8_27), .C2 (n_8_24) );
AOI211_X1 g_12_21 (.ZN (n_12_21), .A (n_11_24), .B (n_10_24), .C1 (n_6_26), .C2 (n_7_26) );
AOI211_X1 g_14_20 (.ZN (n_14_20), .A (n_10_22), .B (n_8_23), .C1 (n_8_25), .C2 (n_6_28) );
AOI211_X1 g_16_19 (.ZN (n_16_19), .A (n_12_21), .B (n_9_25), .C1 (n_10_24), .C2 (n_8_27) );
AOI211_X1 g_18_18 (.ZN (n_18_18), .A (n_14_20), .B (n_11_24), .C1 (n_8_23), .C2 (n_6_26) );
AOI211_X1 g_20_19 (.ZN (n_20_19), .A (n_16_19), .B (n_10_22), .C1 (n_9_25), .C2 (n_8_25) );
AOI211_X1 g_18_20 (.ZN (n_18_20), .A (n_18_18), .B (n_12_21), .C1 (n_11_24), .C2 (n_10_24) );
AOI211_X1 g_16_21 (.ZN (n_16_21), .A (n_20_19), .B (n_14_20), .C1 (n_10_22), .C2 (n_8_23) );
AOI211_X1 g_14_22 (.ZN (n_14_22), .A (n_18_20), .B (n_16_19), .C1 (n_12_21), .C2 (n_9_25) );
AOI211_X1 g_12_23 (.ZN (n_12_23), .A (n_16_21), .B (n_18_18), .C1 (n_14_20), .C2 (n_11_24) );
AOI211_X1 g_11_25 (.ZN (n_11_25), .A (n_14_22), .B (n_20_19), .C1 (n_16_19), .C2 (n_10_22) );
AOI211_X1 g_9_24 (.ZN (n_9_24), .A (n_12_23), .B (n_18_20), .C1 (n_18_18), .C2 (n_12_21) );
AOI211_X1 g_11_23 (.ZN (n_11_23), .A (n_11_25), .B (n_16_21), .C1 (n_20_19), .C2 (n_14_20) );
AOI211_X1 g_13_22 (.ZN (n_13_22), .A (n_9_24), .B (n_14_22), .C1 (n_18_20), .C2 (n_16_19) );
AOI211_X1 g_15_21 (.ZN (n_15_21), .A (n_11_23), .B (n_12_23), .C1 (n_16_21), .C2 (n_18_18) );
AOI211_X1 g_17_20 (.ZN (n_17_20), .A (n_13_22), .B (n_11_25), .C1 (n_14_22), .C2 (n_20_19) );
AOI211_X1 g_19_19 (.ZN (n_19_19), .A (n_15_21), .B (n_9_24), .C1 (n_12_23), .C2 (n_18_20) );
AOI211_X1 g_21_18 (.ZN (n_21_18), .A (n_17_20), .B (n_11_23), .C1 (n_11_25), .C2 (n_16_21) );
AOI211_X1 g_23_17 (.ZN (n_23_17), .A (n_19_19), .B (n_13_22), .C1 (n_9_24), .C2 (n_14_22) );
AOI211_X1 g_25_16 (.ZN (n_25_16), .A (n_21_18), .B (n_15_21), .C1 (n_11_23), .C2 (n_12_23) );
AOI211_X1 g_27_15 (.ZN (n_27_15), .A (n_23_17), .B (n_17_20), .C1 (n_13_22), .C2 (n_11_25) );
AOI211_X1 g_29_14 (.ZN (n_29_14), .A (n_25_16), .B (n_19_19), .C1 (n_15_21), .C2 (n_9_24) );
AOI211_X1 g_31_13 (.ZN (n_31_13), .A (n_27_15), .B (n_21_18), .C1 (n_17_20), .C2 (n_11_23) );
AOI211_X1 g_33_12 (.ZN (n_33_12), .A (n_29_14), .B (n_23_17), .C1 (n_19_19), .C2 (n_13_22) );
AOI211_X1 g_35_11 (.ZN (n_35_11), .A (n_31_13), .B (n_25_16), .C1 (n_21_18), .C2 (n_15_21) );
AOI211_X1 g_37_10 (.ZN (n_37_10), .A (n_33_12), .B (n_27_15), .C1 (n_23_17), .C2 (n_17_20) );
AOI211_X1 g_39_9 (.ZN (n_39_9), .A (n_35_11), .B (n_29_14), .C1 (n_25_16), .C2 (n_19_19) );
AOI211_X1 g_41_8 (.ZN (n_41_8), .A (n_37_10), .B (n_31_13), .C1 (n_27_15), .C2 (n_21_18) );
AOI211_X1 g_43_7 (.ZN (n_43_7), .A (n_39_9), .B (n_33_12), .C1 (n_29_14), .C2 (n_23_17) );
AOI211_X1 g_45_6 (.ZN (n_45_6), .A (n_41_8), .B (n_35_11), .C1 (n_31_13), .C2 (n_25_16) );
AOI211_X1 g_47_5 (.ZN (n_47_5), .A (n_43_7), .B (n_37_10), .C1 (n_33_12), .C2 (n_27_15) );
AOI211_X1 g_49_4 (.ZN (n_49_4), .A (n_45_6), .B (n_39_9), .C1 (n_35_11), .C2 (n_29_14) );
AOI211_X1 g_51_3 (.ZN (n_51_3), .A (n_47_5), .B (n_41_8), .C1 (n_37_10), .C2 (n_31_13) );
AOI211_X1 g_50_5 (.ZN (n_50_5), .A (n_49_4), .B (n_43_7), .C1 (n_39_9), .C2 (n_33_12) );
AOI211_X1 g_48_6 (.ZN (n_48_6), .A (n_51_3), .B (n_45_6), .C1 (n_41_8), .C2 (n_35_11) );
AOI211_X1 g_46_7 (.ZN (n_46_7), .A (n_50_5), .B (n_47_5), .C1 (n_43_7), .C2 (n_37_10) );
AOI211_X1 g_44_8 (.ZN (n_44_8), .A (n_48_6), .B (n_49_4), .C1 (n_45_6), .C2 (n_39_9) );
AOI211_X1 g_42_9 (.ZN (n_42_9), .A (n_46_7), .B (n_51_3), .C1 (n_47_5), .C2 (n_41_8) );
AOI211_X1 g_40_10 (.ZN (n_40_10), .A (n_44_8), .B (n_50_5), .C1 (n_49_4), .C2 (n_43_7) );
AOI211_X1 g_38_11 (.ZN (n_38_11), .A (n_42_9), .B (n_48_6), .C1 (n_51_3), .C2 (n_45_6) );
AOI211_X1 g_36_12 (.ZN (n_36_12), .A (n_40_10), .B (n_46_7), .C1 (n_50_5), .C2 (n_47_5) );
AOI211_X1 g_34_13 (.ZN (n_34_13), .A (n_38_11), .B (n_44_8), .C1 (n_48_6), .C2 (n_49_4) );
AOI211_X1 g_32_14 (.ZN (n_32_14), .A (n_36_12), .B (n_42_9), .C1 (n_46_7), .C2 (n_51_3) );
AOI211_X1 g_30_15 (.ZN (n_30_15), .A (n_34_13), .B (n_40_10), .C1 (n_44_8), .C2 (n_50_5) );
AOI211_X1 g_28_16 (.ZN (n_28_16), .A (n_32_14), .B (n_38_11), .C1 (n_42_9), .C2 (n_48_6) );
AOI211_X1 g_26_17 (.ZN (n_26_17), .A (n_30_15), .B (n_36_12), .C1 (n_40_10), .C2 (n_46_7) );
AOI211_X1 g_24_18 (.ZN (n_24_18), .A (n_28_16), .B (n_34_13), .C1 (n_38_11), .C2 (n_44_8) );
AOI211_X1 g_22_19 (.ZN (n_22_19), .A (n_26_17), .B (n_32_14), .C1 (n_36_12), .C2 (n_42_9) );
AOI211_X1 g_20_20 (.ZN (n_20_20), .A (n_24_18), .B (n_30_15), .C1 (n_34_13), .C2 (n_40_10) );
AOI211_X1 g_18_21 (.ZN (n_18_21), .A (n_22_19), .B (n_28_16), .C1 (n_32_14), .C2 (n_38_11) );
AOI211_X1 g_16_22 (.ZN (n_16_22), .A (n_20_20), .B (n_26_17), .C1 (n_30_15), .C2 (n_36_12) );
AOI211_X1 g_14_23 (.ZN (n_14_23), .A (n_18_21), .B (n_24_18), .C1 (n_28_16), .C2 (n_34_13) );
AOI211_X1 g_12_24 (.ZN (n_12_24), .A (n_16_22), .B (n_22_19), .C1 (n_26_17), .C2 (n_32_14) );
AOI211_X1 g_10_25 (.ZN (n_10_25), .A (n_14_23), .B (n_20_20), .C1 (n_24_18), .C2 (n_30_15) );
AOI211_X1 g_8_26 (.ZN (n_8_26), .A (n_12_24), .B (n_18_21), .C1 (n_22_19), .C2 (n_28_16) );
AOI211_X1 g_6_27 (.ZN (n_6_27), .A (n_10_25), .B (n_16_22), .C1 (n_20_20), .C2 (n_26_17) );
AOI211_X1 g_5_29 (.ZN (n_5_29), .A (n_8_26), .B (n_14_23), .C1 (n_18_21), .C2 (n_24_18) );
AOI211_X1 g_7_28 (.ZN (n_7_28), .A (n_6_27), .B (n_12_24), .C1 (n_16_22), .C2 (n_22_19) );
AOI211_X1 g_9_27 (.ZN (n_9_27), .A (n_5_29), .B (n_10_25), .C1 (n_14_23), .C2 (n_20_20) );
AOI211_X1 g_11_26 (.ZN (n_11_26), .A (n_7_28), .B (n_8_26), .C1 (n_12_24), .C2 (n_18_21) );
AOI211_X1 g_13_25 (.ZN (n_13_25), .A (n_9_27), .B (n_6_27), .C1 (n_10_25), .C2 (n_16_22) );
AOI211_X1 g_15_24 (.ZN (n_15_24), .A (n_11_26), .B (n_5_29), .C1 (n_8_26), .C2 (n_14_23) );
AOI211_X1 g_13_23 (.ZN (n_13_23), .A (n_13_25), .B (n_7_28), .C1 (n_6_27), .C2 (n_12_24) );
AOI211_X1 g_15_22 (.ZN (n_15_22), .A (n_15_24), .B (n_9_27), .C1 (n_5_29), .C2 (n_10_25) );
AOI211_X1 g_17_21 (.ZN (n_17_21), .A (n_13_23), .B (n_11_26), .C1 (n_7_28), .C2 (n_8_26) );
AOI211_X1 g_19_20 (.ZN (n_19_20), .A (n_15_22), .B (n_13_25), .C1 (n_9_27), .C2 (n_6_27) );
AOI211_X1 g_21_19 (.ZN (n_21_19), .A (n_17_21), .B (n_15_24), .C1 (n_11_26), .C2 (n_5_29) );
AOI211_X1 g_20_21 (.ZN (n_20_21), .A (n_19_20), .B (n_13_23), .C1 (n_13_25), .C2 (n_7_28) );
AOI211_X1 g_22_20 (.ZN (n_22_20), .A (n_21_19), .B (n_15_22), .C1 (n_15_24), .C2 (n_9_27) );
AOI211_X1 g_24_19 (.ZN (n_24_19), .A (n_20_21), .B (n_17_21), .C1 (n_13_23), .C2 (n_11_26) );
AOI211_X1 g_26_18 (.ZN (n_26_18), .A (n_22_20), .B (n_19_20), .C1 (n_15_22), .C2 (n_13_25) );
AOI211_X1 g_24_17 (.ZN (n_24_17), .A (n_24_19), .B (n_21_19), .C1 (n_17_21), .C2 (n_15_24) );
AOI211_X1 g_26_16 (.ZN (n_26_16), .A (n_26_18), .B (n_20_21), .C1 (n_19_20), .C2 (n_13_23) );
AOI211_X1 g_28_15 (.ZN (n_28_15), .A (n_24_17), .B (n_22_20), .C1 (n_21_19), .C2 (n_15_22) );
AOI211_X1 g_30_14 (.ZN (n_30_14), .A (n_26_16), .B (n_24_19), .C1 (n_20_21), .C2 (n_17_21) );
AOI211_X1 g_32_13 (.ZN (n_32_13), .A (n_28_15), .B (n_26_18), .C1 (n_22_20), .C2 (n_19_20) );
AOI211_X1 g_34_12 (.ZN (n_34_12), .A (n_30_14), .B (n_24_17), .C1 (n_24_19), .C2 (n_21_19) );
AOI211_X1 g_36_11 (.ZN (n_36_11), .A (n_32_13), .B (n_26_16), .C1 (n_26_18), .C2 (n_20_21) );
AOI211_X1 g_38_10 (.ZN (n_38_10), .A (n_34_12), .B (n_28_15), .C1 (n_24_17), .C2 (n_22_20) );
AOI211_X1 g_40_9 (.ZN (n_40_9), .A (n_36_11), .B (n_30_14), .C1 (n_26_16), .C2 (n_24_19) );
AOI211_X1 g_42_8 (.ZN (n_42_8), .A (n_38_10), .B (n_32_13), .C1 (n_28_15), .C2 (n_26_18) );
AOI211_X1 g_44_7 (.ZN (n_44_7), .A (n_40_9), .B (n_34_12), .C1 (n_30_14), .C2 (n_24_17) );
AOI211_X1 g_46_6 (.ZN (n_46_6), .A (n_42_8), .B (n_36_11), .C1 (n_32_13), .C2 (n_26_16) );
AOI211_X1 g_48_5 (.ZN (n_48_5), .A (n_44_7), .B (n_38_10), .C1 (n_34_12), .C2 (n_28_15) );
AOI211_X1 g_50_4 (.ZN (n_50_4), .A (n_46_6), .B (n_40_9), .C1 (n_36_11), .C2 (n_30_14) );
AOI211_X1 g_51_6 (.ZN (n_51_6), .A (n_48_5), .B (n_42_8), .C1 (n_38_10), .C2 (n_32_13) );
AOI211_X1 g_49_7 (.ZN (n_49_7), .A (n_50_4), .B (n_44_7), .C1 (n_40_9), .C2 (n_34_12) );
AOI211_X1 g_47_8 (.ZN (n_47_8), .A (n_51_6), .B (n_46_6), .C1 (n_42_8), .C2 (n_36_11) );
AOI211_X1 g_45_9 (.ZN (n_45_9), .A (n_49_7), .B (n_48_5), .C1 (n_44_7), .C2 (n_38_10) );
AOI211_X1 g_43_10 (.ZN (n_43_10), .A (n_47_8), .B (n_50_4), .C1 (n_46_6), .C2 (n_40_9) );
AOI211_X1 g_41_11 (.ZN (n_41_11), .A (n_45_9), .B (n_51_6), .C1 (n_48_5), .C2 (n_42_8) );
AOI211_X1 g_39_12 (.ZN (n_39_12), .A (n_43_10), .B (n_49_7), .C1 (n_50_4), .C2 (n_44_7) );
AOI211_X1 g_37_13 (.ZN (n_37_13), .A (n_41_11), .B (n_47_8), .C1 (n_51_6), .C2 (n_46_6) );
AOI211_X1 g_35_14 (.ZN (n_35_14), .A (n_39_12), .B (n_45_9), .C1 (n_49_7), .C2 (n_48_5) );
AOI211_X1 g_33_15 (.ZN (n_33_15), .A (n_37_13), .B (n_43_10), .C1 (n_47_8), .C2 (n_50_4) );
AOI211_X1 g_31_16 (.ZN (n_31_16), .A (n_35_14), .B (n_41_11), .C1 (n_45_9), .C2 (n_51_6) );
AOI211_X1 g_29_17 (.ZN (n_29_17), .A (n_33_15), .B (n_39_12), .C1 (n_43_10), .C2 (n_49_7) );
AOI211_X1 g_27_18 (.ZN (n_27_18), .A (n_31_16), .B (n_37_13), .C1 (n_41_11), .C2 (n_47_8) );
AOI211_X1 g_25_19 (.ZN (n_25_19), .A (n_29_17), .B (n_35_14), .C1 (n_39_12), .C2 (n_45_9) );
AOI211_X1 g_23_20 (.ZN (n_23_20), .A (n_27_18), .B (n_33_15), .C1 (n_37_13), .C2 (n_43_10) );
AOI211_X1 g_21_21 (.ZN (n_21_21), .A (n_25_19), .B (n_31_16), .C1 (n_35_14), .C2 (n_41_11) );
AOI211_X1 g_19_22 (.ZN (n_19_22), .A (n_23_20), .B (n_29_17), .C1 (n_33_15), .C2 (n_39_12) );
AOI211_X1 g_17_23 (.ZN (n_17_23), .A (n_21_21), .B (n_27_18), .C1 (n_31_16), .C2 (n_37_13) );
AOI211_X1 g_16_25 (.ZN (n_16_25), .A (n_19_22), .B (n_25_19), .C1 (n_29_17), .C2 (n_35_14) );
AOI211_X1 g_15_23 (.ZN (n_15_23), .A (n_17_23), .B (n_23_20), .C1 (n_27_18), .C2 (n_33_15) );
AOI211_X1 g_13_24 (.ZN (n_13_24), .A (n_16_25), .B (n_21_21), .C1 (n_25_19), .C2 (n_31_16) );
AOI211_X1 g_12_26 (.ZN (n_12_26), .A (n_15_23), .B (n_19_22), .C1 (n_23_20), .C2 (n_29_17) );
AOI211_X1 g_14_25 (.ZN (n_14_25), .A (n_13_24), .B (n_17_23), .C1 (n_21_21), .C2 (n_27_18) );
AOI211_X1 g_16_24 (.ZN (n_16_24), .A (n_12_26), .B (n_16_25), .C1 (n_19_22), .C2 (n_25_19) );
AOI211_X1 g_17_22 (.ZN (n_17_22), .A (n_14_25), .B (n_15_23), .C1 (n_17_23), .C2 (n_23_20) );
AOI211_X1 g_19_21 (.ZN (n_19_21), .A (n_16_24), .B (n_13_24), .C1 (n_16_25), .C2 (n_21_21) );
AOI211_X1 g_21_20 (.ZN (n_21_20), .A (n_17_22), .B (n_12_26), .C1 (n_15_23), .C2 (n_19_22) );
AOI211_X1 g_23_19 (.ZN (n_23_19), .A (n_19_21), .B (n_14_25), .C1 (n_13_24), .C2 (n_17_23) );
AOI211_X1 g_25_18 (.ZN (n_25_18), .A (n_21_20), .B (n_16_24), .C1 (n_12_26), .C2 (n_16_25) );
AOI211_X1 g_27_17 (.ZN (n_27_17), .A (n_23_19), .B (n_17_22), .C1 (n_14_25), .C2 (n_15_23) );
AOI211_X1 g_29_16 (.ZN (n_29_16), .A (n_25_18), .B (n_19_21), .C1 (n_16_24), .C2 (n_13_24) );
AOI211_X1 g_31_15 (.ZN (n_31_15), .A (n_27_17), .B (n_21_20), .C1 (n_17_22), .C2 (n_12_26) );
AOI211_X1 g_33_14 (.ZN (n_33_14), .A (n_29_16), .B (n_23_19), .C1 (n_19_21), .C2 (n_14_25) );
AOI211_X1 g_35_13 (.ZN (n_35_13), .A (n_31_15), .B (n_25_18), .C1 (n_21_20), .C2 (n_16_24) );
AOI211_X1 g_37_12 (.ZN (n_37_12), .A (n_33_14), .B (n_27_17), .C1 (n_23_19), .C2 (n_17_22) );
AOI211_X1 g_39_11 (.ZN (n_39_11), .A (n_35_13), .B (n_29_16), .C1 (n_25_18), .C2 (n_19_21) );
AOI211_X1 g_41_10 (.ZN (n_41_10), .A (n_37_12), .B (n_31_15), .C1 (n_27_17), .C2 (n_21_20) );
AOI211_X1 g_43_9 (.ZN (n_43_9), .A (n_39_11), .B (n_33_14), .C1 (n_29_16), .C2 (n_23_19) );
AOI211_X1 g_45_8 (.ZN (n_45_8), .A (n_41_10), .B (n_35_13), .C1 (n_31_15), .C2 (n_25_18) );
AOI211_X1 g_47_7 (.ZN (n_47_7), .A (n_43_9), .B (n_37_12), .C1 (n_33_14), .C2 (n_27_17) );
AOI211_X1 g_49_6 (.ZN (n_49_6), .A (n_45_8), .B (n_39_11), .C1 (n_35_13), .C2 (n_29_16) );
AOI211_X1 g_51_5 (.ZN (n_51_5), .A (n_47_7), .B (n_41_10), .C1 (n_37_12), .C2 (n_31_15) );
AOI211_X1 g_53_4 (.ZN (n_53_4), .A (n_49_6), .B (n_43_9), .C1 (n_39_11), .C2 (n_33_14) );
AOI211_X1 g_52_6 (.ZN (n_52_6), .A (n_51_5), .B (n_45_8), .C1 (n_41_10), .C2 (n_35_13) );
AOI211_X1 g_50_7 (.ZN (n_50_7), .A (n_53_4), .B (n_47_7), .C1 (n_43_9), .C2 (n_37_12) );
AOI211_X1 g_48_8 (.ZN (n_48_8), .A (n_52_6), .B (n_49_6), .C1 (n_45_8), .C2 (n_39_11) );
AOI211_X1 g_46_9 (.ZN (n_46_9), .A (n_50_7), .B (n_51_5), .C1 (n_47_7), .C2 (n_41_10) );
AOI211_X1 g_44_10 (.ZN (n_44_10), .A (n_48_8), .B (n_53_4), .C1 (n_49_6), .C2 (n_43_9) );
AOI211_X1 g_42_11 (.ZN (n_42_11), .A (n_46_9), .B (n_52_6), .C1 (n_51_5), .C2 (n_45_8) );
AOI211_X1 g_40_12 (.ZN (n_40_12), .A (n_44_10), .B (n_50_7), .C1 (n_53_4), .C2 (n_47_7) );
AOI211_X1 g_38_13 (.ZN (n_38_13), .A (n_42_11), .B (n_48_8), .C1 (n_52_6), .C2 (n_49_6) );
AOI211_X1 g_36_14 (.ZN (n_36_14), .A (n_40_12), .B (n_46_9), .C1 (n_50_7), .C2 (n_51_5) );
AOI211_X1 g_34_15 (.ZN (n_34_15), .A (n_38_13), .B (n_44_10), .C1 (n_48_8), .C2 (n_53_4) );
AOI211_X1 g_32_16 (.ZN (n_32_16), .A (n_36_14), .B (n_42_11), .C1 (n_46_9), .C2 (n_52_6) );
AOI211_X1 g_30_17 (.ZN (n_30_17), .A (n_34_15), .B (n_40_12), .C1 (n_44_10), .C2 (n_50_7) );
AOI211_X1 g_28_18 (.ZN (n_28_18), .A (n_32_16), .B (n_38_13), .C1 (n_42_11), .C2 (n_48_8) );
AOI211_X1 g_26_19 (.ZN (n_26_19), .A (n_30_17), .B (n_36_14), .C1 (n_40_12), .C2 (n_46_9) );
AOI211_X1 g_24_20 (.ZN (n_24_20), .A (n_28_18), .B (n_34_15), .C1 (n_38_13), .C2 (n_44_10) );
AOI211_X1 g_22_21 (.ZN (n_22_21), .A (n_26_19), .B (n_32_16), .C1 (n_36_14), .C2 (n_42_11) );
AOI211_X1 g_20_22 (.ZN (n_20_22), .A (n_24_20), .B (n_30_17), .C1 (n_34_15), .C2 (n_40_12) );
AOI211_X1 g_18_23 (.ZN (n_18_23), .A (n_22_21), .B (n_28_18), .C1 (n_32_16), .C2 (n_38_13) );
AOI211_X1 g_17_25 (.ZN (n_17_25), .A (n_20_22), .B (n_26_19), .C1 (n_30_17), .C2 (n_36_14) );
AOI211_X1 g_16_23 (.ZN (n_16_23), .A (n_18_23), .B (n_24_20), .C1 (n_28_18), .C2 (n_34_15) );
AOI211_X1 g_18_22 (.ZN (n_18_22), .A (n_17_25), .B (n_22_21), .C1 (n_26_19), .C2 (n_32_16) );
AOI211_X1 g_19_24 (.ZN (n_19_24), .A (n_16_23), .B (n_20_22), .C1 (n_24_20), .C2 (n_30_17) );
AOI211_X1 g_21_23 (.ZN (n_21_23), .A (n_18_22), .B (n_18_23), .C1 (n_22_21), .C2 (n_28_18) );
AOI211_X1 g_23_22 (.ZN (n_23_22), .A (n_19_24), .B (n_17_25), .C1 (n_20_22), .C2 (n_26_19) );
AOI211_X1 g_25_21 (.ZN (n_25_21), .A (n_21_23), .B (n_16_23), .C1 (n_18_23), .C2 (n_24_20) );
AOI211_X1 g_27_20 (.ZN (n_27_20), .A (n_23_22), .B (n_18_22), .C1 (n_17_25), .C2 (n_22_21) );
AOI211_X1 g_29_19 (.ZN (n_29_19), .A (n_25_21), .B (n_19_24), .C1 (n_16_23), .C2 (n_20_22) );
AOI211_X1 g_28_17 (.ZN (n_28_17), .A (n_27_20), .B (n_21_23), .C1 (n_18_22), .C2 (n_18_23) );
AOI211_X1 g_30_16 (.ZN (n_30_16), .A (n_29_19), .B (n_23_22), .C1 (n_19_24), .C2 (n_17_25) );
AOI211_X1 g_32_15 (.ZN (n_32_15), .A (n_28_17), .B (n_25_21), .C1 (n_21_23), .C2 (n_16_23) );
AOI211_X1 g_34_14 (.ZN (n_34_14), .A (n_30_16), .B (n_27_20), .C1 (n_23_22), .C2 (n_18_22) );
AOI211_X1 g_36_13 (.ZN (n_36_13), .A (n_32_15), .B (n_29_19), .C1 (n_25_21), .C2 (n_19_24) );
AOI211_X1 g_38_12 (.ZN (n_38_12), .A (n_34_14), .B (n_28_17), .C1 (n_27_20), .C2 (n_21_23) );
AOI211_X1 g_40_11 (.ZN (n_40_11), .A (n_36_13), .B (n_30_16), .C1 (n_29_19), .C2 (n_23_22) );
AOI211_X1 g_42_10 (.ZN (n_42_10), .A (n_38_12), .B (n_32_15), .C1 (n_28_17), .C2 (n_25_21) );
AOI211_X1 g_44_9 (.ZN (n_44_9), .A (n_40_11), .B (n_34_14), .C1 (n_30_16), .C2 (n_27_20) );
AOI211_X1 g_46_8 (.ZN (n_46_8), .A (n_42_10), .B (n_36_13), .C1 (n_32_15), .C2 (n_29_19) );
AOI211_X1 g_48_7 (.ZN (n_48_7), .A (n_44_9), .B (n_38_12), .C1 (n_34_14), .C2 (n_28_17) );
AOI211_X1 g_50_6 (.ZN (n_50_6), .A (n_46_8), .B (n_40_11), .C1 (n_36_13), .C2 (n_30_16) );
AOI211_X1 g_52_5 (.ZN (n_52_5), .A (n_48_7), .B (n_42_10), .C1 (n_38_12), .C2 (n_32_15) );
AOI211_X1 g_53_7 (.ZN (n_53_7), .A (n_50_6), .B (n_44_9), .C1 (n_40_11), .C2 (n_34_14) );
AOI211_X1 g_51_8 (.ZN (n_51_8), .A (n_52_5), .B (n_46_8), .C1 (n_42_10), .C2 (n_36_13) );
AOI211_X1 g_49_9 (.ZN (n_49_9), .A (n_53_7), .B (n_48_7), .C1 (n_44_9), .C2 (n_38_12) );
AOI211_X1 g_47_10 (.ZN (n_47_10), .A (n_51_8), .B (n_50_6), .C1 (n_46_8), .C2 (n_40_11) );
AOI211_X1 g_45_11 (.ZN (n_45_11), .A (n_49_9), .B (n_52_5), .C1 (n_48_7), .C2 (n_42_10) );
AOI211_X1 g_43_12 (.ZN (n_43_12), .A (n_47_10), .B (n_53_7), .C1 (n_50_6), .C2 (n_44_9) );
AOI211_X1 g_41_13 (.ZN (n_41_13), .A (n_45_11), .B (n_51_8), .C1 (n_52_5), .C2 (n_46_8) );
AOI211_X1 g_39_14 (.ZN (n_39_14), .A (n_43_12), .B (n_49_9), .C1 (n_53_7), .C2 (n_48_7) );
AOI211_X1 g_37_15 (.ZN (n_37_15), .A (n_41_13), .B (n_47_10), .C1 (n_51_8), .C2 (n_50_6) );
AOI211_X1 g_35_16 (.ZN (n_35_16), .A (n_39_14), .B (n_45_11), .C1 (n_49_9), .C2 (n_52_5) );
AOI211_X1 g_33_17 (.ZN (n_33_17), .A (n_37_15), .B (n_43_12), .C1 (n_47_10), .C2 (n_53_7) );
AOI211_X1 g_31_18 (.ZN (n_31_18), .A (n_35_16), .B (n_41_13), .C1 (n_45_11), .C2 (n_51_8) );
AOI211_X1 g_30_20 (.ZN (n_30_20), .A (n_33_17), .B (n_39_14), .C1 (n_43_12), .C2 (n_49_9) );
AOI211_X1 g_29_18 (.ZN (n_29_18), .A (n_31_18), .B (n_37_15), .C1 (n_41_13), .C2 (n_47_10) );
AOI211_X1 g_31_17 (.ZN (n_31_17), .A (n_30_20), .B (n_35_16), .C1 (n_39_14), .C2 (n_45_11) );
AOI211_X1 g_33_16 (.ZN (n_33_16), .A (n_29_18), .B (n_33_17), .C1 (n_37_15), .C2 (n_43_12) );
AOI211_X1 g_35_15 (.ZN (n_35_15), .A (n_31_17), .B (n_31_18), .C1 (n_35_16), .C2 (n_41_13) );
AOI211_X1 g_37_14 (.ZN (n_37_14), .A (n_33_16), .B (n_30_20), .C1 (n_33_17), .C2 (n_39_14) );
AOI211_X1 g_39_13 (.ZN (n_39_13), .A (n_35_15), .B (n_29_18), .C1 (n_31_18), .C2 (n_37_15) );
AOI211_X1 g_41_12 (.ZN (n_41_12), .A (n_37_14), .B (n_31_17), .C1 (n_30_20), .C2 (n_35_16) );
AOI211_X1 g_43_11 (.ZN (n_43_11), .A (n_39_13), .B (n_33_16), .C1 (n_29_18), .C2 (n_33_17) );
AOI211_X1 g_45_10 (.ZN (n_45_10), .A (n_41_12), .B (n_35_15), .C1 (n_31_17), .C2 (n_31_18) );
AOI211_X1 g_47_9 (.ZN (n_47_9), .A (n_43_11), .B (n_37_14), .C1 (n_33_16), .C2 (n_30_20) );
AOI211_X1 g_49_8 (.ZN (n_49_8), .A (n_45_10), .B (n_39_13), .C1 (n_35_15), .C2 (n_29_18) );
AOI211_X1 g_51_7 (.ZN (n_51_7), .A (n_47_9), .B (n_41_12), .C1 (n_37_14), .C2 (n_31_17) );
AOI211_X1 g_53_6 (.ZN (n_53_6), .A (n_49_8), .B (n_43_11), .C1 (n_39_13), .C2 (n_33_16) );
AOI211_X1 g_55_5 (.ZN (n_55_5), .A (n_51_7), .B (n_45_10), .C1 (n_41_12), .C2 (n_35_15) );
AOI211_X1 g_54_7 (.ZN (n_54_7), .A (n_53_6), .B (n_47_9), .C1 (n_43_11), .C2 (n_37_14) );
AOI211_X1 g_52_8 (.ZN (n_52_8), .A (n_55_5), .B (n_49_8), .C1 (n_45_10), .C2 (n_39_13) );
AOI211_X1 g_50_9 (.ZN (n_50_9), .A (n_54_7), .B (n_51_7), .C1 (n_47_9), .C2 (n_41_12) );
AOI211_X1 g_48_10 (.ZN (n_48_10), .A (n_52_8), .B (n_53_6), .C1 (n_49_8), .C2 (n_43_11) );
AOI211_X1 g_46_11 (.ZN (n_46_11), .A (n_50_9), .B (n_55_5), .C1 (n_51_7), .C2 (n_45_10) );
AOI211_X1 g_44_12 (.ZN (n_44_12), .A (n_48_10), .B (n_54_7), .C1 (n_53_6), .C2 (n_47_9) );
AOI211_X1 g_42_13 (.ZN (n_42_13), .A (n_46_11), .B (n_52_8), .C1 (n_55_5), .C2 (n_49_8) );
AOI211_X1 g_40_14 (.ZN (n_40_14), .A (n_44_12), .B (n_50_9), .C1 (n_54_7), .C2 (n_51_7) );
AOI211_X1 g_38_15 (.ZN (n_38_15), .A (n_42_13), .B (n_48_10), .C1 (n_52_8), .C2 (n_53_6) );
AOI211_X1 g_36_16 (.ZN (n_36_16), .A (n_40_14), .B (n_46_11), .C1 (n_50_9), .C2 (n_55_5) );
AOI211_X1 g_34_17 (.ZN (n_34_17), .A (n_38_15), .B (n_44_12), .C1 (n_48_10), .C2 (n_54_7) );
AOI211_X1 g_32_18 (.ZN (n_32_18), .A (n_36_16), .B (n_42_13), .C1 (n_46_11), .C2 (n_52_8) );
AOI211_X1 g_30_19 (.ZN (n_30_19), .A (n_34_17), .B (n_40_14), .C1 (n_44_12), .C2 (n_50_9) );
AOI211_X1 g_28_20 (.ZN (n_28_20), .A (n_32_18), .B (n_38_15), .C1 (n_42_13), .C2 (n_48_10) );
AOI211_X1 g_26_21 (.ZN (n_26_21), .A (n_30_19), .B (n_36_16), .C1 (n_40_14), .C2 (n_46_11) );
AOI211_X1 g_27_19 (.ZN (n_27_19), .A (n_28_20), .B (n_34_17), .C1 (n_38_15), .C2 (n_44_12) );
AOI211_X1 g_25_20 (.ZN (n_25_20), .A (n_26_21), .B (n_32_18), .C1 (n_36_16), .C2 (n_42_13) );
AOI211_X1 g_23_21 (.ZN (n_23_21), .A (n_27_19), .B (n_30_19), .C1 (n_34_17), .C2 (n_40_14) );
AOI211_X1 g_21_22 (.ZN (n_21_22), .A (n_25_20), .B (n_28_20), .C1 (n_32_18), .C2 (n_38_15) );
AOI211_X1 g_19_23 (.ZN (n_19_23), .A (n_23_21), .B (n_26_21), .C1 (n_30_19), .C2 (n_36_16) );
AOI211_X1 g_17_24 (.ZN (n_17_24), .A (n_21_22), .B (n_27_19), .C1 (n_28_20), .C2 (n_34_17) );
AOI211_X1 g_15_25 (.ZN (n_15_25), .A (n_19_23), .B (n_25_20), .C1 (n_26_21), .C2 (n_32_18) );
AOI211_X1 g_13_26 (.ZN (n_13_26), .A (n_17_24), .B (n_23_21), .C1 (n_27_19), .C2 (n_30_19) );
AOI211_X1 g_14_24 (.ZN (n_14_24), .A (n_15_25), .B (n_21_22), .C1 (n_25_20), .C2 (n_28_20) );
AOI211_X1 g_12_25 (.ZN (n_12_25), .A (n_13_26), .B (n_19_23), .C1 (n_23_21), .C2 (n_26_21) );
AOI211_X1 g_10_26 (.ZN (n_10_26), .A (n_14_24), .B (n_17_24), .C1 (n_21_22), .C2 (n_27_19) );
AOI211_X1 g_11_28 (.ZN (n_11_28), .A (n_12_25), .B (n_15_25), .C1 (n_19_23), .C2 (n_25_20) );
AOI211_X1 g_13_27 (.ZN (n_13_27), .A (n_10_26), .B (n_13_26), .C1 (n_17_24), .C2 (n_23_21) );
AOI211_X1 g_15_26 (.ZN (n_15_26), .A (n_11_28), .B (n_14_24), .C1 (n_15_25), .C2 (n_21_22) );
AOI211_X1 g_14_28 (.ZN (n_14_28), .A (n_13_27), .B (n_12_25), .C1 (n_13_26), .C2 (n_19_23) );
AOI211_X1 g_12_27 (.ZN (n_12_27), .A (n_15_26), .B (n_10_26), .C1 (n_14_24), .C2 (n_17_24) );
AOI211_X1 g_14_26 (.ZN (n_14_26), .A (n_14_28), .B (n_11_28), .C1 (n_12_25), .C2 (n_15_25) );
AOI211_X1 g_16_27 (.ZN (n_16_27), .A (n_12_27), .B (n_13_27), .C1 (n_10_26), .C2 (n_13_26) );
AOI211_X1 g_18_26 (.ZN (n_18_26), .A (n_14_26), .B (n_15_26), .C1 (n_11_28), .C2 (n_14_24) );
AOI211_X1 g_20_25 (.ZN (n_20_25), .A (n_16_27), .B (n_14_28), .C1 (n_13_27), .C2 (n_12_25) );
AOI211_X1 g_18_24 (.ZN (n_18_24), .A (n_18_26), .B (n_12_27), .C1 (n_15_26), .C2 (n_10_26) );
AOI211_X1 g_20_23 (.ZN (n_20_23), .A (n_20_25), .B (n_14_26), .C1 (n_14_28), .C2 (n_11_28) );
AOI211_X1 g_22_22 (.ZN (n_22_22), .A (n_18_24), .B (n_16_27), .C1 (n_12_27), .C2 (n_13_27) );
AOI211_X1 g_24_21 (.ZN (n_24_21), .A (n_20_23), .B (n_18_26), .C1 (n_14_26), .C2 (n_15_26) );
AOI211_X1 g_26_20 (.ZN (n_26_20), .A (n_22_22), .B (n_20_25), .C1 (n_16_27), .C2 (n_14_28) );
AOI211_X1 g_28_19 (.ZN (n_28_19), .A (n_24_21), .B (n_18_24), .C1 (n_18_26), .C2 (n_12_27) );
AOI211_X1 g_30_18 (.ZN (n_30_18), .A (n_26_20), .B (n_20_23), .C1 (n_20_25), .C2 (n_14_26) );
AOI211_X1 g_32_17 (.ZN (n_32_17), .A (n_28_19), .B (n_22_22), .C1 (n_18_24), .C2 (n_16_27) );
AOI211_X1 g_34_16 (.ZN (n_34_16), .A (n_30_18), .B (n_24_21), .C1 (n_20_23), .C2 (n_18_26) );
AOI211_X1 g_36_15 (.ZN (n_36_15), .A (n_32_17), .B (n_26_20), .C1 (n_22_22), .C2 (n_20_25) );
AOI211_X1 g_38_14 (.ZN (n_38_14), .A (n_34_16), .B (n_28_19), .C1 (n_24_21), .C2 (n_18_24) );
AOI211_X1 g_40_13 (.ZN (n_40_13), .A (n_36_15), .B (n_30_18), .C1 (n_26_20), .C2 (n_20_23) );
AOI211_X1 g_42_12 (.ZN (n_42_12), .A (n_38_14), .B (n_32_17), .C1 (n_28_19), .C2 (n_22_22) );
AOI211_X1 g_44_11 (.ZN (n_44_11), .A (n_40_13), .B (n_34_16), .C1 (n_30_18), .C2 (n_24_21) );
AOI211_X1 g_46_10 (.ZN (n_46_10), .A (n_42_12), .B (n_36_15), .C1 (n_32_17), .C2 (n_26_20) );
AOI211_X1 g_48_9 (.ZN (n_48_9), .A (n_44_11), .B (n_38_14), .C1 (n_34_16), .C2 (n_28_19) );
AOI211_X1 g_50_8 (.ZN (n_50_8), .A (n_46_10), .B (n_40_13), .C1 (n_36_15), .C2 (n_30_18) );
AOI211_X1 g_52_7 (.ZN (n_52_7), .A (n_48_9), .B (n_42_12), .C1 (n_38_14), .C2 (n_32_17) );
AOI211_X1 g_54_6 (.ZN (n_54_6), .A (n_50_8), .B (n_44_11), .C1 (n_40_13), .C2 (n_34_16) );
AOI211_X1 g_56_7 (.ZN (n_56_7), .A (n_52_7), .B (n_46_10), .C1 (n_42_12), .C2 (n_36_15) );
AOI211_X1 g_54_8 (.ZN (n_54_8), .A (n_54_6), .B (n_48_9), .C1 (n_44_11), .C2 (n_38_14) );
AOI211_X1 g_52_9 (.ZN (n_52_9), .A (n_56_7), .B (n_50_8), .C1 (n_46_10), .C2 (n_40_13) );
AOI211_X1 g_50_10 (.ZN (n_50_10), .A (n_54_8), .B (n_52_7), .C1 (n_48_9), .C2 (n_42_12) );
AOI211_X1 g_48_11 (.ZN (n_48_11), .A (n_52_9), .B (n_54_6), .C1 (n_50_8), .C2 (n_44_11) );
AOI211_X1 g_46_12 (.ZN (n_46_12), .A (n_50_10), .B (n_56_7), .C1 (n_52_7), .C2 (n_46_10) );
AOI211_X1 g_44_13 (.ZN (n_44_13), .A (n_48_11), .B (n_54_8), .C1 (n_54_6), .C2 (n_48_9) );
AOI211_X1 g_42_14 (.ZN (n_42_14), .A (n_46_12), .B (n_52_9), .C1 (n_56_7), .C2 (n_50_8) );
AOI211_X1 g_40_15 (.ZN (n_40_15), .A (n_44_13), .B (n_50_10), .C1 (n_54_8), .C2 (n_52_7) );
AOI211_X1 g_38_16 (.ZN (n_38_16), .A (n_42_14), .B (n_48_11), .C1 (n_52_9), .C2 (n_54_6) );
AOI211_X1 g_36_17 (.ZN (n_36_17), .A (n_40_15), .B (n_46_12), .C1 (n_50_10), .C2 (n_56_7) );
AOI211_X1 g_34_18 (.ZN (n_34_18), .A (n_38_16), .B (n_44_13), .C1 (n_48_11), .C2 (n_54_8) );
AOI211_X1 g_32_19 (.ZN (n_32_19), .A (n_36_17), .B (n_42_14), .C1 (n_46_12), .C2 (n_52_9) );
AOI211_X1 g_31_21 (.ZN (n_31_21), .A (n_34_18), .B (n_40_15), .C1 (n_44_13), .C2 (n_50_10) );
AOI211_X1 g_29_20 (.ZN (n_29_20), .A (n_32_19), .B (n_38_16), .C1 (n_42_14), .C2 (n_48_11) );
AOI211_X1 g_31_19 (.ZN (n_31_19), .A (n_31_21), .B (n_36_17), .C1 (n_40_15), .C2 (n_46_12) );
AOI211_X1 g_33_18 (.ZN (n_33_18), .A (n_29_20), .B (n_34_18), .C1 (n_38_16), .C2 (n_44_13) );
AOI211_X1 g_35_17 (.ZN (n_35_17), .A (n_31_19), .B (n_32_19), .C1 (n_36_17), .C2 (n_42_14) );
AOI211_X1 g_37_16 (.ZN (n_37_16), .A (n_33_18), .B (n_31_21), .C1 (n_34_18), .C2 (n_40_15) );
AOI211_X1 g_39_15 (.ZN (n_39_15), .A (n_35_17), .B (n_29_20), .C1 (n_32_19), .C2 (n_38_16) );
AOI211_X1 g_41_14 (.ZN (n_41_14), .A (n_37_16), .B (n_31_19), .C1 (n_31_21), .C2 (n_36_17) );
AOI211_X1 g_43_13 (.ZN (n_43_13), .A (n_39_15), .B (n_33_18), .C1 (n_29_20), .C2 (n_34_18) );
AOI211_X1 g_45_12 (.ZN (n_45_12), .A (n_41_14), .B (n_35_17), .C1 (n_31_19), .C2 (n_32_19) );
AOI211_X1 g_47_11 (.ZN (n_47_11), .A (n_43_13), .B (n_37_16), .C1 (n_33_18), .C2 (n_31_21) );
AOI211_X1 g_49_10 (.ZN (n_49_10), .A (n_45_12), .B (n_39_15), .C1 (n_35_17), .C2 (n_29_20) );
AOI211_X1 g_51_9 (.ZN (n_51_9), .A (n_47_11), .B (n_41_14), .C1 (n_37_16), .C2 (n_31_19) );
AOI211_X1 g_53_8 (.ZN (n_53_8), .A (n_49_10), .B (n_43_13), .C1 (n_39_15), .C2 (n_33_18) );
AOI211_X1 g_55_7 (.ZN (n_55_7), .A (n_51_9), .B (n_45_12), .C1 (n_41_14), .C2 (n_35_17) );
AOI211_X1 g_57_6 (.ZN (n_57_6), .A (n_53_8), .B (n_47_11), .C1 (n_43_13), .C2 (n_37_16) );
AOI211_X1 g_58_8 (.ZN (n_58_8), .A (n_55_7), .B (n_49_10), .C1 (n_45_12), .C2 (n_39_15) );
AOI211_X1 g_56_9 (.ZN (n_56_9), .A (n_57_6), .B (n_51_9), .C1 (n_47_11), .C2 (n_41_14) );
AOI211_X1 g_54_10 (.ZN (n_54_10), .A (n_58_8), .B (n_53_8), .C1 (n_49_10), .C2 (n_43_13) );
AOI211_X1 g_52_11 (.ZN (n_52_11), .A (n_56_9), .B (n_55_7), .C1 (n_51_9), .C2 (n_45_12) );
AOI211_X1 g_53_9 (.ZN (n_53_9), .A (n_54_10), .B (n_57_6), .C1 (n_53_8), .C2 (n_47_11) );
AOI211_X1 g_51_10 (.ZN (n_51_10), .A (n_52_11), .B (n_58_8), .C1 (n_55_7), .C2 (n_49_10) );
AOI211_X1 g_49_11 (.ZN (n_49_11), .A (n_53_9), .B (n_56_9), .C1 (n_57_6), .C2 (n_51_9) );
AOI211_X1 g_47_12 (.ZN (n_47_12), .A (n_51_10), .B (n_54_10), .C1 (n_58_8), .C2 (n_53_8) );
AOI211_X1 g_45_13 (.ZN (n_45_13), .A (n_49_11), .B (n_52_11), .C1 (n_56_9), .C2 (n_55_7) );
AOI211_X1 g_43_14 (.ZN (n_43_14), .A (n_47_12), .B (n_53_9), .C1 (n_54_10), .C2 (n_57_6) );
AOI211_X1 g_41_15 (.ZN (n_41_15), .A (n_45_13), .B (n_51_10), .C1 (n_52_11), .C2 (n_58_8) );
AOI211_X1 g_39_16 (.ZN (n_39_16), .A (n_43_14), .B (n_49_11), .C1 (n_53_9), .C2 (n_56_9) );
AOI211_X1 g_37_17 (.ZN (n_37_17), .A (n_41_15), .B (n_47_12), .C1 (n_51_10), .C2 (n_54_10) );
AOI211_X1 g_35_18 (.ZN (n_35_18), .A (n_39_16), .B (n_45_13), .C1 (n_49_11), .C2 (n_52_11) );
AOI211_X1 g_33_19 (.ZN (n_33_19), .A (n_37_17), .B (n_43_14), .C1 (n_47_12), .C2 (n_53_9) );
AOI211_X1 g_31_20 (.ZN (n_31_20), .A (n_35_18), .B (n_41_15), .C1 (n_45_13), .C2 (n_51_10) );
AOI211_X1 g_29_21 (.ZN (n_29_21), .A (n_33_19), .B (n_39_16), .C1 (n_43_14), .C2 (n_49_11) );
AOI211_X1 g_27_22 (.ZN (n_27_22), .A (n_31_20), .B (n_37_17), .C1 (n_41_15), .C2 (n_47_12) );
AOI211_X1 g_25_23 (.ZN (n_25_23), .A (n_29_21), .B (n_35_18), .C1 (n_39_16), .C2 (n_45_13) );
AOI211_X1 g_23_24 (.ZN (n_23_24), .A (n_27_22), .B (n_33_19), .C1 (n_37_17), .C2 (n_43_14) );
AOI211_X1 g_24_22 (.ZN (n_24_22), .A (n_25_23), .B (n_31_20), .C1 (n_35_18), .C2 (n_41_15) );
AOI211_X1 g_22_23 (.ZN (n_22_23), .A (n_23_24), .B (n_29_21), .C1 (n_33_19), .C2 (n_39_16) );
AOI211_X1 g_20_24 (.ZN (n_20_24), .A (n_24_22), .B (n_27_22), .C1 (n_31_20), .C2 (n_37_17) );
AOI211_X1 g_18_25 (.ZN (n_18_25), .A (n_22_23), .B (n_25_23), .C1 (n_29_21), .C2 (n_35_18) );
AOI211_X1 g_16_26 (.ZN (n_16_26), .A (n_20_24), .B (n_23_24), .C1 (n_27_22), .C2 (n_33_19) );
AOI211_X1 g_14_27 (.ZN (n_14_27), .A (n_18_25), .B (n_24_22), .C1 (n_25_23), .C2 (n_31_20) );
AOI211_X1 g_12_28 (.ZN (n_12_28), .A (n_16_26), .B (n_22_23), .C1 (n_23_24), .C2 (n_29_21) );
AOI211_X1 g_10_27 (.ZN (n_10_27), .A (n_14_27), .B (n_20_24), .C1 (n_24_22), .C2 (n_27_22) );
AOI211_X1 g_9_29 (.ZN (n_9_29), .A (n_12_28), .B (n_18_25), .C1 (n_22_23), .C2 (n_25_23) );
AOI211_X1 g_7_30 (.ZN (n_7_30), .A (n_10_27), .B (n_16_26), .C1 (n_20_24), .C2 (n_23_24) );
AOI211_X1 g_8_28 (.ZN (n_8_28), .A (n_9_29), .B (n_14_27), .C1 (n_18_25), .C2 (n_24_22) );
AOI211_X1 g_9_26 (.ZN (n_9_26), .A (n_7_30), .B (n_12_28), .C1 (n_16_26), .C2 (n_22_23) );
AOI211_X1 g_7_27 (.ZN (n_7_27), .A (n_8_28), .B (n_10_27), .C1 (n_14_27), .C2 (n_20_24) );
AOI211_X1 g_5_28 (.ZN (n_5_28), .A (n_9_26), .B (n_9_29), .C1 (n_12_28), .C2 (n_18_25) );
AOI211_X1 g_4_30 (.ZN (n_4_30), .A (n_7_27), .B (n_7_30), .C1 (n_10_27), .C2 (n_16_26) );
AOI211_X1 g_6_29 (.ZN (n_6_29), .A (n_5_28), .B (n_8_28), .C1 (n_9_29), .C2 (n_14_27) );
AOI211_X1 g_5_31 (.ZN (n_5_31), .A (n_4_30), .B (n_9_26), .C1 (n_7_30), .C2 (n_12_28) );
AOI211_X1 g_3_32 (.ZN (n_3_32), .A (n_6_29), .B (n_7_27), .C1 (n_8_28), .C2 (n_10_27) );
AOI211_X1 g_2_34 (.ZN (n_2_34), .A (n_5_31), .B (n_5_28), .C1 (n_9_26), .C2 (n_9_29) );
AOI211_X1 g_1_36 (.ZN (n_1_36), .A (n_3_32), .B (n_4_30), .C1 (n_7_27), .C2 (n_7_30) );
AOI211_X1 g_3_35 (.ZN (n_3_35), .A (n_2_34), .B (n_6_29), .C1 (n_5_28), .C2 (n_8_28) );
AOI211_X1 g_4_33 (.ZN (n_4_33), .A (n_1_36), .B (n_5_31), .C1 (n_4_30), .C2 (n_9_26) );
AOI211_X1 g_6_32 (.ZN (n_6_32), .A (n_3_35), .B (n_3_32), .C1 (n_6_29), .C2 (n_7_27) );
AOI211_X1 g_4_31 (.ZN (n_4_31), .A (n_4_33), .B (n_2_34), .C1 (n_5_31), .C2 (n_5_28) );
AOI211_X1 g_3_33 (.ZN (n_3_33), .A (n_6_32), .B (n_1_36), .C1 (n_3_32), .C2 (n_4_30) );
AOI211_X1 g_5_34 (.ZN (n_5_34), .A (n_4_31), .B (n_3_35), .C1 (n_2_34), .C2 (n_6_29) );
AOI211_X1 g_7_33 (.ZN (n_7_33), .A (n_3_33), .B (n_4_33), .C1 (n_1_36), .C2 (n_5_31) );
AOI211_X1 g_6_31 (.ZN (n_6_31), .A (n_5_34), .B (n_6_32), .C1 (n_3_35), .C2 (n_3_32) );
AOI211_X1 g_7_29 (.ZN (n_7_29), .A (n_7_33), .B (n_4_31), .C1 (n_4_33), .C2 (n_2_34) );
AOI211_X1 g_9_28 (.ZN (n_9_28), .A (n_6_31), .B (n_3_33), .C1 (n_6_32), .C2 (n_1_36) );
AOI211_X1 g_11_27 (.ZN (n_11_27), .A (n_7_29), .B (n_5_34), .C1 (n_4_31), .C2 (n_3_35) );
AOI211_X1 g_10_29 (.ZN (n_10_29), .A (n_9_28), .B (n_7_33), .C1 (n_3_33), .C2 (n_4_33) );
AOI211_X1 g_8_30 (.ZN (n_8_30), .A (n_11_27), .B (n_6_31), .C1 (n_5_34), .C2 (n_6_32) );
AOI211_X1 g_7_32 (.ZN (n_7_32), .A (n_10_29), .B (n_7_29), .C1 (n_7_33), .C2 (n_4_31) );
AOI211_X1 g_6_30 (.ZN (n_6_30), .A (n_8_30), .B (n_9_28), .C1 (n_6_31), .C2 (n_3_33) );
AOI211_X1 g_5_32 (.ZN (n_5_32), .A (n_7_32), .B (n_11_27), .C1 (n_7_29), .C2 (n_5_34) );
AOI211_X1 g_4_34 (.ZN (n_4_34), .A (n_6_30), .B (n_10_29), .C1 (n_9_28), .C2 (n_7_33) );
AOI211_X1 g_3_36 (.ZN (n_3_36), .A (n_5_32), .B (n_8_30), .C1 (n_11_27), .C2 (n_6_31) );
AOI211_X1 g_2_38 (.ZN (n_2_38), .A (n_4_34), .B (n_7_32), .C1 (n_10_29), .C2 (n_7_29) );
AOI211_X1 g_1_40 (.ZN (n_1_40), .A (n_3_36), .B (n_6_30), .C1 (n_8_30), .C2 (n_9_28) );
AOI211_X1 g_3_39 (.ZN (n_3_39), .A (n_2_38), .B (n_5_32), .C1 (n_7_32), .C2 (n_11_27) );
AOI211_X1 g_4_37 (.ZN (n_4_37), .A (n_1_40), .B (n_4_34), .C1 (n_6_30), .C2 (n_10_29) );
AOI211_X1 g_5_35 (.ZN (n_5_35), .A (n_3_39), .B (n_3_36), .C1 (n_5_32), .C2 (n_8_30) );
AOI211_X1 g_6_33 (.ZN (n_6_33), .A (n_4_37), .B (n_2_38), .C1 (n_4_34), .C2 (n_7_32) );
AOI211_X1 g_7_31 (.ZN (n_7_31), .A (n_5_35), .B (n_1_40), .C1 (n_3_36), .C2 (n_6_30) );
AOI211_X1 g_8_29 (.ZN (n_8_29), .A (n_6_33), .B (n_3_39), .C1 (n_2_38), .C2 (n_5_32) );
AOI211_X1 g_10_28 (.ZN (n_10_28), .A (n_7_31), .B (n_4_37), .C1 (n_1_40), .C2 (n_4_34) );
AOI211_X1 g_9_30 (.ZN (n_9_30), .A (n_8_29), .B (n_5_35), .C1 (n_3_39), .C2 (n_3_36) );
AOI211_X1 g_11_29 (.ZN (n_11_29), .A (n_10_28), .B (n_6_33), .C1 (n_4_37), .C2 (n_2_38) );
AOI211_X1 g_13_28 (.ZN (n_13_28), .A (n_9_30), .B (n_7_31), .C1 (n_5_35), .C2 (n_1_40) );
AOI211_X1 g_15_27 (.ZN (n_15_27), .A (n_11_29), .B (n_8_29), .C1 (n_6_33), .C2 (n_3_39) );
AOI211_X1 g_17_26 (.ZN (n_17_26), .A (n_13_28), .B (n_10_28), .C1 (n_7_31), .C2 (n_4_37) );
AOI211_X1 g_19_25 (.ZN (n_19_25), .A (n_15_27), .B (n_9_30), .C1 (n_8_29), .C2 (n_5_35) );
AOI211_X1 g_21_24 (.ZN (n_21_24), .A (n_17_26), .B (n_11_29), .C1 (n_10_28), .C2 (n_6_33) );
AOI211_X1 g_23_23 (.ZN (n_23_23), .A (n_19_25), .B (n_13_28), .C1 (n_9_30), .C2 (n_7_31) );
AOI211_X1 g_25_22 (.ZN (n_25_22), .A (n_21_24), .B (n_15_27), .C1 (n_11_29), .C2 (n_8_29) );
AOI211_X1 g_27_21 (.ZN (n_27_21), .A (n_23_23), .B (n_17_26), .C1 (n_13_28), .C2 (n_10_28) );
AOI211_X1 g_29_22 (.ZN (n_29_22), .A (n_25_22), .B (n_19_25), .C1 (n_15_27), .C2 (n_9_30) );
AOI211_X1 g_27_23 (.ZN (n_27_23), .A (n_27_21), .B (n_21_24), .C1 (n_17_26), .C2 (n_11_29) );
AOI211_X1 g_28_21 (.ZN (n_28_21), .A (n_29_22), .B (n_23_23), .C1 (n_19_25), .C2 (n_13_28) );
AOI211_X1 g_26_22 (.ZN (n_26_22), .A (n_27_23), .B (n_25_22), .C1 (n_21_24), .C2 (n_15_27) );
AOI211_X1 g_24_23 (.ZN (n_24_23), .A (n_28_21), .B (n_27_21), .C1 (n_23_23), .C2 (n_17_26) );
AOI211_X1 g_22_24 (.ZN (n_22_24), .A (n_26_22), .B (n_29_22), .C1 (n_25_22), .C2 (n_19_25) );
AOI211_X1 g_21_26 (.ZN (n_21_26), .A (n_24_23), .B (n_27_23), .C1 (n_27_21), .C2 (n_21_24) );
AOI211_X1 g_23_25 (.ZN (n_23_25), .A (n_22_24), .B (n_28_21), .C1 (n_29_22), .C2 (n_23_23) );
AOI211_X1 g_25_24 (.ZN (n_25_24), .A (n_21_26), .B (n_26_22), .C1 (n_27_23), .C2 (n_25_22) );
AOI211_X1 g_24_26 (.ZN (n_24_26), .A (n_23_25), .B (n_24_23), .C1 (n_28_21), .C2 (n_27_21) );
AOI211_X1 g_22_25 (.ZN (n_22_25), .A (n_25_24), .B (n_22_24), .C1 (n_26_22), .C2 (n_29_22) );
AOI211_X1 g_24_24 (.ZN (n_24_24), .A (n_24_26), .B (n_21_26), .C1 (n_24_23), .C2 (n_27_23) );
AOI211_X1 g_26_23 (.ZN (n_26_23), .A (n_22_25), .B (n_23_25), .C1 (n_22_24), .C2 (n_28_21) );
AOI211_X1 g_28_22 (.ZN (n_28_22), .A (n_24_24), .B (n_25_24), .C1 (n_21_26), .C2 (n_26_22) );
AOI211_X1 g_30_21 (.ZN (n_30_21), .A (n_26_23), .B (n_24_26), .C1 (n_23_25), .C2 (n_24_23) );
AOI211_X1 g_32_20 (.ZN (n_32_20), .A (n_28_22), .B (n_22_25), .C1 (n_25_24), .C2 (n_22_24) );
AOI211_X1 g_34_19 (.ZN (n_34_19), .A (n_30_21), .B (n_24_24), .C1 (n_24_26), .C2 (n_21_26) );
AOI211_X1 g_36_18 (.ZN (n_36_18), .A (n_32_20), .B (n_26_23), .C1 (n_22_25), .C2 (n_23_25) );
AOI211_X1 g_38_17 (.ZN (n_38_17), .A (n_34_19), .B (n_28_22), .C1 (n_24_24), .C2 (n_25_24) );
AOI211_X1 g_40_16 (.ZN (n_40_16), .A (n_36_18), .B (n_30_21), .C1 (n_26_23), .C2 (n_24_26) );
AOI211_X1 g_42_15 (.ZN (n_42_15), .A (n_38_17), .B (n_32_20), .C1 (n_28_22), .C2 (n_22_25) );
AOI211_X1 g_44_14 (.ZN (n_44_14), .A (n_40_16), .B (n_34_19), .C1 (n_30_21), .C2 (n_24_24) );
AOI211_X1 g_46_13 (.ZN (n_46_13), .A (n_42_15), .B (n_36_18), .C1 (n_32_20), .C2 (n_26_23) );
AOI211_X1 g_48_12 (.ZN (n_48_12), .A (n_44_14), .B (n_38_17), .C1 (n_34_19), .C2 (n_28_22) );
AOI211_X1 g_50_11 (.ZN (n_50_11), .A (n_46_13), .B (n_40_16), .C1 (n_36_18), .C2 (n_30_21) );
AOI211_X1 g_52_10 (.ZN (n_52_10), .A (n_48_12), .B (n_42_15), .C1 (n_38_17), .C2 (n_32_20) );
AOI211_X1 g_54_9 (.ZN (n_54_9), .A (n_50_11), .B (n_44_14), .C1 (n_40_16), .C2 (n_34_19) );
AOI211_X1 g_56_8 (.ZN (n_56_8), .A (n_52_10), .B (n_46_13), .C1 (n_42_15), .C2 (n_36_18) );
AOI211_X1 g_58_7 (.ZN (n_58_7), .A (n_54_9), .B (n_48_12), .C1 (n_44_14), .C2 (n_38_17) );
AOI211_X1 g_57_9 (.ZN (n_57_9), .A (n_56_8), .B (n_50_11), .C1 (n_46_13), .C2 (n_40_16) );
AOI211_X1 g_55_10 (.ZN (n_55_10), .A (n_58_7), .B (n_52_10), .C1 (n_48_12), .C2 (n_42_15) );
AOI211_X1 g_53_11 (.ZN (n_53_11), .A (n_57_9), .B (n_54_9), .C1 (n_50_11), .C2 (n_44_14) );
AOI211_X1 g_51_12 (.ZN (n_51_12), .A (n_55_10), .B (n_56_8), .C1 (n_52_10), .C2 (n_46_13) );
AOI211_X1 g_49_13 (.ZN (n_49_13), .A (n_53_11), .B (n_58_7), .C1 (n_54_9), .C2 (n_48_12) );
AOI211_X1 g_47_14 (.ZN (n_47_14), .A (n_51_12), .B (n_57_9), .C1 (n_56_8), .C2 (n_50_11) );
AOI211_X1 g_45_15 (.ZN (n_45_15), .A (n_49_13), .B (n_55_10), .C1 (n_58_7), .C2 (n_52_10) );
AOI211_X1 g_43_16 (.ZN (n_43_16), .A (n_47_14), .B (n_53_11), .C1 (n_57_9), .C2 (n_54_9) );
AOI211_X1 g_41_17 (.ZN (n_41_17), .A (n_45_15), .B (n_51_12), .C1 (n_55_10), .C2 (n_56_8) );
AOI211_X1 g_39_18 (.ZN (n_39_18), .A (n_43_16), .B (n_49_13), .C1 (n_53_11), .C2 (n_58_7) );
AOI211_X1 g_37_19 (.ZN (n_37_19), .A (n_41_17), .B (n_47_14), .C1 (n_51_12), .C2 (n_57_9) );
AOI211_X1 g_35_20 (.ZN (n_35_20), .A (n_39_18), .B (n_45_15), .C1 (n_49_13), .C2 (n_55_10) );
AOI211_X1 g_33_21 (.ZN (n_33_21), .A (n_37_19), .B (n_43_16), .C1 (n_47_14), .C2 (n_53_11) );
AOI211_X1 g_31_22 (.ZN (n_31_22), .A (n_35_20), .B (n_41_17), .C1 (n_45_15), .C2 (n_51_12) );
AOI211_X1 g_29_23 (.ZN (n_29_23), .A (n_33_21), .B (n_39_18), .C1 (n_43_16), .C2 (n_49_13) );
AOI211_X1 g_27_24 (.ZN (n_27_24), .A (n_31_22), .B (n_37_19), .C1 (n_41_17), .C2 (n_47_14) );
AOI211_X1 g_25_25 (.ZN (n_25_25), .A (n_29_23), .B (n_35_20), .C1 (n_39_18), .C2 (n_45_15) );
AOI211_X1 g_23_26 (.ZN (n_23_26), .A (n_27_24), .B (n_33_21), .C1 (n_37_19), .C2 (n_43_16) );
AOI211_X1 g_21_25 (.ZN (n_21_25), .A (n_25_25), .B (n_31_22), .C1 (n_35_20), .C2 (n_41_17) );
AOI211_X1 g_19_26 (.ZN (n_19_26), .A (n_23_26), .B (n_29_23), .C1 (n_33_21), .C2 (n_39_18) );
AOI211_X1 g_17_27 (.ZN (n_17_27), .A (n_21_25), .B (n_27_24), .C1 (n_31_22), .C2 (n_37_19) );
AOI211_X1 g_15_28 (.ZN (n_15_28), .A (n_19_26), .B (n_25_25), .C1 (n_29_23), .C2 (n_35_20) );
AOI211_X1 g_13_29 (.ZN (n_13_29), .A (n_17_27), .B (n_23_26), .C1 (n_27_24), .C2 (n_33_21) );
AOI211_X1 g_11_30 (.ZN (n_11_30), .A (n_15_28), .B (n_21_25), .C1 (n_25_25), .C2 (n_31_22) );
AOI211_X1 g_9_31 (.ZN (n_9_31), .A (n_13_29), .B (n_19_26), .C1 (n_23_26), .C2 (n_29_23) );
AOI211_X1 g_8_33 (.ZN (n_8_33), .A (n_11_30), .B (n_17_27), .C1 (n_21_25), .C2 (n_27_24) );
AOI211_X1 g_6_34 (.ZN (n_6_34), .A (n_9_31), .B (n_15_28), .C1 (n_19_26), .C2 (n_25_25) );
AOI211_X1 g_4_35 (.ZN (n_4_35), .A (n_8_33), .B (n_13_29), .C1 (n_17_27), .C2 (n_23_26) );
AOI211_X1 g_5_33 (.ZN (n_5_33), .A (n_6_34), .B (n_11_30), .C1 (n_15_28), .C2 (n_21_25) );
AOI211_X1 g_6_35 (.ZN (n_6_35), .A (n_4_35), .B (n_9_31), .C1 (n_13_29), .C2 (n_19_26) );
AOI211_X1 g_5_37 (.ZN (n_5_37), .A (n_5_33), .B (n_8_33), .C1 (n_11_30), .C2 (n_17_27) );
AOI211_X1 g_7_36 (.ZN (n_7_36), .A (n_6_35), .B (n_6_34), .C1 (n_9_31), .C2 (n_15_28) );
AOI211_X1 g_8_34 (.ZN (n_8_34), .A (n_5_37), .B (n_4_35), .C1 (n_8_33), .C2 (n_13_29) );
AOI211_X1 g_9_32 (.ZN (n_9_32), .A (n_7_36), .B (n_5_33), .C1 (n_6_34), .C2 (n_11_30) );
AOI211_X1 g_10_30 (.ZN (n_10_30), .A (n_8_34), .B (n_6_35), .C1 (n_4_35), .C2 (n_9_31) );
AOI211_X1 g_8_31 (.ZN (n_8_31), .A (n_9_32), .B (n_5_37), .C1 (n_5_33), .C2 (n_8_33) );
AOI211_X1 g_10_32 (.ZN (n_10_32), .A (n_10_30), .B (n_7_36), .C1 (n_6_35), .C2 (n_6_34) );
AOI211_X1 g_12_31 (.ZN (n_12_31), .A (n_8_31), .B (n_8_34), .C1 (n_5_37), .C2 (n_4_35) );
AOI211_X1 g_14_30 (.ZN (n_14_30), .A (n_10_32), .B (n_9_32), .C1 (n_7_36), .C2 (n_5_33) );
AOI211_X1 g_12_29 (.ZN (n_12_29), .A (n_12_31), .B (n_10_30), .C1 (n_8_34), .C2 (n_6_35) );
AOI211_X1 g_11_31 (.ZN (n_11_31), .A (n_14_30), .B (n_8_31), .C1 (n_9_32), .C2 (n_5_37) );
AOI211_X1 g_13_30 (.ZN (n_13_30), .A (n_12_29), .B (n_10_32), .C1 (n_10_30), .C2 (n_7_36) );
AOI211_X1 g_15_29 (.ZN (n_15_29), .A (n_11_31), .B (n_12_31), .C1 (n_8_31), .C2 (n_8_34) );
AOI211_X1 g_17_28 (.ZN (n_17_28), .A (n_13_30), .B (n_14_30), .C1 (n_10_32), .C2 (n_9_32) );
AOI211_X1 g_19_27 (.ZN (n_19_27), .A (n_15_29), .B (n_12_29), .C1 (n_12_31), .C2 (n_10_30) );
AOI211_X1 g_18_29 (.ZN (n_18_29), .A (n_17_28), .B (n_11_31), .C1 (n_14_30), .C2 (n_8_31) );
AOI211_X1 g_16_28 (.ZN (n_16_28), .A (n_19_27), .B (n_13_30), .C1 (n_12_29), .C2 (n_10_32) );
AOI211_X1 g_18_27 (.ZN (n_18_27), .A (n_18_29), .B (n_15_29), .C1 (n_11_31), .C2 (n_12_31) );
AOI211_X1 g_20_26 (.ZN (n_20_26), .A (n_16_28), .B (n_17_28), .C1 (n_13_30), .C2 (n_14_30) );
AOI211_X1 g_22_27 (.ZN (n_22_27), .A (n_18_27), .B (n_19_27), .C1 (n_15_29), .C2 (n_12_29) );
AOI211_X1 g_20_28 (.ZN (n_20_28), .A (n_20_26), .B (n_18_29), .C1 (n_17_28), .C2 (n_11_31) );
AOI211_X1 g_19_30 (.ZN (n_19_30), .A (n_22_27), .B (n_16_28), .C1 (n_19_27), .C2 (n_13_30) );
AOI211_X1 g_18_28 (.ZN (n_18_28), .A (n_20_28), .B (n_18_27), .C1 (n_18_29), .C2 (n_15_29) );
AOI211_X1 g_16_29 (.ZN (n_16_29), .A (n_19_30), .B (n_20_26), .C1 (n_16_28), .C2 (n_17_28) );
AOI211_X1 g_17_31 (.ZN (n_17_31), .A (n_18_28), .B (n_22_27), .C1 (n_18_27), .C2 (n_19_27) );
AOI211_X1 g_15_30 (.ZN (n_15_30), .A (n_16_29), .B (n_20_28), .C1 (n_20_26), .C2 (n_18_29) );
AOI211_X1 g_17_29 (.ZN (n_17_29), .A (n_17_31), .B (n_19_30), .C1 (n_22_27), .C2 (n_16_28) );
AOI211_X1 g_19_28 (.ZN (n_19_28), .A (n_15_30), .B (n_18_28), .C1 (n_20_28), .C2 (n_18_27) );
AOI211_X1 g_21_27 (.ZN (n_21_27), .A (n_17_29), .B (n_16_29), .C1 (n_19_30), .C2 (n_20_26) );
AOI211_X1 g_20_29 (.ZN (n_20_29), .A (n_19_28), .B (n_17_31), .C1 (n_18_28), .C2 (n_22_27) );
AOI211_X1 g_18_30 (.ZN (n_18_30), .A (n_21_27), .B (n_15_30), .C1 (n_16_29), .C2 (n_20_28) );
AOI211_X1 g_16_31 (.ZN (n_16_31), .A (n_20_29), .B (n_17_29), .C1 (n_17_31), .C2 (n_19_30) );
AOI211_X1 g_14_32 (.ZN (n_14_32), .A (n_18_30), .B (n_19_28), .C1 (n_15_30), .C2 (n_18_28) );
AOI211_X1 g_12_33 (.ZN (n_12_33), .A (n_16_31), .B (n_21_27), .C1 (n_17_29), .C2 (n_16_29) );
AOI211_X1 g_13_31 (.ZN (n_13_31), .A (n_14_32), .B (n_20_29), .C1 (n_19_28), .C2 (n_17_31) );
AOI211_X1 g_14_29 (.ZN (n_14_29), .A (n_12_33), .B (n_18_30), .C1 (n_21_27), .C2 (n_15_30) );
AOI211_X1 g_12_30 (.ZN (n_12_30), .A (n_13_31), .B (n_16_31), .C1 (n_20_29), .C2 (n_17_29) );
AOI211_X1 g_10_31 (.ZN (n_10_31), .A (n_14_29), .B (n_14_32), .C1 (n_18_30), .C2 (n_19_28) );
AOI211_X1 g_8_32 (.ZN (n_8_32), .A (n_12_30), .B (n_12_33), .C1 (n_16_31), .C2 (n_21_27) );
AOI211_X1 g_7_34 (.ZN (n_7_34), .A (n_10_31), .B (n_13_31), .C1 (n_14_32), .C2 (n_20_29) );
AOI211_X1 g_9_33 (.ZN (n_9_33), .A (n_8_32), .B (n_14_29), .C1 (n_12_33), .C2 (n_18_30) );
AOI211_X1 g_11_32 (.ZN (n_11_32), .A (n_7_34), .B (n_12_30), .C1 (n_13_31), .C2 (n_16_31) );
AOI211_X1 g_10_34 (.ZN (n_10_34), .A (n_9_33), .B (n_10_31), .C1 (n_14_29), .C2 (n_14_32) );
AOI211_X1 g_8_35 (.ZN (n_8_35), .A (n_11_32), .B (n_8_32), .C1 (n_12_30), .C2 (n_12_33) );
AOI211_X1 g_6_36 (.ZN (n_6_36), .A (n_10_34), .B (n_7_34), .C1 (n_10_31), .C2 (n_13_31) );
AOI211_X1 g_5_38 (.ZN (n_5_38), .A (n_8_35), .B (n_9_33), .C1 (n_8_32), .C2 (n_14_29) );
AOI211_X1 g_3_37 (.ZN (n_3_37), .A (n_6_36), .B (n_11_32), .C1 (n_7_34), .C2 (n_12_30) );
AOI211_X1 g_5_36 (.ZN (n_5_36), .A (n_5_38), .B (n_10_34), .C1 (n_9_33), .C2 (n_10_31) );
AOI211_X1 g_7_35 (.ZN (n_7_35), .A (n_3_37), .B (n_8_35), .C1 (n_11_32), .C2 (n_8_32) );
AOI211_X1 g_9_34 (.ZN (n_9_34), .A (n_5_36), .B (n_6_36), .C1 (n_10_34), .C2 (n_7_34) );
AOI211_X1 g_11_33 (.ZN (n_11_33), .A (n_7_35), .B (n_5_38), .C1 (n_8_35), .C2 (n_9_33) );
AOI211_X1 g_13_32 (.ZN (n_13_32), .A (n_9_34), .B (n_3_37), .C1 (n_6_36), .C2 (n_11_32) );
AOI211_X1 g_15_31 (.ZN (n_15_31), .A (n_11_33), .B (n_5_36), .C1 (n_5_38), .C2 (n_10_34) );
AOI211_X1 g_17_30 (.ZN (n_17_30), .A (n_13_32), .B (n_7_35), .C1 (n_3_37), .C2 (n_8_35) );
AOI211_X1 g_19_29 (.ZN (n_19_29), .A (n_15_31), .B (n_9_34), .C1 (n_5_36), .C2 (n_6_36) );
AOI211_X1 g_20_27 (.ZN (n_20_27), .A (n_17_30), .B (n_11_33), .C1 (n_7_35), .C2 (n_5_38) );
AOI211_X1 g_22_26 (.ZN (n_22_26), .A (n_19_29), .B (n_13_32), .C1 (n_9_34), .C2 (n_3_37) );
AOI211_X1 g_24_25 (.ZN (n_24_25), .A (n_20_27), .B (n_15_31), .C1 (n_11_33), .C2 (n_5_36) );
AOI211_X1 g_26_24 (.ZN (n_26_24), .A (n_22_26), .B (n_17_30), .C1 (n_13_32), .C2 (n_7_35) );
AOI211_X1 g_28_23 (.ZN (n_28_23), .A (n_24_25), .B (n_19_29), .C1 (n_15_31), .C2 (n_9_34) );
AOI211_X1 g_30_22 (.ZN (n_30_22), .A (n_26_24), .B (n_20_27), .C1 (n_17_30), .C2 (n_11_33) );
AOI211_X1 g_32_21 (.ZN (n_32_21), .A (n_28_23), .B (n_22_26), .C1 (n_19_29), .C2 (n_13_32) );
AOI211_X1 g_34_20 (.ZN (n_34_20), .A (n_30_22), .B (n_24_25), .C1 (n_20_27), .C2 (n_15_31) );
AOI211_X1 g_36_19 (.ZN (n_36_19), .A (n_32_21), .B (n_26_24), .C1 (n_22_26), .C2 (n_17_30) );
AOI211_X1 g_38_18 (.ZN (n_38_18), .A (n_34_20), .B (n_28_23), .C1 (n_24_25), .C2 (n_19_29) );
AOI211_X1 g_40_17 (.ZN (n_40_17), .A (n_36_19), .B (n_30_22), .C1 (n_26_24), .C2 (n_20_27) );
AOI211_X1 g_42_16 (.ZN (n_42_16), .A (n_38_18), .B (n_32_21), .C1 (n_28_23), .C2 (n_22_26) );
AOI211_X1 g_44_15 (.ZN (n_44_15), .A (n_40_17), .B (n_34_20), .C1 (n_30_22), .C2 (n_24_25) );
AOI211_X1 g_46_14 (.ZN (n_46_14), .A (n_42_16), .B (n_36_19), .C1 (n_32_21), .C2 (n_26_24) );
AOI211_X1 g_48_13 (.ZN (n_48_13), .A (n_44_15), .B (n_38_18), .C1 (n_34_20), .C2 (n_28_23) );
AOI211_X1 g_50_12 (.ZN (n_50_12), .A (n_46_14), .B (n_40_17), .C1 (n_36_19), .C2 (n_30_22) );
AOI211_X1 g_49_14 (.ZN (n_49_14), .A (n_48_13), .B (n_42_16), .C1 (n_38_18), .C2 (n_32_21) );
AOI211_X1 g_47_13 (.ZN (n_47_13), .A (n_50_12), .B (n_44_15), .C1 (n_40_17), .C2 (n_34_20) );
AOI211_X1 g_49_12 (.ZN (n_49_12), .A (n_49_14), .B (n_46_14), .C1 (n_42_16), .C2 (n_36_19) );
AOI211_X1 g_51_11 (.ZN (n_51_11), .A (n_47_13), .B (n_48_13), .C1 (n_44_15), .C2 (n_38_18) );
AOI211_X1 g_53_10 (.ZN (n_53_10), .A (n_49_12), .B (n_50_12), .C1 (n_46_14), .C2 (n_40_17) );
AOI211_X1 g_55_9 (.ZN (n_55_9), .A (n_51_11), .B (n_49_14), .C1 (n_48_13), .C2 (n_42_16) );
AOI211_X1 g_57_8 (.ZN (n_57_8), .A (n_53_10), .B (n_47_13), .C1 (n_50_12), .C2 (n_44_15) );
AOI211_X1 g_59_7 (.ZN (n_59_7), .A (n_55_9), .B (n_49_12), .C1 (n_49_14), .C2 (n_46_14) );
AOI211_X1 g_61_8 (.ZN (n_61_8), .A (n_57_8), .B (n_51_11), .C1 (n_47_13), .C2 (n_48_13) );
AOI211_X1 g_59_9 (.ZN (n_59_9), .A (n_59_7), .B (n_53_10), .C1 (n_49_12), .C2 (n_50_12) );
AOI211_X1 g_57_10 (.ZN (n_57_10), .A (n_61_8), .B (n_55_9), .C1 (n_51_11), .C2 (n_49_14) );
AOI211_X1 g_55_11 (.ZN (n_55_11), .A (n_59_9), .B (n_57_8), .C1 (n_53_10), .C2 (n_47_13) );
AOI211_X1 g_53_12 (.ZN (n_53_12), .A (n_57_10), .B (n_59_7), .C1 (n_55_9), .C2 (n_49_12) );
AOI211_X1 g_51_13 (.ZN (n_51_13), .A (n_55_11), .B (n_61_8), .C1 (n_57_8), .C2 (n_51_11) );
AOI211_X1 g_50_15 (.ZN (n_50_15), .A (n_53_12), .B (n_59_9), .C1 (n_59_7), .C2 (n_53_10) );
AOI211_X1 g_48_14 (.ZN (n_48_14), .A (n_51_13), .B (n_57_10), .C1 (n_61_8), .C2 (n_55_9) );
AOI211_X1 g_50_13 (.ZN (n_50_13), .A (n_50_15), .B (n_55_11), .C1 (n_59_9), .C2 (n_57_8) );
AOI211_X1 g_52_12 (.ZN (n_52_12), .A (n_48_14), .B (n_53_12), .C1 (n_57_10), .C2 (n_59_7) );
AOI211_X1 g_54_11 (.ZN (n_54_11), .A (n_50_13), .B (n_51_13), .C1 (n_55_11), .C2 (n_61_8) );
AOI211_X1 g_56_10 (.ZN (n_56_10), .A (n_52_12), .B (n_50_15), .C1 (n_53_12), .C2 (n_59_9) );
AOI211_X1 g_58_9 (.ZN (n_58_9), .A (n_54_11), .B (n_48_14), .C1 (n_51_13), .C2 (n_57_10) );
AOI211_X1 g_60_8 (.ZN (n_60_8), .A (n_56_10), .B (n_50_13), .C1 (n_50_15), .C2 (n_55_11) );
AOI211_X1 g_62_9 (.ZN (n_62_9), .A (n_58_9), .B (n_52_12), .C1 (n_48_14), .C2 (n_53_12) );
AOI211_X1 g_60_10 (.ZN (n_60_10), .A (n_60_8), .B (n_54_11), .C1 (n_50_13), .C2 (n_51_13) );
AOI211_X1 g_58_11 (.ZN (n_58_11), .A (n_62_9), .B (n_56_10), .C1 (n_52_12), .C2 (n_50_15) );
AOI211_X1 g_56_12 (.ZN (n_56_12), .A (n_60_10), .B (n_58_9), .C1 (n_54_11), .C2 (n_48_14) );
AOI211_X1 g_54_13 (.ZN (n_54_13), .A (n_58_11), .B (n_60_8), .C1 (n_56_10), .C2 (n_50_13) );
AOI211_X1 g_52_14 (.ZN (n_52_14), .A (n_56_12), .B (n_62_9), .C1 (n_58_9), .C2 (n_52_12) );
AOI211_X1 g_51_16 (.ZN (n_51_16), .A (n_54_13), .B (n_60_10), .C1 (n_60_8), .C2 (n_54_11) );
AOI211_X1 g_50_14 (.ZN (n_50_14), .A (n_52_14), .B (n_58_11), .C1 (n_62_9), .C2 (n_56_10) );
AOI211_X1 g_52_13 (.ZN (n_52_13), .A (n_51_16), .B (n_56_12), .C1 (n_60_10), .C2 (n_58_9) );
AOI211_X1 g_54_12 (.ZN (n_54_12), .A (n_50_14), .B (n_54_13), .C1 (n_58_11), .C2 (n_60_8) );
AOI211_X1 g_56_11 (.ZN (n_56_11), .A (n_52_13), .B (n_52_14), .C1 (n_56_12), .C2 (n_62_9) );
AOI211_X1 g_58_10 (.ZN (n_58_10), .A (n_54_12), .B (n_51_16), .C1 (n_54_13), .C2 (n_60_10) );
AOI211_X1 g_60_9 (.ZN (n_60_9), .A (n_56_11), .B (n_50_14), .C1 (n_52_14), .C2 (n_58_11) );
AOI211_X1 g_62_8 (.ZN (n_62_8), .A (n_58_10), .B (n_52_13), .C1 (n_51_16), .C2 (n_56_12) );
AOI211_X1 g_64_7 (.ZN (n_64_7), .A (n_60_9), .B (n_54_12), .C1 (n_50_14), .C2 (n_54_13) );
AOI211_X1 g_63_9 (.ZN (n_63_9), .A (n_62_8), .B (n_56_11), .C1 (n_52_13), .C2 (n_52_14) );
AOI211_X1 g_61_10 (.ZN (n_61_10), .A (n_64_7), .B (n_58_10), .C1 (n_54_12), .C2 (n_51_16) );
AOI211_X1 g_59_11 (.ZN (n_59_11), .A (n_63_9), .B (n_60_9), .C1 (n_56_11), .C2 (n_50_14) );
AOI211_X1 g_57_12 (.ZN (n_57_12), .A (n_61_10), .B (n_62_8), .C1 (n_58_10), .C2 (n_52_13) );
AOI211_X1 g_55_13 (.ZN (n_55_13), .A (n_59_11), .B (n_64_7), .C1 (n_60_9), .C2 (n_54_12) );
AOI211_X1 g_53_14 (.ZN (n_53_14), .A (n_57_12), .B (n_63_9), .C1 (n_62_8), .C2 (n_56_11) );
AOI211_X1 g_51_15 (.ZN (n_51_15), .A (n_55_13), .B (n_61_10), .C1 (n_64_7), .C2 (n_58_10) );
AOI211_X1 g_49_16 (.ZN (n_49_16), .A (n_53_14), .B (n_59_11), .C1 (n_63_9), .C2 (n_60_9) );
AOI211_X1 g_47_15 (.ZN (n_47_15), .A (n_51_15), .B (n_57_12), .C1 (n_61_10), .C2 (n_62_8) );
AOI211_X1 g_45_14 (.ZN (n_45_14), .A (n_49_16), .B (n_55_13), .C1 (n_59_11), .C2 (n_64_7) );
AOI211_X1 g_43_15 (.ZN (n_43_15), .A (n_47_15), .B (n_53_14), .C1 (n_57_12), .C2 (n_63_9) );
AOI211_X1 g_41_16 (.ZN (n_41_16), .A (n_45_14), .B (n_51_15), .C1 (n_55_13), .C2 (n_61_10) );
AOI211_X1 g_39_17 (.ZN (n_39_17), .A (n_43_15), .B (n_49_16), .C1 (n_53_14), .C2 (n_59_11) );
AOI211_X1 g_37_18 (.ZN (n_37_18), .A (n_41_16), .B (n_47_15), .C1 (n_51_15), .C2 (n_57_12) );
AOI211_X1 g_35_19 (.ZN (n_35_19), .A (n_39_17), .B (n_45_14), .C1 (n_49_16), .C2 (n_55_13) );
AOI211_X1 g_33_20 (.ZN (n_33_20), .A (n_37_18), .B (n_43_15), .C1 (n_47_15), .C2 (n_53_14) );
AOI211_X1 g_32_22 (.ZN (n_32_22), .A (n_35_19), .B (n_41_16), .C1 (n_45_14), .C2 (n_51_15) );
AOI211_X1 g_34_21 (.ZN (n_34_21), .A (n_33_20), .B (n_39_17), .C1 (n_43_15), .C2 (n_49_16) );
AOI211_X1 g_36_20 (.ZN (n_36_20), .A (n_32_22), .B (n_37_18), .C1 (n_41_16), .C2 (n_47_15) );
AOI211_X1 g_38_19 (.ZN (n_38_19), .A (n_34_21), .B (n_35_19), .C1 (n_39_17), .C2 (n_45_14) );
AOI211_X1 g_40_18 (.ZN (n_40_18), .A (n_36_20), .B (n_33_20), .C1 (n_37_18), .C2 (n_43_15) );
AOI211_X1 g_42_17 (.ZN (n_42_17), .A (n_38_19), .B (n_32_22), .C1 (n_35_19), .C2 (n_41_16) );
AOI211_X1 g_44_16 (.ZN (n_44_16), .A (n_40_18), .B (n_34_21), .C1 (n_33_20), .C2 (n_39_17) );
AOI211_X1 g_46_15 (.ZN (n_46_15), .A (n_42_17), .B (n_36_20), .C1 (n_32_22), .C2 (n_37_18) );
AOI211_X1 g_48_16 (.ZN (n_48_16), .A (n_44_16), .B (n_38_19), .C1 (n_34_21), .C2 (n_35_19) );
AOI211_X1 g_46_17 (.ZN (n_46_17), .A (n_46_15), .B (n_40_18), .C1 (n_36_20), .C2 (n_33_20) );
AOI211_X1 g_44_18 (.ZN (n_44_18), .A (n_48_16), .B (n_42_17), .C1 (n_38_19), .C2 (n_32_22) );
AOI211_X1 g_45_16 (.ZN (n_45_16), .A (n_46_17), .B (n_44_16), .C1 (n_40_18), .C2 (n_34_21) );
AOI211_X1 g_43_17 (.ZN (n_43_17), .A (n_44_18), .B (n_46_15), .C1 (n_42_17), .C2 (n_36_20) );
AOI211_X1 g_41_18 (.ZN (n_41_18), .A (n_45_16), .B (n_48_16), .C1 (n_44_16), .C2 (n_38_19) );
AOI211_X1 g_39_19 (.ZN (n_39_19), .A (n_43_17), .B (n_46_17), .C1 (n_46_15), .C2 (n_40_18) );
AOI211_X1 g_37_20 (.ZN (n_37_20), .A (n_41_18), .B (n_44_18), .C1 (n_48_16), .C2 (n_42_17) );
AOI211_X1 g_35_21 (.ZN (n_35_21), .A (n_39_19), .B (n_45_16), .C1 (n_46_17), .C2 (n_44_16) );
AOI211_X1 g_33_22 (.ZN (n_33_22), .A (n_37_20), .B (n_43_17), .C1 (n_44_18), .C2 (n_46_15) );
AOI211_X1 g_31_23 (.ZN (n_31_23), .A (n_35_21), .B (n_41_18), .C1 (n_45_16), .C2 (n_48_16) );
AOI211_X1 g_29_24 (.ZN (n_29_24), .A (n_33_22), .B (n_39_19), .C1 (n_43_17), .C2 (n_46_17) );
AOI211_X1 g_27_25 (.ZN (n_27_25), .A (n_31_23), .B (n_37_20), .C1 (n_41_18), .C2 (n_44_18) );
AOI211_X1 g_25_26 (.ZN (n_25_26), .A (n_29_24), .B (n_35_21), .C1 (n_39_19), .C2 (n_45_16) );
AOI211_X1 g_23_27 (.ZN (n_23_27), .A (n_27_25), .B (n_33_22), .C1 (n_37_20), .C2 (n_43_17) );
AOI211_X1 g_21_28 (.ZN (n_21_28), .A (n_25_26), .B (n_31_23), .C1 (n_35_21), .C2 (n_41_18) );
AOI211_X1 g_20_30 (.ZN (n_20_30), .A (n_23_27), .B (n_29_24), .C1 (n_33_22), .C2 (n_39_19) );
AOI211_X1 g_22_29 (.ZN (n_22_29), .A (n_21_28), .B (n_27_25), .C1 (n_31_23), .C2 (n_37_20) );
AOI211_X1 g_24_28 (.ZN (n_24_28), .A (n_20_30), .B (n_25_26), .C1 (n_29_24), .C2 (n_35_21) );
AOI211_X1 g_26_27 (.ZN (n_26_27), .A (n_22_29), .B (n_23_27), .C1 (n_27_25), .C2 (n_33_22) );
AOI211_X1 g_28_26 (.ZN (n_28_26), .A (n_24_28), .B (n_21_28), .C1 (n_25_26), .C2 (n_31_23) );
AOI211_X1 g_26_25 (.ZN (n_26_25), .A (n_26_27), .B (n_20_30), .C1 (n_23_27), .C2 (n_29_24) );
AOI211_X1 g_28_24 (.ZN (n_28_24), .A (n_28_26), .B (n_22_29), .C1 (n_21_28), .C2 (n_27_25) );
AOI211_X1 g_30_23 (.ZN (n_30_23), .A (n_26_25), .B (n_24_28), .C1 (n_20_30), .C2 (n_25_26) );
AOI211_X1 g_29_25 (.ZN (n_29_25), .A (n_28_24), .B (n_26_27), .C1 (n_22_29), .C2 (n_23_27) );
AOI211_X1 g_31_24 (.ZN (n_31_24), .A (n_30_23), .B (n_28_26), .C1 (n_24_28), .C2 (n_21_28) );
AOI211_X1 g_33_23 (.ZN (n_33_23), .A (n_29_25), .B (n_26_25), .C1 (n_26_27), .C2 (n_20_30) );
AOI211_X1 g_35_22 (.ZN (n_35_22), .A (n_31_24), .B (n_28_24), .C1 (n_28_26), .C2 (n_22_29) );
AOI211_X1 g_37_21 (.ZN (n_37_21), .A (n_33_23), .B (n_30_23), .C1 (n_26_25), .C2 (n_24_28) );
AOI211_X1 g_39_20 (.ZN (n_39_20), .A (n_35_22), .B (n_29_25), .C1 (n_28_24), .C2 (n_26_27) );
AOI211_X1 g_41_19 (.ZN (n_41_19), .A (n_37_21), .B (n_31_24), .C1 (n_30_23), .C2 (n_28_26) );
AOI211_X1 g_43_18 (.ZN (n_43_18), .A (n_39_20), .B (n_33_23), .C1 (n_29_25), .C2 (n_26_25) );
AOI211_X1 g_45_17 (.ZN (n_45_17), .A (n_41_19), .B (n_35_22), .C1 (n_31_24), .C2 (n_28_24) );
AOI211_X1 g_47_16 (.ZN (n_47_16), .A (n_43_18), .B (n_37_21), .C1 (n_33_23), .C2 (n_30_23) );
AOI211_X1 g_49_15 (.ZN (n_49_15), .A (n_45_17), .B (n_39_20), .C1 (n_35_22), .C2 (n_29_25) );
AOI211_X1 g_51_14 (.ZN (n_51_14), .A (n_47_16), .B (n_41_19), .C1 (n_37_21), .C2 (n_31_24) );
AOI211_X1 g_53_13 (.ZN (n_53_13), .A (n_49_15), .B (n_43_18), .C1 (n_39_20), .C2 (n_33_23) );
AOI211_X1 g_55_12 (.ZN (n_55_12), .A (n_51_14), .B (n_45_17), .C1 (n_41_19), .C2 (n_35_22) );
AOI211_X1 g_57_11 (.ZN (n_57_11), .A (n_53_13), .B (n_47_16), .C1 (n_43_18), .C2 (n_37_21) );
AOI211_X1 g_59_10 (.ZN (n_59_10), .A (n_55_12), .B (n_49_15), .C1 (n_45_17), .C2 (n_39_20) );
AOI211_X1 g_58_12 (.ZN (n_58_12), .A (n_57_11), .B (n_51_14), .C1 (n_47_16), .C2 (n_41_19) );
AOI211_X1 g_60_11 (.ZN (n_60_11), .A (n_59_10), .B (n_53_13), .C1 (n_49_15), .C2 (n_43_18) );
AOI211_X1 g_62_10 (.ZN (n_62_10), .A (n_58_12), .B (n_55_12), .C1 (n_51_14), .C2 (n_45_17) );
AOI211_X1 g_64_9 (.ZN (n_64_9), .A (n_60_11), .B (n_57_11), .C1 (n_53_13), .C2 (n_47_16) );
AOI211_X1 g_66_8 (.ZN (n_66_8), .A (n_62_10), .B (n_59_10), .C1 (n_55_12), .C2 (n_49_15) );
AOI211_X1 g_65_10 (.ZN (n_65_10), .A (n_64_9), .B (n_58_12), .C1 (n_57_11), .C2 (n_51_14) );
AOI211_X1 g_63_11 (.ZN (n_63_11), .A (n_66_8), .B (n_60_11), .C1 (n_59_10), .C2 (n_53_13) );
AOI211_X1 g_61_12 (.ZN (n_61_12), .A (n_65_10), .B (n_62_10), .C1 (n_58_12), .C2 (n_55_12) );
AOI211_X1 g_59_13 (.ZN (n_59_13), .A (n_63_11), .B (n_64_9), .C1 (n_60_11), .C2 (n_57_11) );
AOI211_X1 g_57_14 (.ZN (n_57_14), .A (n_61_12), .B (n_66_8), .C1 (n_62_10), .C2 (n_59_10) );
AOI211_X1 g_55_15 (.ZN (n_55_15), .A (n_59_13), .B (n_65_10), .C1 (n_64_9), .C2 (n_58_12) );
AOI211_X1 g_56_13 (.ZN (n_56_13), .A (n_57_14), .B (n_63_11), .C1 (n_66_8), .C2 (n_60_11) );
AOI211_X1 g_54_14 (.ZN (n_54_14), .A (n_55_15), .B (n_61_12), .C1 (n_65_10), .C2 (n_62_10) );
AOI211_X1 g_52_15 (.ZN (n_52_15), .A (n_56_13), .B (n_59_13), .C1 (n_63_11), .C2 (n_64_9) );
AOI211_X1 g_50_16 (.ZN (n_50_16), .A (n_54_14), .B (n_57_14), .C1 (n_61_12), .C2 (n_66_8) );
AOI211_X1 g_48_15 (.ZN (n_48_15), .A (n_52_15), .B (n_55_15), .C1 (n_59_13), .C2 (n_65_10) );
AOI211_X1 g_46_16 (.ZN (n_46_16), .A (n_50_16), .B (n_56_13), .C1 (n_57_14), .C2 (n_63_11) );
AOI211_X1 g_44_17 (.ZN (n_44_17), .A (n_48_15), .B (n_54_14), .C1 (n_55_15), .C2 (n_61_12) );
AOI211_X1 g_42_18 (.ZN (n_42_18), .A (n_46_16), .B (n_52_15), .C1 (n_56_13), .C2 (n_59_13) );
AOI211_X1 g_40_19 (.ZN (n_40_19), .A (n_44_17), .B (n_50_16), .C1 (n_54_14), .C2 (n_57_14) );
AOI211_X1 g_38_20 (.ZN (n_38_20), .A (n_42_18), .B (n_48_15), .C1 (n_52_15), .C2 (n_55_15) );
AOI211_X1 g_36_21 (.ZN (n_36_21), .A (n_40_19), .B (n_46_16), .C1 (n_50_16), .C2 (n_56_13) );
AOI211_X1 g_34_22 (.ZN (n_34_22), .A (n_38_20), .B (n_44_17), .C1 (n_48_15), .C2 (n_54_14) );
AOI211_X1 g_32_23 (.ZN (n_32_23), .A (n_36_21), .B (n_42_18), .C1 (n_46_16), .C2 (n_52_15) );
AOI211_X1 g_30_24 (.ZN (n_30_24), .A (n_34_22), .B (n_40_19), .C1 (n_44_17), .C2 (n_50_16) );
AOI211_X1 g_28_25 (.ZN (n_28_25), .A (n_32_23), .B (n_38_20), .C1 (n_42_18), .C2 (n_48_15) );
AOI211_X1 g_26_26 (.ZN (n_26_26), .A (n_30_24), .B (n_36_21), .C1 (n_40_19), .C2 (n_46_16) );
AOI211_X1 g_24_27 (.ZN (n_24_27), .A (n_28_25), .B (n_34_22), .C1 (n_38_20), .C2 (n_44_17) );
AOI211_X1 g_22_28 (.ZN (n_22_28), .A (n_26_26), .B (n_32_23), .C1 (n_36_21), .C2 (n_42_18) );
AOI211_X1 g_21_30 (.ZN (n_21_30), .A (n_24_27), .B (n_30_24), .C1 (n_34_22), .C2 (n_40_19) );
AOI211_X1 g_23_29 (.ZN (n_23_29), .A (n_22_28), .B (n_28_25), .C1 (n_32_23), .C2 (n_38_20) );
AOI211_X1 g_25_28 (.ZN (n_25_28), .A (n_21_30), .B (n_26_26), .C1 (n_30_24), .C2 (n_36_21) );
AOI211_X1 g_27_27 (.ZN (n_27_27), .A (n_23_29), .B (n_24_27), .C1 (n_28_25), .C2 (n_34_22) );
AOI211_X1 g_29_26 (.ZN (n_29_26), .A (n_25_28), .B (n_22_28), .C1 (n_26_26), .C2 (n_32_23) );
AOI211_X1 g_31_25 (.ZN (n_31_25), .A (n_27_27), .B (n_21_30), .C1 (n_24_27), .C2 (n_30_24) );
AOI211_X1 g_33_24 (.ZN (n_33_24), .A (n_29_26), .B (n_23_29), .C1 (n_22_28), .C2 (n_28_25) );
AOI211_X1 g_35_23 (.ZN (n_35_23), .A (n_31_25), .B (n_25_28), .C1 (n_21_30), .C2 (n_26_26) );
AOI211_X1 g_37_22 (.ZN (n_37_22), .A (n_33_24), .B (n_27_27), .C1 (n_23_29), .C2 (n_24_27) );
AOI211_X1 g_39_21 (.ZN (n_39_21), .A (n_35_23), .B (n_29_26), .C1 (n_25_28), .C2 (n_22_28) );
AOI211_X1 g_41_20 (.ZN (n_41_20), .A (n_37_22), .B (n_31_25), .C1 (n_27_27), .C2 (n_21_30) );
AOI211_X1 g_43_19 (.ZN (n_43_19), .A (n_39_21), .B (n_33_24), .C1 (n_29_26), .C2 (n_23_29) );
AOI211_X1 g_45_18 (.ZN (n_45_18), .A (n_41_20), .B (n_35_23), .C1 (n_31_25), .C2 (n_25_28) );
AOI211_X1 g_47_17 (.ZN (n_47_17), .A (n_43_19), .B (n_37_22), .C1 (n_33_24), .C2 (n_27_27) );
AOI211_X1 g_46_19 (.ZN (n_46_19), .A (n_45_18), .B (n_39_21), .C1 (n_35_23), .C2 (n_29_26) );
AOI211_X1 g_48_18 (.ZN (n_48_18), .A (n_47_17), .B (n_41_20), .C1 (n_37_22), .C2 (n_31_25) );
AOI211_X1 g_50_17 (.ZN (n_50_17), .A (n_46_19), .B (n_43_19), .C1 (n_39_21), .C2 (n_33_24) );
AOI211_X1 g_52_16 (.ZN (n_52_16), .A (n_48_18), .B (n_45_18), .C1 (n_41_20), .C2 (n_35_23) );
AOI211_X1 g_54_15 (.ZN (n_54_15), .A (n_50_17), .B (n_47_17), .C1 (n_43_19), .C2 (n_37_22) );
AOI211_X1 g_56_14 (.ZN (n_56_14), .A (n_52_16), .B (n_46_19), .C1 (n_45_18), .C2 (n_39_21) );
AOI211_X1 g_58_13 (.ZN (n_58_13), .A (n_54_15), .B (n_48_18), .C1 (n_47_17), .C2 (n_41_20) );
AOI211_X1 g_60_12 (.ZN (n_60_12), .A (n_56_14), .B (n_50_17), .C1 (n_46_19), .C2 (n_43_19) );
AOI211_X1 g_62_11 (.ZN (n_62_11), .A (n_58_13), .B (n_52_16), .C1 (n_48_18), .C2 (n_45_18) );
AOI211_X1 g_61_13 (.ZN (n_61_13), .A (n_60_12), .B (n_54_15), .C1 (n_50_17), .C2 (n_47_17) );
AOI211_X1 g_59_12 (.ZN (n_59_12), .A (n_62_11), .B (n_56_14), .C1 (n_52_16), .C2 (n_46_19) );
AOI211_X1 g_61_11 (.ZN (n_61_11), .A (n_61_13), .B (n_58_13), .C1 (n_54_15), .C2 (n_48_18) );
AOI211_X1 g_63_10 (.ZN (n_63_10), .A (n_59_12), .B (n_60_12), .C1 (n_56_14), .C2 (n_50_17) );
AOI211_X1 g_65_9 (.ZN (n_65_9), .A (n_61_11), .B (n_62_11), .C1 (n_58_13), .C2 (n_52_16) );
AOI211_X1 g_66_11 (.ZN (n_66_11), .A (n_63_10), .B (n_61_13), .C1 (n_60_12), .C2 (n_54_15) );
AOI211_X1 g_64_12 (.ZN (n_64_12), .A (n_65_9), .B (n_59_12), .C1 (n_62_11), .C2 (n_56_14) );
AOI211_X1 g_62_13 (.ZN (n_62_13), .A (n_66_11), .B (n_61_11), .C1 (n_61_13), .C2 (n_58_13) );
AOI211_X1 g_60_14 (.ZN (n_60_14), .A (n_64_12), .B (n_63_10), .C1 (n_59_12), .C2 (n_60_12) );
AOI211_X1 g_58_15 (.ZN (n_58_15), .A (n_62_13), .B (n_65_9), .C1 (n_61_11), .C2 (n_62_11) );
AOI211_X1 g_57_13 (.ZN (n_57_13), .A (n_60_14), .B (n_66_11), .C1 (n_63_10), .C2 (n_61_13) );
AOI211_X1 g_55_14 (.ZN (n_55_14), .A (n_58_15), .B (n_64_12), .C1 (n_65_9), .C2 (n_59_12) );
AOI211_X1 g_53_15 (.ZN (n_53_15), .A (n_57_13), .B (n_62_13), .C1 (n_66_11), .C2 (n_61_11) );
AOI211_X1 g_52_17 (.ZN (n_52_17), .A (n_55_14), .B (n_60_14), .C1 (n_64_12), .C2 (n_63_10) );
AOI211_X1 g_54_16 (.ZN (n_54_16), .A (n_53_15), .B (n_58_15), .C1 (n_62_13), .C2 (n_65_9) );
AOI211_X1 g_56_15 (.ZN (n_56_15), .A (n_52_17), .B (n_57_13), .C1 (n_60_14), .C2 (n_66_11) );
AOI211_X1 g_58_14 (.ZN (n_58_14), .A (n_54_16), .B (n_55_14), .C1 (n_58_15), .C2 (n_64_12) );
AOI211_X1 g_60_13 (.ZN (n_60_13), .A (n_56_15), .B (n_53_15), .C1 (n_57_13), .C2 (n_62_13) );
AOI211_X1 g_62_12 (.ZN (n_62_12), .A (n_58_14), .B (n_52_17), .C1 (n_55_14), .C2 (n_60_14) );
AOI211_X1 g_64_11 (.ZN (n_64_11), .A (n_60_13), .B (n_54_16), .C1 (n_53_15), .C2 (n_58_15) );
AOI211_X1 g_66_10 (.ZN (n_66_10), .A (n_62_12), .B (n_56_15), .C1 (n_52_17), .C2 (n_57_13) );
AOI211_X1 g_68_9 (.ZN (n_68_9), .A (n_64_11), .B (n_58_14), .C1 (n_54_16), .C2 (n_55_14) );
AOI211_X1 g_70_10 (.ZN (n_70_10), .A (n_66_10), .B (n_60_13), .C1 (n_56_15), .C2 (n_53_15) );
AOI211_X1 g_68_11 (.ZN (n_68_11), .A (n_68_9), .B (n_62_12), .C1 (n_58_14), .C2 (n_52_17) );
AOI211_X1 g_70_12 (.ZN (n_70_12), .A (n_70_10), .B (n_64_11), .C1 (n_60_13), .C2 (n_54_16) );
AOI211_X1 g_72_13 (.ZN (n_72_13), .A (n_68_11), .B (n_66_10), .C1 (n_62_12), .C2 (n_56_15) );
AOI211_X1 g_73_11 (.ZN (n_73_11), .A (n_70_12), .B (n_68_9), .C1 (n_64_11), .C2 (n_58_14) );
AOI211_X1 g_74_13 (.ZN (n_74_13), .A (n_72_13), .B (n_70_10), .C1 (n_66_10), .C2 (n_60_13) );
AOI211_X1 g_72_14 (.ZN (n_72_14), .A (n_73_11), .B (n_68_11), .C1 (n_68_9), .C2 (n_62_12) );
AOI211_X1 g_71_12 (.ZN (n_71_12), .A (n_74_13), .B (n_70_12), .C1 (n_70_10), .C2 (n_64_11) );
AOI211_X1 g_69_11 (.ZN (n_69_11), .A (n_72_14), .B (n_72_13), .C1 (n_68_11), .C2 (n_66_10) );
AOI211_X1 g_67_10 (.ZN (n_67_10), .A (n_71_12), .B (n_73_11), .C1 (n_70_12), .C2 (n_68_9) );
AOI211_X1 g_65_11 (.ZN (n_65_11), .A (n_69_11), .B (n_74_13), .C1 (n_72_13), .C2 (n_70_10) );
AOI211_X1 g_63_12 (.ZN (n_63_12), .A (n_67_10), .B (n_72_14), .C1 (n_73_11), .C2 (n_68_11) );
AOI211_X1 g_62_14 (.ZN (n_62_14), .A (n_65_11), .B (n_71_12), .C1 (n_74_13), .C2 (n_70_12) );
AOI211_X1 g_64_13 (.ZN (n_64_13), .A (n_63_12), .B (n_69_11), .C1 (n_72_14), .C2 (n_72_13) );
AOI211_X1 g_66_12 (.ZN (n_66_12), .A (n_62_14), .B (n_67_10), .C1 (n_71_12), .C2 (n_73_11) );
AOI211_X1 g_68_13 (.ZN (n_68_13), .A (n_64_13), .B (n_65_11), .C1 (n_69_11), .C2 (n_74_13) );
AOI211_X1 g_67_11 (.ZN (n_67_11), .A (n_66_12), .B (n_63_12), .C1 (n_67_10), .C2 (n_72_14) );
AOI211_X1 g_69_12 (.ZN (n_69_12), .A (n_68_13), .B (n_62_14), .C1 (n_65_11), .C2 (n_71_12) );
AOI211_X1 g_70_14 (.ZN (n_70_14), .A (n_67_11), .B (n_64_13), .C1 (n_63_12), .C2 (n_69_11) );
AOI211_X1 g_71_16 (.ZN (n_71_16), .A (n_69_12), .B (n_66_12), .C1 (n_62_14), .C2 (n_67_10) );
AOI211_X1 g_73_15 (.ZN (n_73_15), .A (n_70_14), .B (n_68_13), .C1 (n_64_13), .C2 (n_65_11) );
AOI211_X1 g_75_14 (.ZN (n_75_14), .A (n_71_16), .B (n_67_11), .C1 (n_66_12), .C2 (n_63_12) );
AOI211_X1 g_73_13 (.ZN (n_73_13), .A (n_73_15), .B (n_69_12), .C1 (n_68_13), .C2 (n_62_14) );
AOI211_X1 g_75_12 (.ZN (n_75_12), .A (n_75_14), .B (n_70_14), .C1 (n_67_11), .C2 (n_64_13) );
AOI211_X1 g_77_11 (.ZN (n_77_11), .A (n_73_13), .B (n_71_16), .C1 (n_69_12), .C2 (n_66_12) );
AOI211_X1 g_78_13 (.ZN (n_78_13), .A (n_75_12), .B (n_73_15), .C1 (n_70_14), .C2 (n_68_13) );
AOI211_X1 g_76_14 (.ZN (n_76_14), .A (n_77_11), .B (n_75_14), .C1 (n_71_16), .C2 (n_67_11) );
AOI211_X1 g_74_15 (.ZN (n_74_15), .A (n_78_13), .B (n_73_13), .C1 (n_73_15), .C2 (n_69_12) );
AOI211_X1 g_72_16 (.ZN (n_72_16), .A (n_76_14), .B (n_75_12), .C1 (n_75_14), .C2 (n_70_14) );
AOI211_X1 g_71_14 (.ZN (n_71_14), .A (n_74_15), .B (n_77_11), .C1 (n_73_13), .C2 (n_71_16) );
AOI211_X1 g_69_13 (.ZN (n_69_13), .A (n_72_16), .B (n_78_13), .C1 (n_75_12), .C2 (n_73_15) );
AOI211_X1 g_67_12 (.ZN (n_67_12), .A (n_71_14), .B (n_76_14), .C1 (n_77_11), .C2 (n_75_14) );
AOI211_X1 g_65_13 (.ZN (n_65_13), .A (n_69_13), .B (n_74_15), .C1 (n_78_13), .C2 (n_73_13) );
AOI211_X1 g_63_14 (.ZN (n_63_14), .A (n_67_12), .B (n_72_16), .C1 (n_76_14), .C2 (n_75_12) );
AOI211_X1 g_61_15 (.ZN (n_61_15), .A (n_65_13), .B (n_71_14), .C1 (n_74_15), .C2 (n_77_11) );
AOI211_X1 g_59_14 (.ZN (n_59_14), .A (n_63_14), .B (n_69_13), .C1 (n_72_16), .C2 (n_78_13) );
AOI211_X1 g_57_15 (.ZN (n_57_15), .A (n_61_15), .B (n_67_12), .C1 (n_71_14), .C2 (n_76_14) );
AOI211_X1 g_55_16 (.ZN (n_55_16), .A (n_59_14), .B (n_65_13), .C1 (n_69_13), .C2 (n_74_15) );
AOI211_X1 g_53_17 (.ZN (n_53_17), .A (n_57_15), .B (n_63_14), .C1 (n_67_12), .C2 (n_72_16) );
AOI211_X1 g_51_18 (.ZN (n_51_18), .A (n_55_16), .B (n_61_15), .C1 (n_65_13), .C2 (n_71_14) );
AOI211_X1 g_49_17 (.ZN (n_49_17), .A (n_53_17), .B (n_59_14), .C1 (n_63_14), .C2 (n_69_13) );
AOI211_X1 g_47_18 (.ZN (n_47_18), .A (n_51_18), .B (n_57_15), .C1 (n_61_15), .C2 (n_67_12) );
AOI211_X1 g_45_19 (.ZN (n_45_19), .A (n_49_17), .B (n_55_16), .C1 (n_59_14), .C2 (n_65_13) );
AOI211_X1 g_43_20 (.ZN (n_43_20), .A (n_47_18), .B (n_53_17), .C1 (n_57_15), .C2 (n_63_14) );
AOI211_X1 g_41_21 (.ZN (n_41_21), .A (n_45_19), .B (n_51_18), .C1 (n_55_16), .C2 (n_61_15) );
AOI211_X1 g_42_19 (.ZN (n_42_19), .A (n_43_20), .B (n_49_17), .C1 (n_53_17), .C2 (n_59_14) );
AOI211_X1 g_40_20 (.ZN (n_40_20), .A (n_41_21), .B (n_47_18), .C1 (n_51_18), .C2 (n_57_15) );
AOI211_X1 g_38_21 (.ZN (n_38_21), .A (n_42_19), .B (n_45_19), .C1 (n_49_17), .C2 (n_55_16) );
AOI211_X1 g_36_22 (.ZN (n_36_22), .A (n_40_20), .B (n_43_20), .C1 (n_47_18), .C2 (n_53_17) );
AOI211_X1 g_34_23 (.ZN (n_34_23), .A (n_38_21), .B (n_41_21), .C1 (n_45_19), .C2 (n_51_18) );
AOI211_X1 g_32_24 (.ZN (n_32_24), .A (n_36_22), .B (n_42_19), .C1 (n_43_20), .C2 (n_49_17) );
AOI211_X1 g_30_25 (.ZN (n_30_25), .A (n_34_23), .B (n_40_20), .C1 (n_41_21), .C2 (n_47_18) );
AOI211_X1 g_32_26 (.ZN (n_32_26), .A (n_32_24), .B (n_38_21), .C1 (n_42_19), .C2 (n_45_19) );
AOI211_X1 g_34_25 (.ZN (n_34_25), .A (n_30_25), .B (n_36_22), .C1 (n_40_20), .C2 (n_43_20) );
AOI211_X1 g_36_24 (.ZN (n_36_24), .A (n_32_26), .B (n_34_23), .C1 (n_38_21), .C2 (n_41_21) );
AOI211_X1 g_38_23 (.ZN (n_38_23), .A (n_34_25), .B (n_32_24), .C1 (n_36_22), .C2 (n_42_19) );
AOI211_X1 g_40_22 (.ZN (n_40_22), .A (n_36_24), .B (n_30_25), .C1 (n_34_23), .C2 (n_40_20) );
AOI211_X1 g_42_21 (.ZN (n_42_21), .A (n_38_23), .B (n_32_26), .C1 (n_32_24), .C2 (n_38_21) );
AOI211_X1 g_44_20 (.ZN (n_44_20), .A (n_40_22), .B (n_34_25), .C1 (n_30_25), .C2 (n_36_22) );
AOI211_X1 g_43_22 (.ZN (n_43_22), .A (n_42_21), .B (n_36_24), .C1 (n_32_26), .C2 (n_34_23) );
AOI211_X1 g_42_20 (.ZN (n_42_20), .A (n_44_20), .B (n_38_23), .C1 (n_34_25), .C2 (n_32_24) );
AOI211_X1 g_44_19 (.ZN (n_44_19), .A (n_43_22), .B (n_40_22), .C1 (n_36_24), .C2 (n_30_25) );
AOI211_X1 g_46_18 (.ZN (n_46_18), .A (n_42_20), .B (n_42_21), .C1 (n_38_23), .C2 (n_32_26) );
AOI211_X1 g_48_17 (.ZN (n_48_17), .A (n_44_19), .B (n_44_20), .C1 (n_40_22), .C2 (n_34_25) );
AOI211_X1 g_49_19 (.ZN (n_49_19), .A (n_46_18), .B (n_43_22), .C1 (n_42_21), .C2 (n_36_24) );
AOI211_X1 g_47_20 (.ZN (n_47_20), .A (n_48_17), .B (n_42_20), .C1 (n_44_20), .C2 (n_38_23) );
AOI211_X1 g_45_21 (.ZN (n_45_21), .A (n_49_19), .B (n_44_19), .C1 (n_43_22), .C2 (n_40_22) );
AOI211_X1 g_44_23 (.ZN (n_44_23), .A (n_47_20), .B (n_46_18), .C1 (n_42_20), .C2 (n_42_21) );
AOI211_X1 g_43_21 (.ZN (n_43_21), .A (n_45_21), .B (n_48_17), .C1 (n_44_19), .C2 (n_44_20) );
AOI211_X1 g_45_20 (.ZN (n_45_20), .A (n_44_23), .B (n_49_19), .C1 (n_46_18), .C2 (n_43_22) );
AOI211_X1 g_47_19 (.ZN (n_47_19), .A (n_43_21), .B (n_47_20), .C1 (n_48_17), .C2 (n_42_20) );
AOI211_X1 g_49_18 (.ZN (n_49_18), .A (n_45_20), .B (n_45_21), .C1 (n_49_19), .C2 (n_44_19) );
AOI211_X1 g_51_17 (.ZN (n_51_17), .A (n_47_19), .B (n_44_23), .C1 (n_47_20), .C2 (n_46_18) );
AOI211_X1 g_53_16 (.ZN (n_53_16), .A (n_49_18), .B (n_43_21), .C1 (n_45_21), .C2 (n_48_17) );
AOI211_X1 g_52_18 (.ZN (n_52_18), .A (n_51_17), .B (n_45_20), .C1 (n_44_23), .C2 (n_49_19) );
AOI211_X1 g_54_17 (.ZN (n_54_17), .A (n_53_16), .B (n_47_19), .C1 (n_43_21), .C2 (n_47_20) );
AOI211_X1 g_56_16 (.ZN (n_56_16), .A (n_52_18), .B (n_49_18), .C1 (n_45_20), .C2 (n_45_21) );
AOI211_X1 g_55_18 (.ZN (n_55_18), .A (n_54_17), .B (n_51_17), .C1 (n_47_19), .C2 (n_44_23) );
AOI211_X1 g_57_17 (.ZN (n_57_17), .A (n_56_16), .B (n_53_16), .C1 (n_49_18), .C2 (n_43_21) );
AOI211_X1 g_59_16 (.ZN (n_59_16), .A (n_55_18), .B (n_52_18), .C1 (n_51_17), .C2 (n_45_20) );
AOI211_X1 g_58_18 (.ZN (n_58_18), .A (n_57_17), .B (n_54_17), .C1 (n_53_16), .C2 (n_47_19) );
AOI211_X1 g_57_16 (.ZN (n_57_16), .A (n_59_16), .B (n_56_16), .C1 (n_52_18), .C2 (n_49_18) );
AOI211_X1 g_59_15 (.ZN (n_59_15), .A (n_58_18), .B (n_55_18), .C1 (n_54_17), .C2 (n_51_17) );
AOI211_X1 g_61_14 (.ZN (n_61_14), .A (n_57_16), .B (n_57_17), .C1 (n_56_16), .C2 (n_53_16) );
AOI211_X1 g_63_13 (.ZN (n_63_13), .A (n_59_15), .B (n_59_16), .C1 (n_55_18), .C2 (n_52_18) );
AOI211_X1 g_65_12 (.ZN (n_65_12), .A (n_61_14), .B (n_58_18), .C1 (n_57_17), .C2 (n_54_17) );
AOI211_X1 g_66_14 (.ZN (n_66_14), .A (n_63_13), .B (n_57_16), .C1 (n_59_16), .C2 (n_56_16) );
AOI211_X1 g_64_15 (.ZN (n_64_15), .A (n_65_12), .B (n_59_15), .C1 (n_58_18), .C2 (n_55_18) );
AOI211_X1 g_62_16 (.ZN (n_62_16), .A (n_66_14), .B (n_61_14), .C1 (n_57_16), .C2 (n_57_17) );
AOI211_X1 g_60_15 (.ZN (n_60_15), .A (n_64_15), .B (n_63_13), .C1 (n_59_15), .C2 (n_59_16) );
AOI211_X1 g_58_16 (.ZN (n_58_16), .A (n_62_16), .B (n_65_12), .C1 (n_61_14), .C2 (n_58_18) );
AOI211_X1 g_56_17 (.ZN (n_56_17), .A (n_60_15), .B (n_66_14), .C1 (n_63_13), .C2 (n_57_16) );
AOI211_X1 g_54_18 (.ZN (n_54_18), .A (n_58_16), .B (n_64_15), .C1 (n_65_12), .C2 (n_59_15) );
AOI211_X1 g_52_19 (.ZN (n_52_19), .A (n_56_17), .B (n_62_16), .C1 (n_66_14), .C2 (n_61_14) );
AOI211_X1 g_50_18 (.ZN (n_50_18), .A (n_54_18), .B (n_60_15), .C1 (n_64_15), .C2 (n_63_13) );
AOI211_X1 g_48_19 (.ZN (n_48_19), .A (n_52_19), .B (n_58_16), .C1 (n_62_16), .C2 (n_65_12) );
AOI211_X1 g_46_20 (.ZN (n_46_20), .A (n_50_18), .B (n_56_17), .C1 (n_60_15), .C2 (n_66_14) );
AOI211_X1 g_44_21 (.ZN (n_44_21), .A (n_48_19), .B (n_54_18), .C1 (n_58_16), .C2 (n_64_15) );
AOI211_X1 g_42_22 (.ZN (n_42_22), .A (n_46_20), .B (n_52_19), .C1 (n_56_17), .C2 (n_62_16) );
AOI211_X1 g_40_21 (.ZN (n_40_21), .A (n_44_21), .B (n_50_18), .C1 (n_54_18), .C2 (n_60_15) );
AOI211_X1 g_38_22 (.ZN (n_38_22), .A (n_42_22), .B (n_48_19), .C1 (n_52_19), .C2 (n_58_16) );
AOI211_X1 g_36_23 (.ZN (n_36_23), .A (n_40_21), .B (n_46_20), .C1 (n_50_18), .C2 (n_56_17) );
AOI211_X1 g_34_24 (.ZN (n_34_24), .A (n_38_22), .B (n_44_21), .C1 (n_48_19), .C2 (n_54_18) );
AOI211_X1 g_32_25 (.ZN (n_32_25), .A (n_36_23), .B (n_42_22), .C1 (n_46_20), .C2 (n_52_19) );
AOI211_X1 g_30_26 (.ZN (n_30_26), .A (n_34_24), .B (n_40_21), .C1 (n_44_21), .C2 (n_50_18) );
AOI211_X1 g_28_27 (.ZN (n_28_27), .A (n_32_25), .B (n_38_22), .C1 (n_42_22), .C2 (n_48_19) );
AOI211_X1 g_26_28 (.ZN (n_26_28), .A (n_30_26), .B (n_36_23), .C1 (n_40_21), .C2 (n_46_20) );
AOI211_X1 g_27_26 (.ZN (n_27_26), .A (n_28_27), .B (n_34_24), .C1 (n_38_22), .C2 (n_44_21) );
AOI211_X1 g_25_27 (.ZN (n_25_27), .A (n_26_28), .B (n_32_25), .C1 (n_36_23), .C2 (n_42_22) );
AOI211_X1 g_23_28 (.ZN (n_23_28), .A (n_27_26), .B (n_30_26), .C1 (n_34_24), .C2 (n_40_21) );
AOI211_X1 g_21_29 (.ZN (n_21_29), .A (n_25_27), .B (n_28_27), .C1 (n_32_25), .C2 (n_38_22) );
AOI211_X1 g_20_31 (.ZN (n_20_31), .A (n_23_28), .B (n_26_28), .C1 (n_30_26), .C2 (n_36_23) );
AOI211_X1 g_22_30 (.ZN (n_22_30), .A (n_21_29), .B (n_27_26), .C1 (n_28_27), .C2 (n_34_24) );
AOI211_X1 g_24_29 (.ZN (n_24_29), .A (n_20_31), .B (n_25_27), .C1 (n_26_28), .C2 (n_32_25) );
AOI211_X1 g_23_31 (.ZN (n_23_31), .A (n_22_30), .B (n_23_28), .C1 (n_27_26), .C2 (n_30_26) );
AOI211_X1 g_25_30 (.ZN (n_25_30), .A (n_24_29), .B (n_21_29), .C1 (n_25_27), .C2 (n_28_27) );
AOI211_X1 g_27_29 (.ZN (n_27_29), .A (n_23_31), .B (n_20_31), .C1 (n_23_28), .C2 (n_26_28) );
AOI211_X1 g_29_28 (.ZN (n_29_28), .A (n_25_30), .B (n_22_30), .C1 (n_21_29), .C2 (n_27_26) );
AOI211_X1 g_31_27 (.ZN (n_31_27), .A (n_27_29), .B (n_24_29), .C1 (n_20_31), .C2 (n_25_27) );
AOI211_X1 g_33_26 (.ZN (n_33_26), .A (n_29_28), .B (n_23_31), .C1 (n_22_30), .C2 (n_23_28) );
AOI211_X1 g_35_25 (.ZN (n_35_25), .A (n_31_27), .B (n_25_30), .C1 (n_24_29), .C2 (n_21_29) );
AOI211_X1 g_37_24 (.ZN (n_37_24), .A (n_33_26), .B (n_27_29), .C1 (n_23_31), .C2 (n_20_31) );
AOI211_X1 g_39_23 (.ZN (n_39_23), .A (n_35_25), .B (n_29_28), .C1 (n_25_30), .C2 (n_22_30) );
AOI211_X1 g_41_22 (.ZN (n_41_22), .A (n_37_24), .B (n_31_27), .C1 (n_27_29), .C2 (n_24_29) );
AOI211_X1 g_42_24 (.ZN (n_42_24), .A (n_39_23), .B (n_33_26), .C1 (n_29_28), .C2 (n_23_31) );
AOI211_X1 g_40_23 (.ZN (n_40_23), .A (n_41_22), .B (n_35_25), .C1 (n_31_27), .C2 (n_25_30) );
AOI211_X1 g_38_24 (.ZN (n_38_24), .A (n_42_24), .B (n_37_24), .C1 (n_33_26), .C2 (n_27_29) );
AOI211_X1 g_39_22 (.ZN (n_39_22), .A (n_40_23), .B (n_39_23), .C1 (n_35_25), .C2 (n_29_28) );
AOI211_X1 g_37_23 (.ZN (n_37_23), .A (n_38_24), .B (n_41_22), .C1 (n_37_24), .C2 (n_31_27) );
AOI211_X1 g_35_24 (.ZN (n_35_24), .A (n_39_22), .B (n_42_24), .C1 (n_39_23), .C2 (n_33_26) );
AOI211_X1 g_33_25 (.ZN (n_33_25), .A (n_37_23), .B (n_40_23), .C1 (n_41_22), .C2 (n_35_25) );
AOI211_X1 g_31_26 (.ZN (n_31_26), .A (n_35_24), .B (n_38_24), .C1 (n_42_24), .C2 (n_37_24) );
AOI211_X1 g_29_27 (.ZN (n_29_27), .A (n_33_25), .B (n_39_22), .C1 (n_40_23), .C2 (n_39_23) );
AOI211_X1 g_27_28 (.ZN (n_27_28), .A (n_31_26), .B (n_37_23), .C1 (n_38_24), .C2 (n_41_22) );
AOI211_X1 g_25_29 (.ZN (n_25_29), .A (n_29_27), .B (n_35_24), .C1 (n_39_22), .C2 (n_42_24) );
AOI211_X1 g_23_30 (.ZN (n_23_30), .A (n_27_28), .B (n_33_25), .C1 (n_37_23), .C2 (n_40_23) );
AOI211_X1 g_21_31 (.ZN (n_21_31), .A (n_25_29), .B (n_31_26), .C1 (n_35_24), .C2 (n_38_24) );
AOI211_X1 g_19_32 (.ZN (n_19_32), .A (n_23_30), .B (n_29_27), .C1 (n_33_25), .C2 (n_39_22) );
AOI211_X1 g_17_33 (.ZN (n_17_33), .A (n_21_31), .B (n_27_28), .C1 (n_31_26), .C2 (n_37_23) );
AOI211_X1 g_18_31 (.ZN (n_18_31), .A (n_19_32), .B (n_25_29), .C1 (n_29_27), .C2 (n_35_24) );
AOI211_X1 g_16_30 (.ZN (n_16_30), .A (n_17_33), .B (n_23_30), .C1 (n_27_28), .C2 (n_33_25) );
AOI211_X1 g_15_32 (.ZN (n_15_32), .A (n_18_31), .B (n_21_31), .C1 (n_25_29), .C2 (n_31_26) );
AOI211_X1 g_13_33 (.ZN (n_13_33), .A (n_16_30), .B (n_19_32), .C1 (n_23_30), .C2 (n_29_27) );
AOI211_X1 g_14_31 (.ZN (n_14_31), .A (n_15_32), .B (n_17_33), .C1 (n_21_31), .C2 (n_27_28) );
AOI211_X1 g_12_32 (.ZN (n_12_32), .A (n_13_33), .B (n_18_31), .C1 (n_19_32), .C2 (n_25_29) );
AOI211_X1 g_10_33 (.ZN (n_10_33), .A (n_14_31), .B (n_16_30), .C1 (n_17_33), .C2 (n_23_30) );
AOI211_X1 g_9_35 (.ZN (n_9_35), .A (n_12_32), .B (n_15_32), .C1 (n_18_31), .C2 (n_21_31) );
AOI211_X1 g_11_34 (.ZN (n_11_34), .A (n_10_33), .B (n_13_33), .C1 (n_16_30), .C2 (n_19_32) );
AOI211_X1 g_10_36 (.ZN (n_10_36), .A (n_9_35), .B (n_14_31), .C1 (n_15_32), .C2 (n_17_33) );
AOI211_X1 g_12_35 (.ZN (n_12_35), .A (n_11_34), .B (n_12_32), .C1 (n_13_33), .C2 (n_18_31) );
AOI211_X1 g_14_34 (.ZN (n_14_34), .A (n_10_36), .B (n_10_33), .C1 (n_14_31), .C2 (n_16_30) );
AOI211_X1 g_16_33 (.ZN (n_16_33), .A (n_12_35), .B (n_9_35), .C1 (n_12_32), .C2 (n_15_32) );
AOI211_X1 g_18_32 (.ZN (n_18_32), .A (n_14_34), .B (n_11_34), .C1 (n_10_33), .C2 (n_13_33) );
AOI211_X1 g_19_34 (.ZN (n_19_34), .A (n_16_33), .B (n_10_36), .C1 (n_9_35), .C2 (n_14_31) );
AOI211_X1 g_20_32 (.ZN (n_20_32), .A (n_18_32), .B (n_12_35), .C1 (n_11_34), .C2 (n_12_32) );
AOI211_X1 g_22_31 (.ZN (n_22_31), .A (n_19_34), .B (n_14_34), .C1 (n_10_36), .C2 (n_10_33) );
AOI211_X1 g_24_30 (.ZN (n_24_30), .A (n_20_32), .B (n_16_33), .C1 (n_12_35), .C2 (n_9_35) );
AOI211_X1 g_26_29 (.ZN (n_26_29), .A (n_22_31), .B (n_18_32), .C1 (n_14_34), .C2 (n_11_34) );
AOI211_X1 g_28_28 (.ZN (n_28_28), .A (n_24_30), .B (n_19_34), .C1 (n_16_33), .C2 (n_10_36) );
AOI211_X1 g_30_27 (.ZN (n_30_27), .A (n_26_29), .B (n_20_32), .C1 (n_18_32), .C2 (n_12_35) );
AOI211_X1 g_29_29 (.ZN (n_29_29), .A (n_28_28), .B (n_22_31), .C1 (n_19_34), .C2 (n_14_34) );
AOI211_X1 g_31_28 (.ZN (n_31_28), .A (n_30_27), .B (n_24_30), .C1 (n_20_32), .C2 (n_16_33) );
AOI211_X1 g_33_27 (.ZN (n_33_27), .A (n_29_29), .B (n_26_29), .C1 (n_22_31), .C2 (n_18_32) );
AOI211_X1 g_35_26 (.ZN (n_35_26), .A (n_31_28), .B (n_28_28), .C1 (n_24_30), .C2 (n_19_34) );
AOI211_X1 g_37_25 (.ZN (n_37_25), .A (n_33_27), .B (n_30_27), .C1 (n_26_29), .C2 (n_20_32) );
AOI211_X1 g_39_24 (.ZN (n_39_24), .A (n_35_26), .B (n_29_29), .C1 (n_28_28), .C2 (n_22_31) );
AOI211_X1 g_41_23 (.ZN (n_41_23), .A (n_37_25), .B (n_31_28), .C1 (n_30_27), .C2 (n_24_30) );
AOI211_X1 g_40_25 (.ZN (n_40_25), .A (n_39_24), .B (n_33_27), .C1 (n_29_29), .C2 (n_26_29) );
AOI211_X1 g_38_26 (.ZN (n_38_26), .A (n_41_23), .B (n_35_26), .C1 (n_31_28), .C2 (n_28_28) );
AOI211_X1 g_36_25 (.ZN (n_36_25), .A (n_40_25), .B (n_37_25), .C1 (n_33_27), .C2 (n_30_27) );
AOI211_X1 g_34_26 (.ZN (n_34_26), .A (n_38_26), .B (n_39_24), .C1 (n_35_26), .C2 (n_29_29) );
AOI211_X1 g_32_27 (.ZN (n_32_27), .A (n_36_25), .B (n_41_23), .C1 (n_37_25), .C2 (n_31_28) );
AOI211_X1 g_30_28 (.ZN (n_30_28), .A (n_34_26), .B (n_40_25), .C1 (n_39_24), .C2 (n_33_27) );
AOI211_X1 g_28_29 (.ZN (n_28_29), .A (n_32_27), .B (n_38_26), .C1 (n_41_23), .C2 (n_35_26) );
AOI211_X1 g_26_30 (.ZN (n_26_30), .A (n_30_28), .B (n_36_25), .C1 (n_40_25), .C2 (n_37_25) );
AOI211_X1 g_24_31 (.ZN (n_24_31), .A (n_28_29), .B (n_34_26), .C1 (n_38_26), .C2 (n_39_24) );
AOI211_X1 g_22_32 (.ZN (n_22_32), .A (n_26_30), .B (n_32_27), .C1 (n_36_25), .C2 (n_41_23) );
AOI211_X1 g_20_33 (.ZN (n_20_33), .A (n_24_31), .B (n_30_28), .C1 (n_34_26), .C2 (n_40_25) );
AOI211_X1 g_19_31 (.ZN (n_19_31), .A (n_22_32), .B (n_28_29), .C1 (n_32_27), .C2 (n_38_26) );
AOI211_X1 g_17_32 (.ZN (n_17_32), .A (n_20_33), .B (n_26_30), .C1 (n_30_28), .C2 (n_36_25) );
AOI211_X1 g_15_33 (.ZN (n_15_33), .A (n_19_31), .B (n_24_31), .C1 (n_28_29), .C2 (n_34_26) );
AOI211_X1 g_13_34 (.ZN (n_13_34), .A (n_17_32), .B (n_22_32), .C1 (n_26_30), .C2 (n_32_27) );
AOI211_X1 g_11_35 (.ZN (n_11_35), .A (n_15_33), .B (n_20_33), .C1 (n_24_31), .C2 (n_30_28) );
AOI211_X1 g_9_36 (.ZN (n_9_36), .A (n_13_34), .B (n_19_31), .C1 (n_22_32), .C2 (n_28_29) );
AOI211_X1 g_7_37 (.ZN (n_7_37), .A (n_11_35), .B (n_17_32), .C1 (n_20_33), .C2 (n_26_30) );
AOI211_X1 g_6_39 (.ZN (n_6_39), .A (n_9_36), .B (n_15_33), .C1 (n_19_31), .C2 (n_24_31) );
AOI211_X1 g_4_38 (.ZN (n_4_38), .A (n_7_37), .B (n_13_34), .C1 (n_17_32), .C2 (n_22_32) );
AOI211_X1 g_6_37 (.ZN (n_6_37), .A (n_6_39), .B (n_11_35), .C1 (n_15_33), .C2 (n_20_33) );
AOI211_X1 g_8_36 (.ZN (n_8_36), .A (n_4_38), .B (n_9_36), .C1 (n_13_34), .C2 (n_19_31) );
AOI211_X1 g_10_35 (.ZN (n_10_35), .A (n_6_37), .B (n_7_37), .C1 (n_11_35), .C2 (n_17_32) );
AOI211_X1 g_12_34 (.ZN (n_12_34), .A (n_8_36), .B (n_6_39), .C1 (n_9_36), .C2 (n_15_33) );
AOI211_X1 g_14_33 (.ZN (n_14_33), .A (n_10_35), .B (n_4_38), .C1 (n_7_37), .C2 (n_13_34) );
AOI211_X1 g_16_32 (.ZN (n_16_32), .A (n_12_34), .B (n_6_37), .C1 (n_6_39), .C2 (n_11_35) );
AOI211_X1 g_15_34 (.ZN (n_15_34), .A (n_14_33), .B (n_8_36), .C1 (n_4_38), .C2 (n_9_36) );
AOI211_X1 g_13_35 (.ZN (n_13_35), .A (n_16_32), .B (n_10_35), .C1 (n_6_37), .C2 (n_7_37) );
AOI211_X1 g_11_36 (.ZN (n_11_36), .A (n_15_34), .B (n_12_34), .C1 (n_8_36), .C2 (n_6_39) );
AOI211_X1 g_9_37 (.ZN (n_9_37), .A (n_13_35), .B (n_14_33), .C1 (n_10_35), .C2 (n_4_38) );
AOI211_X1 g_7_38 (.ZN (n_7_38), .A (n_11_36), .B (n_16_32), .C1 (n_12_34), .C2 (n_6_37) );
AOI211_X1 g_5_39 (.ZN (n_5_39), .A (n_9_37), .B (n_15_34), .C1 (n_14_33), .C2 (n_8_36) );
AOI211_X1 g_3_40 (.ZN (n_3_40), .A (n_7_38), .B (n_13_35), .C1 (n_16_32), .C2 (n_10_35) );
AOI211_X1 g_2_42 (.ZN (n_2_42), .A (n_5_39), .B (n_11_36), .C1 (n_15_34), .C2 (n_12_34) );
AOI211_X1 g_1_44 (.ZN (n_1_44), .A (n_3_40), .B (n_9_37), .C1 (n_13_35), .C2 (n_14_33) );
AOI211_X1 g_3_43 (.ZN (n_3_43), .A (n_2_42), .B (n_7_38), .C1 (n_11_36), .C2 (n_16_32) );
AOI211_X1 g_4_41 (.ZN (n_4_41), .A (n_1_44), .B (n_5_39), .C1 (n_9_37), .C2 (n_15_34) );
AOI211_X1 g_6_40 (.ZN (n_6_40), .A (n_3_43), .B (n_3_40), .C1 (n_7_38), .C2 (n_13_35) );
AOI211_X1 g_4_39 (.ZN (n_4_39), .A (n_4_41), .B (n_2_42), .C1 (n_5_39), .C2 (n_11_36) );
AOI211_X1 g_3_41 (.ZN (n_3_41), .A (n_6_40), .B (n_1_44), .C1 (n_3_40), .C2 (n_9_37) );
AOI211_X1 g_5_42 (.ZN (n_5_42), .A (n_4_39), .B (n_3_43), .C1 (n_2_42), .C2 (n_7_38) );
AOI211_X1 g_7_41 (.ZN (n_7_41), .A (n_3_41), .B (n_4_41), .C1 (n_1_44), .C2 (n_5_39) );
AOI211_X1 g_8_39 (.ZN (n_8_39), .A (n_5_42), .B (n_6_40), .C1 (n_3_43), .C2 (n_3_40) );
AOI211_X1 g_6_38 (.ZN (n_6_38), .A (n_7_41), .B (n_4_39), .C1 (n_4_41), .C2 (n_2_42) );
AOI211_X1 g_8_37 (.ZN (n_8_37), .A (n_8_39), .B (n_3_41), .C1 (n_6_40), .C2 (n_1_44) );
AOI211_X1 g_10_38 (.ZN (n_10_38), .A (n_6_38), .B (n_5_42), .C1 (n_4_39), .C2 (n_3_43) );
AOI211_X1 g_12_37 (.ZN (n_12_37), .A (n_8_37), .B (n_7_41), .C1 (n_3_41), .C2 (n_4_41) );
AOI211_X1 g_14_36 (.ZN (n_14_36), .A (n_10_38), .B (n_8_39), .C1 (n_5_42), .C2 (n_6_40) );
AOI211_X1 g_16_35 (.ZN (n_16_35), .A (n_12_37), .B (n_6_38), .C1 (n_7_41), .C2 (n_4_39) );
AOI211_X1 g_18_34 (.ZN (n_18_34), .A (n_14_36), .B (n_8_37), .C1 (n_8_39), .C2 (n_3_41) );
AOI211_X1 g_17_36 (.ZN (n_17_36), .A (n_16_35), .B (n_10_38), .C1 (n_6_38), .C2 (n_5_42) );
AOI211_X1 g_16_34 (.ZN (n_16_34), .A (n_18_34), .B (n_12_37), .C1 (n_8_37), .C2 (n_7_41) );
AOI211_X1 g_18_33 (.ZN (n_18_33), .A (n_17_36), .B (n_14_36), .C1 (n_10_38), .C2 (n_8_39) );
AOI211_X1 g_17_35 (.ZN (n_17_35), .A (n_16_34), .B (n_16_35), .C1 (n_12_37), .C2 (n_6_38) );
AOI211_X1 g_15_36 (.ZN (n_15_36), .A (n_18_33), .B (n_18_34), .C1 (n_14_36), .C2 (n_8_37) );
AOI211_X1 g_13_37 (.ZN (n_13_37), .A (n_17_35), .B (n_17_36), .C1 (n_16_35), .C2 (n_10_38) );
AOI211_X1 g_14_35 (.ZN (n_14_35), .A (n_15_36), .B (n_16_34), .C1 (n_18_34), .C2 (n_12_37) );
AOI211_X1 g_12_36 (.ZN (n_12_36), .A (n_13_37), .B (n_18_33), .C1 (n_17_36), .C2 (n_14_36) );
AOI211_X1 g_10_37 (.ZN (n_10_37), .A (n_14_35), .B (n_17_35), .C1 (n_16_34), .C2 (n_16_35) );
AOI211_X1 g_8_38 (.ZN (n_8_38), .A (n_12_36), .B (n_15_36), .C1 (n_18_33), .C2 (n_18_34) );
AOI211_X1 g_7_40 (.ZN (n_7_40), .A (n_10_37), .B (n_13_37), .C1 (n_17_35), .C2 (n_17_36) );
AOI211_X1 g_5_41 (.ZN (n_5_41), .A (n_8_38), .B (n_14_35), .C1 (n_15_36), .C2 (n_16_34) );
AOI211_X1 g_4_43 (.ZN (n_4_43), .A (n_7_40), .B (n_12_36), .C1 (n_13_37), .C2 (n_18_33) );
AOI211_X1 g_3_45 (.ZN (n_3_45), .A (n_5_41), .B (n_10_37), .C1 (n_14_35), .C2 (n_17_35) );
AOI211_X1 g_5_46 (.ZN (n_5_46), .A (n_4_43), .B (n_8_38), .C1 (n_12_36), .C2 (n_15_36) );
AOI211_X1 g_3_47 (.ZN (n_3_47), .A (n_3_45), .B (n_7_40), .C1 (n_10_37), .C2 (n_13_37) );
AOI211_X1 g_1_48 (.ZN (n_1_48), .A (n_5_46), .B (n_5_41), .C1 (n_8_38), .C2 (n_14_35) );
AOI211_X1 g_2_46 (.ZN (n_2_46), .A (n_3_47), .B (n_4_43), .C1 (n_7_40), .C2 (n_12_36) );
AOI211_X1 g_4_45 (.ZN (n_4_45), .A (n_1_48), .B (n_3_45), .C1 (n_5_41), .C2 (n_10_37) );
AOI211_X1 g_6_44 (.ZN (n_6_44), .A (n_2_46), .B (n_5_46), .C1 (n_4_43), .C2 (n_8_38) );
AOI211_X1 g_7_42 (.ZN (n_7_42), .A (n_4_45), .B (n_3_47), .C1 (n_3_45), .C2 (n_7_40) );
AOI211_X1 g_5_43 (.ZN (n_5_43), .A (n_6_44), .B (n_1_48), .C1 (n_5_46), .C2 (n_5_41) );
AOI211_X1 g_3_44 (.ZN (n_3_44), .A (n_7_42), .B (n_2_46), .C1 (n_3_47), .C2 (n_4_43) );
AOI211_X1 g_4_42 (.ZN (n_4_42), .A (n_5_43), .B (n_4_45), .C1 (n_1_48), .C2 (n_3_45) );
AOI211_X1 g_5_40 (.ZN (n_5_40), .A (n_3_44), .B (n_6_44), .C1 (n_2_46), .C2 (n_5_46) );
AOI211_X1 g_7_39 (.ZN (n_7_39), .A (n_4_42), .B (n_7_42), .C1 (n_4_45), .C2 (n_3_47) );
AOI211_X1 g_6_41 (.ZN (n_6_41), .A (n_5_40), .B (n_5_43), .C1 (n_6_44), .C2 (n_1_48) );
AOI211_X1 g_8_40 (.ZN (n_8_40), .A (n_7_39), .B (n_3_44), .C1 (n_7_42), .C2 (n_2_46) );
AOI211_X1 g_9_38 (.ZN (n_9_38), .A (n_6_41), .B (n_4_42), .C1 (n_5_43), .C2 (n_4_45) );
AOI211_X1 g_11_37 (.ZN (n_11_37), .A (n_8_40), .B (n_5_40), .C1 (n_3_44), .C2 (n_6_44) );
AOI211_X1 g_13_36 (.ZN (n_13_36), .A (n_9_38), .B (n_7_39), .C1 (n_4_42), .C2 (n_7_42) );
AOI211_X1 g_15_35 (.ZN (n_15_35), .A (n_11_37), .B (n_6_41), .C1 (n_5_40), .C2 (n_5_43) );
AOI211_X1 g_17_34 (.ZN (n_17_34), .A (n_13_36), .B (n_8_40), .C1 (n_7_39), .C2 (n_3_44) );
AOI211_X1 g_19_33 (.ZN (n_19_33), .A (n_15_35), .B (n_9_38), .C1 (n_6_41), .C2 (n_4_42) );
AOI211_X1 g_21_32 (.ZN (n_21_32), .A (n_17_34), .B (n_11_37), .C1 (n_8_40), .C2 (n_5_40) );
AOI211_X1 g_20_34 (.ZN (n_20_34), .A (n_19_33), .B (n_13_36), .C1 (n_9_38), .C2 (n_7_39) );
AOI211_X1 g_22_33 (.ZN (n_22_33), .A (n_21_32), .B (n_15_35), .C1 (n_11_37), .C2 (n_6_41) );
AOI211_X1 g_24_32 (.ZN (n_24_32), .A (n_20_34), .B (n_17_34), .C1 (n_13_36), .C2 (n_8_40) );
AOI211_X1 g_26_31 (.ZN (n_26_31), .A (n_22_33), .B (n_19_33), .C1 (n_15_35), .C2 (n_9_38) );
AOI211_X1 g_28_30 (.ZN (n_28_30), .A (n_24_32), .B (n_21_32), .C1 (n_17_34), .C2 (n_11_37) );
AOI211_X1 g_30_29 (.ZN (n_30_29), .A (n_26_31), .B (n_20_34), .C1 (n_19_33), .C2 (n_13_36) );
AOI211_X1 g_32_28 (.ZN (n_32_28), .A (n_28_30), .B (n_22_33), .C1 (n_21_32), .C2 (n_15_35) );
AOI211_X1 g_34_27 (.ZN (n_34_27), .A (n_30_29), .B (n_24_32), .C1 (n_20_34), .C2 (n_17_34) );
AOI211_X1 g_36_26 (.ZN (n_36_26), .A (n_32_28), .B (n_26_31), .C1 (n_22_33), .C2 (n_19_33) );
AOI211_X1 g_38_25 (.ZN (n_38_25), .A (n_34_27), .B (n_28_30), .C1 (n_24_32), .C2 (n_21_32) );
AOI211_X1 g_40_24 (.ZN (n_40_24), .A (n_36_26), .B (n_30_29), .C1 (n_26_31), .C2 (n_20_34) );
AOI211_X1 g_42_23 (.ZN (n_42_23), .A (n_38_25), .B (n_32_28), .C1 (n_28_30), .C2 (n_22_33) );
AOI211_X1 g_44_22 (.ZN (n_44_22), .A (n_40_24), .B (n_34_27), .C1 (n_30_29), .C2 (n_24_32) );
AOI211_X1 g_46_21 (.ZN (n_46_21), .A (n_42_23), .B (n_36_26), .C1 (n_32_28), .C2 (n_26_31) );
AOI211_X1 g_48_20 (.ZN (n_48_20), .A (n_44_22), .B (n_38_25), .C1 (n_34_27), .C2 (n_28_30) );
AOI211_X1 g_50_19 (.ZN (n_50_19), .A (n_46_21), .B (n_40_24), .C1 (n_36_26), .C2 (n_30_29) );
AOI211_X1 g_49_21 (.ZN (n_49_21), .A (n_48_20), .B (n_42_23), .C1 (n_38_25), .C2 (n_32_28) );
AOI211_X1 g_51_20 (.ZN (n_51_20), .A (n_50_19), .B (n_44_22), .C1 (n_40_24), .C2 (n_34_27) );
AOI211_X1 g_53_19 (.ZN (n_53_19), .A (n_49_21), .B (n_46_21), .C1 (n_42_23), .C2 (n_36_26) );
AOI211_X1 g_55_20 (.ZN (n_55_20), .A (n_51_20), .B (n_48_20), .C1 (n_44_22), .C2 (n_38_25) );
AOI211_X1 g_56_18 (.ZN (n_56_18), .A (n_53_19), .B (n_50_19), .C1 (n_46_21), .C2 (n_40_24) );
AOI211_X1 g_58_17 (.ZN (n_58_17), .A (n_55_20), .B (n_49_21), .C1 (n_48_20), .C2 (n_42_23) );
AOI211_X1 g_60_16 (.ZN (n_60_16), .A (n_56_18), .B (n_51_20), .C1 (n_50_19), .C2 (n_44_22) );
AOI211_X1 g_62_15 (.ZN (n_62_15), .A (n_58_17), .B (n_53_19), .C1 (n_49_21), .C2 (n_46_21) );
AOI211_X1 g_64_14 (.ZN (n_64_14), .A (n_60_16), .B (n_55_20), .C1 (n_51_20), .C2 (n_48_20) );
AOI211_X1 g_66_13 (.ZN (n_66_13), .A (n_62_15), .B (n_56_18), .C1 (n_53_19), .C2 (n_50_19) );
AOI211_X1 g_68_12 (.ZN (n_68_12), .A (n_64_14), .B (n_58_17), .C1 (n_55_20), .C2 (n_49_21) );
AOI211_X1 g_70_13 (.ZN (n_70_13), .A (n_66_13), .B (n_60_16), .C1 (n_56_18), .C2 (n_51_20) );
AOI211_X1 g_68_14 (.ZN (n_68_14), .A (n_68_12), .B (n_62_15), .C1 (n_58_17), .C2 (n_53_19) );
AOI211_X1 g_70_15 (.ZN (n_70_15), .A (n_70_13), .B (n_64_14), .C1 (n_60_16), .C2 (n_55_20) );
AOI211_X1 g_69_17 (.ZN (n_69_17), .A (n_68_14), .B (n_66_13), .C1 (n_62_15), .C2 (n_56_18) );
AOI211_X1 g_68_15 (.ZN (n_68_15), .A (n_70_15), .B (n_68_12), .C1 (n_64_14), .C2 (n_58_17) );
AOI211_X1 g_67_13 (.ZN (n_67_13), .A (n_69_17), .B (n_70_13), .C1 (n_66_13), .C2 (n_60_16) );
AOI211_X1 g_65_14 (.ZN (n_65_14), .A (n_68_15), .B (n_68_14), .C1 (n_68_12), .C2 (n_62_15) );
AOI211_X1 g_63_15 (.ZN (n_63_15), .A (n_67_13), .B (n_70_15), .C1 (n_70_13), .C2 (n_64_14) );
AOI211_X1 g_61_16 (.ZN (n_61_16), .A (n_65_14), .B (n_69_17), .C1 (n_68_14), .C2 (n_66_13) );
AOI211_X1 g_59_17 (.ZN (n_59_17), .A (n_63_15), .B (n_68_15), .C1 (n_70_15), .C2 (n_68_12) );
AOI211_X1 g_57_18 (.ZN (n_57_18), .A (n_61_16), .B (n_67_13), .C1 (n_69_17), .C2 (n_70_13) );
AOI211_X1 g_55_17 (.ZN (n_55_17), .A (n_59_17), .B (n_65_14), .C1 (n_68_15), .C2 (n_68_14) );
AOI211_X1 g_53_18 (.ZN (n_53_18), .A (n_57_18), .B (n_63_15), .C1 (n_67_13), .C2 (n_70_15) );
AOI211_X1 g_51_19 (.ZN (n_51_19), .A (n_55_17), .B (n_61_16), .C1 (n_65_14), .C2 (n_69_17) );
AOI211_X1 g_49_20 (.ZN (n_49_20), .A (n_53_18), .B (n_59_17), .C1 (n_63_15), .C2 (n_68_15) );
AOI211_X1 g_47_21 (.ZN (n_47_21), .A (n_51_19), .B (n_57_18), .C1 (n_61_16), .C2 (n_67_13) );
AOI211_X1 g_45_22 (.ZN (n_45_22), .A (n_49_20), .B (n_55_17), .C1 (n_59_17), .C2 (n_65_14) );
AOI211_X1 g_43_23 (.ZN (n_43_23), .A (n_47_21), .B (n_53_18), .C1 (n_57_18), .C2 (n_63_15) );
AOI211_X1 g_41_24 (.ZN (n_41_24), .A (n_45_22), .B (n_51_19), .C1 (n_55_17), .C2 (n_61_16) );
AOI211_X1 g_39_25 (.ZN (n_39_25), .A (n_43_23), .B (n_49_20), .C1 (n_53_18), .C2 (n_59_17) );
AOI211_X1 g_37_26 (.ZN (n_37_26), .A (n_41_24), .B (n_47_21), .C1 (n_51_19), .C2 (n_57_18) );
AOI211_X1 g_35_27 (.ZN (n_35_27), .A (n_39_25), .B (n_45_22), .C1 (n_49_20), .C2 (n_55_17) );
AOI211_X1 g_33_28 (.ZN (n_33_28), .A (n_37_26), .B (n_43_23), .C1 (n_47_21), .C2 (n_53_18) );
AOI211_X1 g_31_29 (.ZN (n_31_29), .A (n_35_27), .B (n_41_24), .C1 (n_45_22), .C2 (n_51_19) );
AOI211_X1 g_29_30 (.ZN (n_29_30), .A (n_33_28), .B (n_39_25), .C1 (n_43_23), .C2 (n_49_20) );
AOI211_X1 g_27_31 (.ZN (n_27_31), .A (n_31_29), .B (n_37_26), .C1 (n_41_24), .C2 (n_47_21) );
AOI211_X1 g_25_32 (.ZN (n_25_32), .A (n_29_30), .B (n_35_27), .C1 (n_39_25), .C2 (n_45_22) );
AOI211_X1 g_23_33 (.ZN (n_23_33), .A (n_27_31), .B (n_33_28), .C1 (n_37_26), .C2 (n_43_23) );
AOI211_X1 g_21_34 (.ZN (n_21_34), .A (n_25_32), .B (n_31_29), .C1 (n_35_27), .C2 (n_41_24) );
AOI211_X1 g_19_35 (.ZN (n_19_35), .A (n_23_33), .B (n_29_30), .C1 (n_33_28), .C2 (n_39_25) );
AOI211_X1 g_18_37 (.ZN (n_18_37), .A (n_21_34), .B (n_27_31), .C1 (n_31_29), .C2 (n_37_26) );
AOI211_X1 g_16_36 (.ZN (n_16_36), .A (n_19_35), .B (n_25_32), .C1 (n_29_30), .C2 (n_35_27) );
AOI211_X1 g_18_35 (.ZN (n_18_35), .A (n_18_37), .B (n_23_33), .C1 (n_27_31), .C2 (n_33_28) );
AOI211_X1 g_20_36 (.ZN (n_20_36), .A (n_16_36), .B (n_21_34), .C1 (n_25_32), .C2 (n_31_29) );
AOI211_X1 g_22_35 (.ZN (n_22_35), .A (n_18_35), .B (n_19_35), .C1 (n_23_33), .C2 (n_29_30) );
AOI211_X1 g_21_33 (.ZN (n_21_33), .A (n_20_36), .B (n_18_37), .C1 (n_21_34), .C2 (n_27_31) );
AOI211_X1 g_23_32 (.ZN (n_23_32), .A (n_22_35), .B (n_16_36), .C1 (n_19_35), .C2 (n_25_32) );
AOI211_X1 g_25_31 (.ZN (n_25_31), .A (n_21_33), .B (n_18_35), .C1 (n_18_37), .C2 (n_23_33) );
AOI211_X1 g_27_30 (.ZN (n_27_30), .A (n_23_32), .B (n_20_36), .C1 (n_16_36), .C2 (n_21_34) );
AOI211_X1 g_26_32 (.ZN (n_26_32), .A (n_25_31), .B (n_22_35), .C1 (n_18_35), .C2 (n_19_35) );
AOI211_X1 g_28_31 (.ZN (n_28_31), .A (n_27_30), .B (n_21_33), .C1 (n_20_36), .C2 (n_18_37) );
AOI211_X1 g_30_30 (.ZN (n_30_30), .A (n_26_32), .B (n_23_32), .C1 (n_22_35), .C2 (n_16_36) );
AOI211_X1 g_32_29 (.ZN (n_32_29), .A (n_28_31), .B (n_25_31), .C1 (n_21_33), .C2 (n_18_35) );
AOI211_X1 g_34_28 (.ZN (n_34_28), .A (n_30_30), .B (n_27_30), .C1 (n_23_32), .C2 (n_20_36) );
AOI211_X1 g_36_27 (.ZN (n_36_27), .A (n_32_29), .B (n_26_32), .C1 (n_25_31), .C2 (n_22_35) );
AOI211_X1 g_35_29 (.ZN (n_35_29), .A (n_34_28), .B (n_28_31), .C1 (n_27_30), .C2 (n_21_33) );
AOI211_X1 g_37_28 (.ZN (n_37_28), .A (n_36_27), .B (n_30_30), .C1 (n_26_32), .C2 (n_23_32) );
AOI211_X1 g_39_27 (.ZN (n_39_27), .A (n_35_29), .B (n_32_29), .C1 (n_28_31), .C2 (n_25_31) );
AOI211_X1 g_41_26 (.ZN (n_41_26), .A (n_37_28), .B (n_34_28), .C1 (n_30_30), .C2 (n_27_30) );
AOI211_X1 g_43_25 (.ZN (n_43_25), .A (n_39_27), .B (n_36_27), .C1 (n_32_29), .C2 (n_26_32) );
AOI211_X1 g_45_24 (.ZN (n_45_24), .A (n_41_26), .B (n_35_29), .C1 (n_34_28), .C2 (n_28_31) );
AOI211_X1 g_46_22 (.ZN (n_46_22), .A (n_43_25), .B (n_37_28), .C1 (n_36_27), .C2 (n_30_30) );
AOI211_X1 g_48_21 (.ZN (n_48_21), .A (n_45_24), .B (n_39_27), .C1 (n_35_29), .C2 (n_32_29) );
AOI211_X1 g_50_20 (.ZN (n_50_20), .A (n_46_22), .B (n_41_26), .C1 (n_37_28), .C2 (n_34_28) );
AOI211_X1 g_49_22 (.ZN (n_49_22), .A (n_48_21), .B (n_43_25), .C1 (n_39_27), .C2 (n_36_27) );
AOI211_X1 g_47_23 (.ZN (n_47_23), .A (n_50_20), .B (n_45_24), .C1 (n_41_26), .C2 (n_35_29) );
AOI211_X1 g_46_25 (.ZN (n_46_25), .A (n_49_22), .B (n_46_22), .C1 (n_43_25), .C2 (n_37_28) );
AOI211_X1 g_45_23 (.ZN (n_45_23), .A (n_47_23), .B (n_48_21), .C1 (n_45_24), .C2 (n_39_27) );
AOI211_X1 g_47_22 (.ZN (n_47_22), .A (n_46_25), .B (n_50_20), .C1 (n_46_22), .C2 (n_41_26) );
AOI211_X1 g_46_24 (.ZN (n_46_24), .A (n_45_23), .B (n_49_22), .C1 (n_48_21), .C2 (n_43_25) );
AOI211_X1 g_48_23 (.ZN (n_48_23), .A (n_47_22), .B (n_47_23), .C1 (n_50_20), .C2 (n_45_24) );
AOI211_X1 g_50_22 (.ZN (n_50_22), .A (n_46_24), .B (n_46_25), .C1 (n_49_22), .C2 (n_46_22) );
AOI211_X1 g_52_21 (.ZN (n_52_21), .A (n_48_23), .B (n_45_23), .C1 (n_47_23), .C2 (n_48_21) );
AOI211_X1 g_54_20 (.ZN (n_54_20), .A (n_50_22), .B (n_47_22), .C1 (n_46_25), .C2 (n_50_20) );
AOI211_X1 g_56_19 (.ZN (n_56_19), .A (n_52_21), .B (n_46_24), .C1 (n_45_23), .C2 (n_49_22) );
AOI211_X1 g_57_21 (.ZN (n_57_21), .A (n_54_20), .B (n_48_23), .C1 (n_47_22), .C2 (n_47_23) );
AOI211_X1 g_58_19 (.ZN (n_58_19), .A (n_56_19), .B (n_50_22), .C1 (n_46_24), .C2 (n_46_25) );
AOI211_X1 g_60_18 (.ZN (n_60_18), .A (n_57_21), .B (n_52_21), .C1 (n_48_23), .C2 (n_45_23) );
AOI211_X1 g_62_17 (.ZN (n_62_17), .A (n_58_19), .B (n_54_20), .C1 (n_50_22), .C2 (n_47_22) );
AOI211_X1 g_64_16 (.ZN (n_64_16), .A (n_60_18), .B (n_56_19), .C1 (n_52_21), .C2 (n_46_24) );
AOI211_X1 g_66_15 (.ZN (n_66_15), .A (n_62_17), .B (n_57_21), .C1 (n_54_20), .C2 (n_48_23) );
AOI211_X1 g_65_17 (.ZN (n_65_17), .A (n_64_16), .B (n_58_19), .C1 (n_56_19), .C2 (n_50_22) );
AOI211_X1 g_67_16 (.ZN (n_67_16), .A (n_66_15), .B (n_60_18), .C1 (n_57_21), .C2 (n_52_21) );
AOI211_X1 g_69_15 (.ZN (n_69_15), .A (n_65_17), .B (n_62_17), .C1 (n_58_19), .C2 (n_54_20) );
AOI211_X1 g_67_14 (.ZN (n_67_14), .A (n_67_16), .B (n_64_16), .C1 (n_60_18), .C2 (n_56_19) );
AOI211_X1 g_65_15 (.ZN (n_65_15), .A (n_69_15), .B (n_66_15), .C1 (n_62_17), .C2 (n_57_21) );
AOI211_X1 g_63_16 (.ZN (n_63_16), .A (n_67_14), .B (n_65_17), .C1 (n_64_16), .C2 (n_58_19) );
AOI211_X1 g_61_17 (.ZN (n_61_17), .A (n_65_15), .B (n_67_16), .C1 (n_66_15), .C2 (n_60_18) );
AOI211_X1 g_59_18 (.ZN (n_59_18), .A (n_63_16), .B (n_69_15), .C1 (n_65_17), .C2 (n_62_17) );
AOI211_X1 g_57_19 (.ZN (n_57_19), .A (n_61_17), .B (n_67_14), .C1 (n_67_16), .C2 (n_64_16) );
AOI211_X1 g_59_20 (.ZN (n_59_20), .A (n_59_18), .B (n_65_15), .C1 (n_69_15), .C2 (n_66_15) );
AOI211_X1 g_61_19 (.ZN (n_61_19), .A (n_57_19), .B (n_63_16), .C1 (n_67_14), .C2 (n_65_17) );
AOI211_X1 g_60_17 (.ZN (n_60_17), .A (n_59_20), .B (n_61_17), .C1 (n_65_15), .C2 (n_67_16) );
AOI211_X1 g_59_19 (.ZN (n_59_19), .A (n_61_19), .B (n_59_18), .C1 (n_63_16), .C2 (n_69_15) );
AOI211_X1 g_61_18 (.ZN (n_61_18), .A (n_60_17), .B (n_57_19), .C1 (n_61_17), .C2 (n_67_14) );
AOI211_X1 g_63_17 (.ZN (n_63_17), .A (n_59_19), .B (n_59_20), .C1 (n_59_18), .C2 (n_65_15) );
AOI211_X1 g_65_16 (.ZN (n_65_16), .A (n_61_18), .B (n_61_19), .C1 (n_57_19), .C2 (n_63_16) );
AOI211_X1 g_67_15 (.ZN (n_67_15), .A (n_63_17), .B (n_60_17), .C1 (n_59_20), .C2 (n_61_17) );
AOI211_X1 g_69_14 (.ZN (n_69_14), .A (n_65_16), .B (n_59_19), .C1 (n_61_19), .C2 (n_59_18) );
AOI211_X1 g_68_16 (.ZN (n_68_16), .A (n_67_15), .B (n_61_18), .C1 (n_60_17), .C2 (n_57_19) );
AOI211_X1 g_66_17 (.ZN (n_66_17), .A (n_69_14), .B (n_63_17), .C1 (n_59_19), .C2 (n_59_20) );
AOI211_X1 g_64_18 (.ZN (n_64_18), .A (n_68_16), .B (n_65_16), .C1 (n_61_18), .C2 (n_61_19) );
AOI211_X1 g_62_19 (.ZN (n_62_19), .A (n_66_17), .B (n_67_15), .C1 (n_63_17), .C2 (n_60_17) );
AOI211_X1 g_60_20 (.ZN (n_60_20), .A (n_64_18), .B (n_69_14), .C1 (n_65_16), .C2 (n_59_19) );
AOI211_X1 g_58_21 (.ZN (n_58_21), .A (n_62_19), .B (n_68_16), .C1 (n_67_15), .C2 (n_61_18) );
AOI211_X1 g_56_20 (.ZN (n_56_20), .A (n_60_20), .B (n_66_17), .C1 (n_69_14), .C2 (n_63_17) );
AOI211_X1 g_54_19 (.ZN (n_54_19), .A (n_58_21), .B (n_64_18), .C1 (n_68_16), .C2 (n_65_16) );
AOI211_X1 g_52_20 (.ZN (n_52_20), .A (n_56_20), .B (n_62_19), .C1 (n_66_17), .C2 (n_67_15) );
AOI211_X1 g_50_21 (.ZN (n_50_21), .A (n_54_19), .B (n_60_20), .C1 (n_64_18), .C2 (n_69_14) );
AOI211_X1 g_48_22 (.ZN (n_48_22), .A (n_52_20), .B (n_58_21), .C1 (n_62_19), .C2 (n_68_16) );
AOI211_X1 g_46_23 (.ZN (n_46_23), .A (n_50_21), .B (n_56_20), .C1 (n_60_20), .C2 (n_66_17) );
AOI211_X1 g_44_24 (.ZN (n_44_24), .A (n_48_22), .B (n_54_19), .C1 (n_58_21), .C2 (n_64_18) );
AOI211_X1 g_42_25 (.ZN (n_42_25), .A (n_46_23), .B (n_52_20), .C1 (n_56_20), .C2 (n_62_19) );
AOI211_X1 g_40_26 (.ZN (n_40_26), .A (n_44_24), .B (n_50_21), .C1 (n_54_19), .C2 (n_60_20) );
AOI211_X1 g_38_27 (.ZN (n_38_27), .A (n_42_25), .B (n_48_22), .C1 (n_52_20), .C2 (n_58_21) );
AOI211_X1 g_36_28 (.ZN (n_36_28), .A (n_40_26), .B (n_46_23), .C1 (n_50_21), .C2 (n_56_20) );
AOI211_X1 g_34_29 (.ZN (n_34_29), .A (n_38_27), .B (n_44_24), .C1 (n_48_22), .C2 (n_54_19) );
AOI211_X1 g_32_30 (.ZN (n_32_30), .A (n_36_28), .B (n_42_25), .C1 (n_46_23), .C2 (n_52_20) );
AOI211_X1 g_30_31 (.ZN (n_30_31), .A (n_34_29), .B (n_40_26), .C1 (n_44_24), .C2 (n_50_21) );
AOI211_X1 g_28_32 (.ZN (n_28_32), .A (n_32_30), .B (n_38_27), .C1 (n_42_25), .C2 (n_48_22) );
AOI211_X1 g_26_33 (.ZN (n_26_33), .A (n_30_31), .B (n_36_28), .C1 (n_40_26), .C2 (n_46_23) );
AOI211_X1 g_24_34 (.ZN (n_24_34), .A (n_28_32), .B (n_34_29), .C1 (n_38_27), .C2 (n_44_24) );
AOI211_X1 g_23_36 (.ZN (n_23_36), .A (n_26_33), .B (n_32_30), .C1 (n_36_28), .C2 (n_42_25) );
AOI211_X1 g_22_34 (.ZN (n_22_34), .A (n_24_34), .B (n_30_31), .C1 (n_34_29), .C2 (n_40_26) );
AOI211_X1 g_24_33 (.ZN (n_24_33), .A (n_23_36), .B (n_28_32), .C1 (n_32_30), .C2 (n_38_27) );
AOI211_X1 g_23_35 (.ZN (n_23_35), .A (n_22_34), .B (n_26_33), .C1 (n_30_31), .C2 (n_36_28) );
AOI211_X1 g_25_34 (.ZN (n_25_34), .A (n_24_33), .B (n_24_34), .C1 (n_28_32), .C2 (n_34_29) );
AOI211_X1 g_27_33 (.ZN (n_27_33), .A (n_23_35), .B (n_23_36), .C1 (n_26_33), .C2 (n_32_30) );
AOI211_X1 g_29_32 (.ZN (n_29_32), .A (n_25_34), .B (n_22_34), .C1 (n_24_34), .C2 (n_30_31) );
AOI211_X1 g_31_31 (.ZN (n_31_31), .A (n_27_33), .B (n_24_33), .C1 (n_23_36), .C2 (n_28_32) );
AOI211_X1 g_33_30 (.ZN (n_33_30), .A (n_29_32), .B (n_23_35), .C1 (n_22_34), .C2 (n_26_33) );
AOI211_X1 g_32_32 (.ZN (n_32_32), .A (n_31_31), .B (n_25_34), .C1 (n_24_33), .C2 (n_24_34) );
AOI211_X1 g_31_30 (.ZN (n_31_30), .A (n_33_30), .B (n_27_33), .C1 (n_23_35), .C2 (n_23_36) );
AOI211_X1 g_33_29 (.ZN (n_33_29), .A (n_32_32), .B (n_29_32), .C1 (n_25_34), .C2 (n_22_34) );
AOI211_X1 g_35_28 (.ZN (n_35_28), .A (n_31_30), .B (n_31_31), .C1 (n_27_33), .C2 (n_24_33) );
AOI211_X1 g_37_27 (.ZN (n_37_27), .A (n_33_29), .B (n_33_30), .C1 (n_29_32), .C2 (n_23_35) );
AOI211_X1 g_39_26 (.ZN (n_39_26), .A (n_35_28), .B (n_32_32), .C1 (n_31_31), .C2 (n_25_34) );
AOI211_X1 g_41_25 (.ZN (n_41_25), .A (n_37_27), .B (n_31_30), .C1 (n_33_30), .C2 (n_27_33) );
AOI211_X1 g_43_24 (.ZN (n_43_24), .A (n_39_26), .B (n_33_29), .C1 (n_32_32), .C2 (n_29_32) );
AOI211_X1 g_44_26 (.ZN (n_44_26), .A (n_41_25), .B (n_35_28), .C1 (n_31_30), .C2 (n_31_31) );
AOI211_X1 g_42_27 (.ZN (n_42_27), .A (n_43_24), .B (n_37_27), .C1 (n_33_29), .C2 (n_33_30) );
AOI211_X1 g_40_28 (.ZN (n_40_28), .A (n_44_26), .B (n_39_26), .C1 (n_35_28), .C2 (n_32_32) );
AOI211_X1 g_38_29 (.ZN (n_38_29), .A (n_42_27), .B (n_41_25), .C1 (n_37_27), .C2 (n_31_30) );
AOI211_X1 g_36_30 (.ZN (n_36_30), .A (n_40_28), .B (n_43_24), .C1 (n_39_26), .C2 (n_33_29) );
AOI211_X1 g_34_31 (.ZN (n_34_31), .A (n_38_29), .B (n_44_26), .C1 (n_41_25), .C2 (n_35_28) );
AOI211_X1 g_33_33 (.ZN (n_33_33), .A (n_36_30), .B (n_42_27), .C1 (n_43_24), .C2 (n_37_27) );
AOI211_X1 g_32_31 (.ZN (n_32_31), .A (n_34_31), .B (n_40_28), .C1 (n_44_26), .C2 (n_39_26) );
AOI211_X1 g_34_30 (.ZN (n_34_30), .A (n_33_33), .B (n_38_29), .C1 (n_42_27), .C2 (n_41_25) );
AOI211_X1 g_36_29 (.ZN (n_36_29), .A (n_32_31), .B (n_36_30), .C1 (n_40_28), .C2 (n_43_24) );
AOI211_X1 g_38_28 (.ZN (n_38_28), .A (n_34_30), .B (n_34_31), .C1 (n_38_29), .C2 (n_44_26) );
AOI211_X1 g_40_27 (.ZN (n_40_27), .A (n_36_29), .B (n_33_33), .C1 (n_36_30), .C2 (n_42_27) );
AOI211_X1 g_42_26 (.ZN (n_42_26), .A (n_38_28), .B (n_32_31), .C1 (n_34_31), .C2 (n_40_28) );
AOI211_X1 g_44_25 (.ZN (n_44_25), .A (n_40_27), .B (n_34_30), .C1 (n_33_33), .C2 (n_38_29) );
AOI211_X1 g_43_27 (.ZN (n_43_27), .A (n_42_26), .B (n_36_29), .C1 (n_32_31), .C2 (n_36_30) );
AOI211_X1 g_45_26 (.ZN (n_45_26), .A (n_44_25), .B (n_38_28), .C1 (n_34_30), .C2 (n_34_31) );
AOI211_X1 g_47_25 (.ZN (n_47_25), .A (n_43_27), .B (n_40_27), .C1 (n_36_29), .C2 (n_33_33) );
AOI211_X1 g_49_24 (.ZN (n_49_24), .A (n_45_26), .B (n_42_26), .C1 (n_38_28), .C2 (n_32_31) );
AOI211_X1 g_51_23 (.ZN (n_51_23), .A (n_47_25), .B (n_44_25), .C1 (n_40_27), .C2 (n_34_30) );
AOI211_X1 g_53_22 (.ZN (n_53_22), .A (n_49_24), .B (n_43_27), .C1 (n_42_26), .C2 (n_36_29) );
AOI211_X1 g_51_21 (.ZN (n_51_21), .A (n_51_23), .B (n_45_26), .C1 (n_44_25), .C2 (n_38_28) );
AOI211_X1 g_53_20 (.ZN (n_53_20), .A (n_53_22), .B (n_47_25), .C1 (n_43_27), .C2 (n_40_27) );
AOI211_X1 g_55_19 (.ZN (n_55_19), .A (n_51_21), .B (n_49_24), .C1 (n_45_26), .C2 (n_42_26) );
AOI211_X1 g_54_21 (.ZN (n_54_21), .A (n_53_20), .B (n_51_23), .C1 (n_47_25), .C2 (n_44_25) );
AOI211_X1 g_52_22 (.ZN (n_52_22), .A (n_55_19), .B (n_53_22), .C1 (n_49_24), .C2 (n_43_27) );
AOI211_X1 g_50_23 (.ZN (n_50_23), .A (n_54_21), .B (n_51_21), .C1 (n_51_23), .C2 (n_45_26) );
AOI211_X1 g_48_24 (.ZN (n_48_24), .A (n_52_22), .B (n_53_20), .C1 (n_53_22), .C2 (n_47_25) );
AOI211_X1 g_47_26 (.ZN (n_47_26), .A (n_50_23), .B (n_55_19), .C1 (n_51_21), .C2 (n_49_24) );
AOI211_X1 g_45_25 (.ZN (n_45_25), .A (n_48_24), .B (n_54_21), .C1 (n_53_20), .C2 (n_51_23) );
AOI211_X1 g_47_24 (.ZN (n_47_24), .A (n_47_26), .B (n_52_22), .C1 (n_55_19), .C2 (n_53_22) );
AOI211_X1 g_49_23 (.ZN (n_49_23), .A (n_45_25), .B (n_50_23), .C1 (n_54_21), .C2 (n_51_21) );
AOI211_X1 g_51_22 (.ZN (n_51_22), .A (n_47_24), .B (n_48_24), .C1 (n_52_22), .C2 (n_53_20) );
AOI211_X1 g_53_21 (.ZN (n_53_21), .A (n_49_23), .B (n_47_26), .C1 (n_50_23), .C2 (n_55_19) );
AOI211_X1 g_55_22 (.ZN (n_55_22), .A (n_51_22), .B (n_45_25), .C1 (n_48_24), .C2 (n_54_21) );
AOI211_X1 g_53_23 (.ZN (n_53_23), .A (n_53_21), .B (n_47_24), .C1 (n_47_26), .C2 (n_52_22) );
AOI211_X1 g_51_24 (.ZN (n_51_24), .A (n_55_22), .B (n_49_23), .C1 (n_45_25), .C2 (n_50_23) );
AOI211_X1 g_49_25 (.ZN (n_49_25), .A (n_53_23), .B (n_51_22), .C1 (n_47_24), .C2 (n_48_24) );
AOI211_X1 g_48_27 (.ZN (n_48_27), .A (n_51_24), .B (n_53_21), .C1 (n_49_23), .C2 (n_47_26) );
AOI211_X1 g_46_26 (.ZN (n_46_26), .A (n_49_25), .B (n_55_22), .C1 (n_51_22), .C2 (n_45_25) );
AOI211_X1 g_48_25 (.ZN (n_48_25), .A (n_48_27), .B (n_53_23), .C1 (n_53_21), .C2 (n_47_24) );
AOI211_X1 g_50_24 (.ZN (n_50_24), .A (n_46_26), .B (n_51_24), .C1 (n_55_22), .C2 (n_49_23) );
AOI211_X1 g_52_23 (.ZN (n_52_23), .A (n_48_25), .B (n_49_25), .C1 (n_53_23), .C2 (n_51_22) );
AOI211_X1 g_54_22 (.ZN (n_54_22), .A (n_50_24), .B (n_48_27), .C1 (n_51_24), .C2 (n_53_21) );
AOI211_X1 g_56_21 (.ZN (n_56_21), .A (n_52_23), .B (n_46_26), .C1 (n_49_25), .C2 (n_55_22) );
AOI211_X1 g_58_20 (.ZN (n_58_20), .A (n_54_22), .B (n_48_25), .C1 (n_48_27), .C2 (n_53_23) );
AOI211_X1 g_60_19 (.ZN (n_60_19), .A (n_56_21), .B (n_50_24), .C1 (n_46_26), .C2 (n_51_24) );
AOI211_X1 g_62_18 (.ZN (n_62_18), .A (n_58_20), .B (n_52_23), .C1 (n_48_25), .C2 (n_49_25) );
AOI211_X1 g_64_17 (.ZN (n_64_17), .A (n_60_19), .B (n_54_22), .C1 (n_50_24), .C2 (n_48_27) );
AOI211_X1 g_66_16 (.ZN (n_66_16), .A (n_62_18), .B (n_56_21), .C1 (n_52_23), .C2 (n_46_26) );
AOI211_X1 g_67_18 (.ZN (n_67_18), .A (n_64_17), .B (n_58_20), .C1 (n_54_22), .C2 (n_48_25) );
AOI211_X1 g_65_19 (.ZN (n_65_19), .A (n_66_16), .B (n_60_19), .C1 (n_56_21), .C2 (n_50_24) );
AOI211_X1 g_63_18 (.ZN (n_63_18), .A (n_67_18), .B (n_62_18), .C1 (n_58_20), .C2 (n_52_23) );
AOI211_X1 g_62_20 (.ZN (n_62_20), .A (n_65_19), .B (n_64_17), .C1 (n_60_19), .C2 (n_54_22) );
AOI211_X1 g_64_19 (.ZN (n_64_19), .A (n_63_18), .B (n_66_16), .C1 (n_62_18), .C2 (n_56_21) );
AOI211_X1 g_66_18 (.ZN (n_66_18), .A (n_62_20), .B (n_67_18), .C1 (n_64_17), .C2 (n_58_20) );
AOI211_X1 g_68_17 (.ZN (n_68_17), .A (n_64_19), .B (n_65_19), .C1 (n_66_16), .C2 (n_60_19) );
AOI211_X1 g_70_16 (.ZN (n_70_16), .A (n_66_18), .B (n_63_18), .C1 (n_67_18), .C2 (n_62_18) );
AOI211_X1 g_72_15 (.ZN (n_72_15), .A (n_68_17), .B (n_62_20), .C1 (n_65_19), .C2 (n_64_17) );
AOI211_X1 g_74_14 (.ZN (n_74_14), .A (n_70_16), .B (n_64_19), .C1 (n_63_18), .C2 (n_66_16) );
AOI211_X1 g_76_13 (.ZN (n_76_13), .A (n_72_15), .B (n_66_18), .C1 (n_62_20), .C2 (n_67_18) );
AOI211_X1 g_78_12 (.ZN (n_78_12), .A (n_74_14), .B (n_68_17), .C1 (n_64_19), .C2 (n_65_19) );
AOI211_X1 g_77_14 (.ZN (n_77_14), .A (n_76_13), .B (n_70_16), .C1 (n_66_18), .C2 (n_63_18) );
AOI211_X1 g_75_15 (.ZN (n_75_15), .A (n_78_12), .B (n_72_15), .C1 (n_68_17), .C2 (n_62_20) );
AOI211_X1 g_73_16 (.ZN (n_73_16), .A (n_77_14), .B (n_74_14), .C1 (n_70_16), .C2 (n_64_19) );
AOI211_X1 g_71_15 (.ZN (n_71_15), .A (n_75_15), .B (n_76_13), .C1 (n_72_15), .C2 (n_66_18) );
AOI211_X1 g_69_16 (.ZN (n_69_16), .A (n_73_16), .B (n_78_12), .C1 (n_74_14), .C2 (n_68_17) );
AOI211_X1 g_67_17 (.ZN (n_67_17), .A (n_71_15), .B (n_77_14), .C1 (n_76_13), .C2 (n_70_16) );
AOI211_X1 g_65_18 (.ZN (n_65_18), .A (n_69_16), .B (n_75_15), .C1 (n_78_12), .C2 (n_72_15) );
AOI211_X1 g_63_19 (.ZN (n_63_19), .A (n_67_17), .B (n_73_16), .C1 (n_77_14), .C2 (n_74_14) );
AOI211_X1 g_61_20 (.ZN (n_61_20), .A (n_65_18), .B (n_71_15), .C1 (n_75_15), .C2 (n_76_13) );
AOI211_X1 g_59_21 (.ZN (n_59_21), .A (n_63_19), .B (n_69_16), .C1 (n_73_16), .C2 (n_78_12) );
AOI211_X1 g_57_20 (.ZN (n_57_20), .A (n_61_20), .B (n_67_17), .C1 (n_71_15), .C2 (n_77_14) );
AOI211_X1 g_55_21 (.ZN (n_55_21), .A (n_59_21), .B (n_65_18), .C1 (n_69_16), .C2 (n_75_15) );
AOI211_X1 g_57_22 (.ZN (n_57_22), .A (n_57_20), .B (n_63_19), .C1 (n_67_17), .C2 (n_73_16) );
AOI211_X1 g_55_23 (.ZN (n_55_23), .A (n_55_21), .B (n_61_20), .C1 (n_65_18), .C2 (n_71_15) );
AOI211_X1 g_53_24 (.ZN (n_53_24), .A (n_57_22), .B (n_59_21), .C1 (n_63_19), .C2 (n_69_16) );
AOI211_X1 g_51_25 (.ZN (n_51_25), .A (n_55_23), .B (n_57_20), .C1 (n_61_20), .C2 (n_67_17) );
AOI211_X1 g_49_26 (.ZN (n_49_26), .A (n_53_24), .B (n_55_21), .C1 (n_59_21), .C2 (n_65_18) );
AOI211_X1 g_47_27 (.ZN (n_47_27), .A (n_51_25), .B (n_57_22), .C1 (n_57_20), .C2 (n_63_19) );
AOI211_X1 g_45_28 (.ZN (n_45_28), .A (n_49_26), .B (n_55_23), .C1 (n_55_21), .C2 (n_61_20) );
AOI211_X1 g_43_29 (.ZN (n_43_29), .A (n_47_27), .B (n_53_24), .C1 (n_57_22), .C2 (n_59_21) );
AOI211_X1 g_44_27 (.ZN (n_44_27), .A (n_45_28), .B (n_51_25), .C1 (n_55_23), .C2 (n_57_20) );
AOI211_X1 g_46_28 (.ZN (n_46_28), .A (n_43_29), .B (n_49_26), .C1 (n_53_24), .C2 (n_55_21) );
AOI211_X1 g_44_29 (.ZN (n_44_29), .A (n_44_27), .B (n_47_27), .C1 (n_51_25), .C2 (n_57_22) );
AOI211_X1 g_45_27 (.ZN (n_45_27), .A (n_46_28), .B (n_45_28), .C1 (n_49_26), .C2 (n_55_23) );
AOI211_X1 g_43_26 (.ZN (n_43_26), .A (n_44_29), .B (n_43_29), .C1 (n_47_27), .C2 (n_53_24) );
AOI211_X1 g_42_28 (.ZN (n_42_28), .A (n_45_27), .B (n_44_27), .C1 (n_45_28), .C2 (n_51_25) );
AOI211_X1 g_40_29 (.ZN (n_40_29), .A (n_43_26), .B (n_46_28), .C1 (n_43_29), .C2 (n_49_26) );
AOI211_X1 g_41_27 (.ZN (n_41_27), .A (n_42_28), .B (n_44_29), .C1 (n_44_27), .C2 (n_47_27) );
AOI211_X1 g_39_28 (.ZN (n_39_28), .A (n_40_29), .B (n_45_27), .C1 (n_46_28), .C2 (n_45_28) );
AOI211_X1 g_37_29 (.ZN (n_37_29), .A (n_41_27), .B (n_43_26), .C1 (n_44_29), .C2 (n_43_29) );
AOI211_X1 g_35_30 (.ZN (n_35_30), .A (n_39_28), .B (n_42_28), .C1 (n_45_27), .C2 (n_44_27) );
AOI211_X1 g_33_31 (.ZN (n_33_31), .A (n_37_29), .B (n_40_29), .C1 (n_43_26), .C2 (n_46_28) );
AOI211_X1 g_31_32 (.ZN (n_31_32), .A (n_35_30), .B (n_41_27), .C1 (n_42_28), .C2 (n_44_29) );
AOI211_X1 g_29_31 (.ZN (n_29_31), .A (n_33_31), .B (n_39_28), .C1 (n_40_29), .C2 (n_45_27) );
AOI211_X1 g_27_32 (.ZN (n_27_32), .A (n_31_32), .B (n_37_29), .C1 (n_41_27), .C2 (n_43_26) );
AOI211_X1 g_25_33 (.ZN (n_25_33), .A (n_29_31), .B (n_35_30), .C1 (n_39_28), .C2 (n_42_28) );
AOI211_X1 g_23_34 (.ZN (n_23_34), .A (n_27_32), .B (n_33_31), .C1 (n_37_29), .C2 (n_40_29) );
AOI211_X1 g_21_35 (.ZN (n_21_35), .A (n_25_33), .B (n_31_32), .C1 (n_35_30), .C2 (n_41_27) );
AOI211_X1 g_19_36 (.ZN (n_19_36), .A (n_23_34), .B (n_29_31), .C1 (n_33_31), .C2 (n_39_28) );
AOI211_X1 g_17_37 (.ZN (n_17_37), .A (n_21_35), .B (n_27_32), .C1 (n_31_32), .C2 (n_37_29) );
AOI211_X1 g_15_38 (.ZN (n_15_38), .A (n_19_36), .B (n_25_33), .C1 (n_29_31), .C2 (n_35_30) );
AOI211_X1 g_13_39 (.ZN (n_13_39), .A (n_17_37), .B (n_23_34), .C1 (n_27_32), .C2 (n_33_31) );
AOI211_X1 g_14_37 (.ZN (n_14_37), .A (n_15_38), .B (n_21_35), .C1 (n_25_33), .C2 (n_31_32) );
AOI211_X1 g_12_38 (.ZN (n_12_38), .A (n_13_39), .B (n_19_36), .C1 (n_23_34), .C2 (n_29_31) );
AOI211_X1 g_10_39 (.ZN (n_10_39), .A (n_14_37), .B (n_17_37), .C1 (n_21_35), .C2 (n_27_32) );
AOI211_X1 g_9_41 (.ZN (n_9_41), .A (n_12_38), .B (n_15_38), .C1 (n_19_36), .C2 (n_25_33) );
AOI211_X1 g_11_40 (.ZN (n_11_40), .A (n_10_39), .B (n_13_39), .C1 (n_17_37), .C2 (n_23_34) );
AOI211_X1 g_9_39 (.ZN (n_9_39), .A (n_9_41), .B (n_14_37), .C1 (n_15_38), .C2 (n_21_35) );
AOI211_X1 g_11_38 (.ZN (n_11_38), .A (n_11_40), .B (n_12_38), .C1 (n_13_39), .C2 (n_19_36) );
AOI211_X1 g_10_40 (.ZN (n_10_40), .A (n_9_39), .B (n_10_39), .C1 (n_14_37), .C2 (n_17_37) );
AOI211_X1 g_12_39 (.ZN (n_12_39), .A (n_11_38), .B (n_9_41), .C1 (n_12_38), .C2 (n_15_38) );
AOI211_X1 g_14_38 (.ZN (n_14_38), .A (n_10_40), .B (n_11_40), .C1 (n_10_39), .C2 (n_13_39) );
AOI211_X1 g_16_37 (.ZN (n_16_37), .A (n_12_39), .B (n_9_39), .C1 (n_9_41), .C2 (n_14_37) );
AOI211_X1 g_18_36 (.ZN (n_18_36), .A (n_14_38), .B (n_11_38), .C1 (n_11_40), .C2 (n_12_38) );
AOI211_X1 g_20_35 (.ZN (n_20_35), .A (n_16_37), .B (n_10_40), .C1 (n_9_39), .C2 (n_10_39) );
AOI211_X1 g_21_37 (.ZN (n_21_37), .A (n_18_36), .B (n_12_39), .C1 (n_11_38), .C2 (n_9_41) );
AOI211_X1 g_19_38 (.ZN (n_19_38), .A (n_20_35), .B (n_14_38), .C1 (n_10_40), .C2 (n_11_40) );
AOI211_X1 g_17_39 (.ZN (n_17_39), .A (n_21_37), .B (n_16_37), .C1 (n_12_39), .C2 (n_9_39) );
AOI211_X1 g_15_40 (.ZN (n_15_40), .A (n_19_38), .B (n_18_36), .C1 (n_14_38), .C2 (n_11_38) );
AOI211_X1 g_16_38 (.ZN (n_16_38), .A (n_17_39), .B (n_20_35), .C1 (n_16_37), .C2 (n_10_40) );
AOI211_X1 g_14_39 (.ZN (n_14_39), .A (n_15_40), .B (n_21_37), .C1 (n_18_36), .C2 (n_12_39) );
AOI211_X1 g_15_37 (.ZN (n_15_37), .A (n_16_38), .B (n_19_38), .C1 (n_20_35), .C2 (n_14_38) );
AOI211_X1 g_13_38 (.ZN (n_13_38), .A (n_14_39), .B (n_17_39), .C1 (n_21_37), .C2 (n_16_37) );
AOI211_X1 g_11_39 (.ZN (n_11_39), .A (n_15_37), .B (n_15_40), .C1 (n_19_38), .C2 (n_18_36) );
AOI211_X1 g_9_40 (.ZN (n_9_40), .A (n_13_38), .B (n_16_38), .C1 (n_17_39), .C2 (n_20_35) );
AOI211_X1 g_8_42 (.ZN (n_8_42), .A (n_11_39), .B (n_14_39), .C1 (n_15_40), .C2 (n_21_37) );
AOI211_X1 g_6_43 (.ZN (n_6_43), .A (n_9_40), .B (n_15_37), .C1 (n_16_38), .C2 (n_19_38) );
AOI211_X1 g_5_45 (.ZN (n_5_45), .A (n_8_42), .B (n_13_38), .C1 (n_14_39), .C2 (n_17_39) );
AOI211_X1 g_4_47 (.ZN (n_4_47), .A (n_6_43), .B (n_11_39), .C1 (n_15_37), .C2 (n_15_40) );
AOI211_X1 g_3_49 (.ZN (n_3_49), .A (n_5_45), .B (n_9_40), .C1 (n_13_38), .C2 (n_16_38) );
AOI211_X1 g_5_50 (.ZN (n_5_50), .A (n_4_47), .B (n_8_42), .C1 (n_11_39), .C2 (n_14_39) );
AOI211_X1 g_3_51 (.ZN (n_3_51), .A (n_3_49), .B (n_6_43), .C1 (n_9_40), .C2 (n_15_37) );
AOI211_X1 g_1_52 (.ZN (n_1_52), .A (n_5_50), .B (n_5_45), .C1 (n_8_42), .C2 (n_13_38) );
AOI211_X1 g_2_50 (.ZN (n_2_50), .A (n_3_51), .B (n_4_47), .C1 (n_6_43), .C2 (n_11_39) );
AOI211_X1 g_4_49 (.ZN (n_4_49), .A (n_1_52), .B (n_3_49), .C1 (n_5_45), .C2 (n_9_40) );
AOI211_X1 g_6_48 (.ZN (n_6_48), .A (n_2_50), .B (n_5_50), .C1 (n_4_47), .C2 (n_8_42) );
AOI211_X1 g_7_46 (.ZN (n_7_46), .A (n_4_49), .B (n_3_51), .C1 (n_3_49), .C2 (n_6_43) );
AOI211_X1 g_5_47 (.ZN (n_5_47), .A (n_6_48), .B (n_1_52), .C1 (n_5_50), .C2 (n_5_45) );
AOI211_X1 g_3_48 (.ZN (n_3_48), .A (n_7_46), .B (n_2_50), .C1 (n_3_51), .C2 (n_4_47) );
AOI211_X1 g_4_46 (.ZN (n_4_46), .A (n_5_47), .B (n_4_49), .C1 (n_1_52), .C2 (n_3_49) );
AOI211_X1 g_6_45 (.ZN (n_6_45), .A (n_3_48), .B (n_6_48), .C1 (n_2_50), .C2 (n_5_50) );
AOI211_X1 g_8_44 (.ZN (n_8_44), .A (n_4_46), .B (n_7_46), .C1 (n_4_49), .C2 (n_3_51) );
AOI211_X1 g_9_42 (.ZN (n_9_42), .A (n_6_45), .B (n_5_47), .C1 (n_6_48), .C2 (n_1_52) );
AOI211_X1 g_11_41 (.ZN (n_11_41), .A (n_8_44), .B (n_3_48), .C1 (n_7_46), .C2 (n_2_50) );
AOI211_X1 g_13_40 (.ZN (n_13_40), .A (n_9_42), .B (n_4_46), .C1 (n_5_47), .C2 (n_4_49) );
AOI211_X1 g_15_39 (.ZN (n_15_39), .A (n_11_41), .B (n_6_45), .C1 (n_3_48), .C2 (n_6_48) );
AOI211_X1 g_17_38 (.ZN (n_17_38), .A (n_13_40), .B (n_8_44), .C1 (n_4_46), .C2 (n_7_46) );
AOI211_X1 g_19_37 (.ZN (n_19_37), .A (n_15_39), .B (n_9_42), .C1 (n_6_45), .C2 (n_5_47) );
AOI211_X1 g_21_36 (.ZN (n_21_36), .A (n_17_38), .B (n_11_41), .C1 (n_8_44), .C2 (n_3_48) );
AOI211_X1 g_20_38 (.ZN (n_20_38), .A (n_19_37), .B (n_13_40), .C1 (n_9_42), .C2 (n_4_46) );
AOI211_X1 g_22_37 (.ZN (n_22_37), .A (n_21_36), .B (n_15_39), .C1 (n_11_41), .C2 (n_6_45) );
AOI211_X1 g_24_36 (.ZN (n_24_36), .A (n_20_38), .B (n_17_38), .C1 (n_13_40), .C2 (n_8_44) );
AOI211_X1 g_26_35 (.ZN (n_26_35), .A (n_22_37), .B (n_19_37), .C1 (n_15_39), .C2 (n_9_42) );
AOI211_X1 g_28_34 (.ZN (n_28_34), .A (n_24_36), .B (n_21_36), .C1 (n_17_38), .C2 (n_11_41) );
AOI211_X1 g_30_33 (.ZN (n_30_33), .A (n_26_35), .B (n_20_38), .C1 (n_19_37), .C2 (n_13_40) );
AOI211_X1 g_32_34 (.ZN (n_32_34), .A (n_28_34), .B (n_22_37), .C1 (n_21_36), .C2 (n_15_39) );
AOI211_X1 g_33_32 (.ZN (n_33_32), .A (n_30_33), .B (n_24_36), .C1 (n_20_38), .C2 (n_17_38) );
AOI211_X1 g_35_31 (.ZN (n_35_31), .A (n_32_34), .B (n_26_35), .C1 (n_22_37), .C2 (n_19_37) );
AOI211_X1 g_37_30 (.ZN (n_37_30), .A (n_33_32), .B (n_28_34), .C1 (n_24_36), .C2 (n_21_36) );
AOI211_X1 g_39_29 (.ZN (n_39_29), .A (n_35_31), .B (n_30_33), .C1 (n_26_35), .C2 (n_20_38) );
AOI211_X1 g_41_28 (.ZN (n_41_28), .A (n_37_30), .B (n_32_34), .C1 (n_28_34), .C2 (n_22_37) );
AOI211_X1 g_40_30 (.ZN (n_40_30), .A (n_39_29), .B (n_33_32), .C1 (n_30_33), .C2 (n_24_36) );
AOI211_X1 g_42_29 (.ZN (n_42_29), .A (n_41_28), .B (n_35_31), .C1 (n_32_34), .C2 (n_26_35) );
AOI211_X1 g_44_28 (.ZN (n_44_28), .A (n_40_30), .B (n_37_30), .C1 (n_33_32), .C2 (n_28_34) );
AOI211_X1 g_46_27 (.ZN (n_46_27), .A (n_42_29), .B (n_39_29), .C1 (n_35_31), .C2 (n_30_33) );
AOI211_X1 g_48_26 (.ZN (n_48_26), .A (n_44_28), .B (n_41_28), .C1 (n_37_30), .C2 (n_32_34) );
AOI211_X1 g_50_25 (.ZN (n_50_25), .A (n_46_27), .B (n_40_30), .C1 (n_39_29), .C2 (n_33_32) );
AOI211_X1 g_52_24 (.ZN (n_52_24), .A (n_48_26), .B (n_42_29), .C1 (n_41_28), .C2 (n_35_31) );
AOI211_X1 g_54_23 (.ZN (n_54_23), .A (n_50_25), .B (n_44_28), .C1 (n_40_30), .C2 (n_37_30) );
AOI211_X1 g_56_22 (.ZN (n_56_22), .A (n_52_24), .B (n_46_27), .C1 (n_42_29), .C2 (n_39_29) );
AOI211_X1 g_55_24 (.ZN (n_55_24), .A (n_54_23), .B (n_48_26), .C1 (n_44_28), .C2 (n_41_28) );
AOI211_X1 g_57_23 (.ZN (n_57_23), .A (n_56_22), .B (n_50_25), .C1 (n_46_27), .C2 (n_40_30) );
AOI211_X1 g_59_22 (.ZN (n_59_22), .A (n_55_24), .B (n_52_24), .C1 (n_48_26), .C2 (n_42_29) );
AOI211_X1 g_61_21 (.ZN (n_61_21), .A (n_57_23), .B (n_54_23), .C1 (n_50_25), .C2 (n_44_28) );
AOI211_X1 g_63_20 (.ZN (n_63_20), .A (n_59_22), .B (n_56_22), .C1 (n_52_24), .C2 (n_46_27) );
AOI211_X1 g_62_22 (.ZN (n_62_22), .A (n_61_21), .B (n_55_24), .C1 (n_54_23), .C2 (n_48_26) );
AOI211_X1 g_60_21 (.ZN (n_60_21), .A (n_63_20), .B (n_57_23), .C1 (n_56_22), .C2 (n_50_25) );
AOI211_X1 g_58_22 (.ZN (n_58_22), .A (n_62_22), .B (n_59_22), .C1 (n_55_24), .C2 (n_52_24) );
AOI211_X1 g_56_23 (.ZN (n_56_23), .A (n_60_21), .B (n_61_21), .C1 (n_57_23), .C2 (n_54_23) );
AOI211_X1 g_54_24 (.ZN (n_54_24), .A (n_58_22), .B (n_63_20), .C1 (n_59_22), .C2 (n_56_22) );
AOI211_X1 g_52_25 (.ZN (n_52_25), .A (n_56_23), .B (n_62_22), .C1 (n_61_21), .C2 (n_55_24) );
AOI211_X1 g_50_26 (.ZN (n_50_26), .A (n_54_24), .B (n_60_21), .C1 (n_63_20), .C2 (n_57_23) );
AOI211_X1 g_49_28 (.ZN (n_49_28), .A (n_52_25), .B (n_58_22), .C1 (n_62_22), .C2 (n_59_22) );
AOI211_X1 g_51_27 (.ZN (n_51_27), .A (n_50_26), .B (n_56_23), .C1 (n_60_21), .C2 (n_61_21) );
AOI211_X1 g_53_26 (.ZN (n_53_26), .A (n_49_28), .B (n_54_24), .C1 (n_58_22), .C2 (n_63_20) );
AOI211_X1 g_55_25 (.ZN (n_55_25), .A (n_51_27), .B (n_52_25), .C1 (n_56_23), .C2 (n_62_22) );
AOI211_X1 g_57_24 (.ZN (n_57_24), .A (n_53_26), .B (n_50_26), .C1 (n_54_24), .C2 (n_60_21) );
AOI211_X1 g_59_23 (.ZN (n_59_23), .A (n_55_25), .B (n_49_28), .C1 (n_52_25), .C2 (n_58_22) );
AOI211_X1 g_61_22 (.ZN (n_61_22), .A (n_57_24), .B (n_51_27), .C1 (n_50_26), .C2 (n_56_23) );
AOI211_X1 g_63_21 (.ZN (n_63_21), .A (n_59_23), .B (n_53_26), .C1 (n_49_28), .C2 (n_54_24) );
AOI211_X1 g_65_20 (.ZN (n_65_20), .A (n_61_22), .B (n_55_25), .C1 (n_51_27), .C2 (n_52_25) );
AOI211_X1 g_67_19 (.ZN (n_67_19), .A (n_63_21), .B (n_57_24), .C1 (n_53_26), .C2 (n_50_26) );
AOI211_X1 g_69_18 (.ZN (n_69_18), .A (n_65_20), .B (n_59_23), .C1 (n_55_25), .C2 (n_49_28) );
AOI211_X1 g_71_17 (.ZN (n_71_17), .A (n_67_19), .B (n_61_22), .C1 (n_57_24), .C2 (n_51_27) );
AOI211_X1 g_70_19 (.ZN (n_70_19), .A (n_69_18), .B (n_63_21), .C1 (n_59_23), .C2 (n_53_26) );
AOI211_X1 g_68_18 (.ZN (n_68_18), .A (n_71_17), .B (n_65_20), .C1 (n_61_22), .C2 (n_55_25) );
AOI211_X1 g_70_17 (.ZN (n_70_17), .A (n_70_19), .B (n_67_19), .C1 (n_63_21), .C2 (n_57_24) );
AOI211_X1 g_72_18 (.ZN (n_72_18), .A (n_68_18), .B (n_69_18), .C1 (n_65_20), .C2 (n_59_23) );
AOI211_X1 g_74_17 (.ZN (n_74_17), .A (n_70_17), .B (n_71_17), .C1 (n_67_19), .C2 (n_61_22) );
AOI211_X1 g_76_16 (.ZN (n_76_16), .A (n_72_18), .B (n_70_19), .C1 (n_69_18), .C2 (n_63_21) );
AOI211_X1 g_78_15 (.ZN (n_78_15), .A (n_74_17), .B (n_68_18), .C1 (n_71_17), .C2 (n_65_20) );
AOI211_X1 g_77_13 (.ZN (n_77_13), .A (n_76_16), .B (n_70_17), .C1 (n_70_19), .C2 (n_67_19) );
AOI211_X1 g_79_12 (.ZN (n_79_12), .A (n_78_15), .B (n_72_18), .C1 (n_68_18), .C2 (n_69_18) );
AOI211_X1 g_81_11 (.ZN (n_81_11), .A (n_77_13), .B (n_74_17), .C1 (n_70_17), .C2 (n_71_17) );
AOI211_X1 g_82_13 (.ZN (n_82_13), .A (n_79_12), .B (n_76_16), .C1 (n_72_18), .C2 (n_70_19) );
AOI211_X1 g_80_14 (.ZN (n_80_14), .A (n_81_11), .B (n_78_15), .C1 (n_74_17), .C2 (n_68_18) );
AOI211_X1 g_82_15 (.ZN (n_82_15), .A (n_82_13), .B (n_77_13), .C1 (n_76_16), .C2 (n_70_17) );
AOI211_X1 g_81_13 (.ZN (n_81_13), .A (n_80_14), .B (n_79_12), .C1 (n_78_15), .C2 (n_72_18) );
AOI211_X1 g_83_12 (.ZN (n_83_12), .A (n_82_15), .B (n_81_11), .C1 (n_77_13), .C2 (n_74_17) );
AOI211_X1 g_85_11 (.ZN (n_85_11), .A (n_81_13), .B (n_82_13), .C1 (n_79_12), .C2 (n_76_16) );
AOI211_X1 g_86_13 (.ZN (n_86_13), .A (n_83_12), .B (n_80_14), .C1 (n_81_11), .C2 (n_78_15) );
AOI211_X1 g_84_14 (.ZN (n_84_14), .A (n_85_11), .B (n_82_15), .C1 (n_82_13), .C2 (n_77_13) );
AOI211_X1 g_86_15 (.ZN (n_86_15), .A (n_86_13), .B (n_81_13), .C1 (n_80_14), .C2 (n_79_12) );
AOI211_X1 g_85_13 (.ZN (n_85_13), .A (n_84_14), .B (n_83_12), .C1 (n_82_15), .C2 (n_81_11) );
AOI211_X1 g_87_12 (.ZN (n_87_12), .A (n_86_15), .B (n_85_11), .C1 (n_81_13), .C2 (n_82_13) );
AOI211_X1 g_89_11 (.ZN (n_89_11), .A (n_85_13), .B (n_86_13), .C1 (n_83_12), .C2 (n_80_14) );
AOI211_X1 g_90_13 (.ZN (n_90_13), .A (n_87_12), .B (n_84_14), .C1 (n_85_11), .C2 (n_82_15) );
AOI211_X1 g_88_14 (.ZN (n_88_14), .A (n_89_11), .B (n_86_15), .C1 (n_86_13), .C2 (n_81_13) );
AOI211_X1 g_90_15 (.ZN (n_90_15), .A (n_90_13), .B (n_85_13), .C1 (n_84_14), .C2 (n_83_12) );
AOI211_X1 g_89_13 (.ZN (n_89_13), .A (n_88_14), .B (n_87_12), .C1 (n_86_15), .C2 (n_85_11) );
AOI211_X1 g_91_12 (.ZN (n_91_12), .A (n_90_15), .B (n_89_11), .C1 (n_85_13), .C2 (n_86_13) );
AOI211_X1 g_93_11 (.ZN (n_93_11), .A (n_89_13), .B (n_90_13), .C1 (n_87_12), .C2 (n_84_14) );
AOI211_X1 g_94_13 (.ZN (n_94_13), .A (n_91_12), .B (n_88_14), .C1 (n_89_11), .C2 (n_86_15) );
AOI211_X1 g_92_14 (.ZN (n_92_14), .A (n_93_11), .B (n_90_15), .C1 (n_90_13), .C2 (n_85_13) );
AOI211_X1 g_94_15 (.ZN (n_94_15), .A (n_94_13), .B (n_89_13), .C1 (n_88_14), .C2 (n_87_12) );
AOI211_X1 g_93_13 (.ZN (n_93_13), .A (n_92_14), .B (n_91_12), .C1 (n_90_15), .C2 (n_89_11) );
AOI211_X1 g_95_12 (.ZN (n_95_12), .A (n_94_15), .B (n_93_11), .C1 (n_89_13), .C2 (n_90_13) );
AOI211_X1 g_97_11 (.ZN (n_97_11), .A (n_93_13), .B (n_94_13), .C1 (n_91_12), .C2 (n_88_14) );
AOI211_X1 g_98_13 (.ZN (n_98_13), .A (n_95_12), .B (n_92_14), .C1 (n_93_11), .C2 (n_90_15) );
AOI211_X1 g_96_14 (.ZN (n_96_14), .A (n_97_11), .B (n_94_15), .C1 (n_94_13), .C2 (n_89_13) );
AOI211_X1 g_98_15 (.ZN (n_98_15), .A (n_98_13), .B (n_93_13), .C1 (n_92_14), .C2 (n_91_12) );
AOI211_X1 g_97_13 (.ZN (n_97_13), .A (n_96_14), .B (n_95_12), .C1 (n_94_15), .C2 (n_93_11) );
AOI211_X1 g_99_12 (.ZN (n_99_12), .A (n_98_15), .B (n_97_11), .C1 (n_93_13), .C2 (n_94_13) );
AOI211_X1 g_101_11 (.ZN (n_101_11), .A (n_97_13), .B (n_98_13), .C1 (n_95_12), .C2 (n_92_14) );
AOI211_X1 g_102_13 (.ZN (n_102_13), .A (n_99_12), .B (n_96_14), .C1 (n_97_11), .C2 (n_94_15) );
AOI211_X1 g_100_14 (.ZN (n_100_14), .A (n_101_11), .B (n_98_15), .C1 (n_98_13), .C2 (n_93_13) );
AOI211_X1 g_102_15 (.ZN (n_102_15), .A (n_102_13), .B (n_97_13), .C1 (n_96_14), .C2 (n_95_12) );
AOI211_X1 g_101_13 (.ZN (n_101_13), .A (n_100_14), .B (n_99_12), .C1 (n_98_15), .C2 (n_97_11) );
AOI211_X1 g_103_12 (.ZN (n_103_12), .A (n_102_15), .B (n_101_11), .C1 (n_97_13), .C2 (n_98_13) );
AOI211_X1 g_105_11 (.ZN (n_105_11), .A (n_101_13), .B (n_102_13), .C1 (n_99_12), .C2 (n_96_14) );
AOI211_X1 g_106_13 (.ZN (n_106_13), .A (n_103_12), .B (n_100_14), .C1 (n_101_11), .C2 (n_98_15) );
AOI211_X1 g_104_14 (.ZN (n_104_14), .A (n_105_11), .B (n_102_15), .C1 (n_102_13), .C2 (n_97_13) );
AOI211_X1 g_106_15 (.ZN (n_106_15), .A (n_106_13), .B (n_101_13), .C1 (n_100_14), .C2 (n_99_12) );
AOI211_X1 g_105_13 (.ZN (n_105_13), .A (n_104_14), .B (n_103_12), .C1 (n_102_15), .C2 (n_101_11) );
AOI211_X1 g_107_12 (.ZN (n_107_12), .A (n_106_15), .B (n_105_11), .C1 (n_101_13), .C2 (n_102_13) );
AOI211_X1 g_109_11 (.ZN (n_109_11), .A (n_105_13), .B (n_106_13), .C1 (n_103_12), .C2 (n_100_14) );
AOI211_X1 g_110_13 (.ZN (n_110_13), .A (n_107_12), .B (n_104_14), .C1 (n_105_11), .C2 (n_102_15) );
AOI211_X1 g_108_14 (.ZN (n_108_14), .A (n_109_11), .B (n_106_15), .C1 (n_106_13), .C2 (n_101_13) );
AOI211_X1 g_110_15 (.ZN (n_110_15), .A (n_110_13), .B (n_105_13), .C1 (n_104_14), .C2 (n_103_12) );
AOI211_X1 g_109_13 (.ZN (n_109_13), .A (n_108_14), .B (n_107_12), .C1 (n_106_15), .C2 (n_105_11) );
AOI211_X1 g_111_12 (.ZN (n_111_12), .A (n_110_15), .B (n_109_11), .C1 (n_105_13), .C2 (n_106_13) );
AOI211_X1 g_113_11 (.ZN (n_113_11), .A (n_109_13), .B (n_110_13), .C1 (n_107_12), .C2 (n_104_14) );
AOI211_X1 g_114_13 (.ZN (n_114_13), .A (n_111_12), .B (n_108_14), .C1 (n_109_11), .C2 (n_106_15) );
AOI211_X1 g_112_14 (.ZN (n_112_14), .A (n_113_11), .B (n_110_15), .C1 (n_110_13), .C2 (n_105_13) );
AOI211_X1 g_114_15 (.ZN (n_114_15), .A (n_114_13), .B (n_109_13), .C1 (n_108_14), .C2 (n_107_12) );
AOI211_X1 g_113_13 (.ZN (n_113_13), .A (n_112_14), .B (n_111_12), .C1 (n_110_15), .C2 (n_109_11) );
AOI211_X1 g_115_12 (.ZN (n_115_12), .A (n_114_15), .B (n_113_11), .C1 (n_109_13), .C2 (n_110_13) );
AOI211_X1 g_117_11 (.ZN (n_117_11), .A (n_113_13), .B (n_114_13), .C1 (n_111_12), .C2 (n_108_14) );
AOI211_X1 g_118_13 (.ZN (n_118_13), .A (n_115_12), .B (n_112_14), .C1 (n_113_11), .C2 (n_110_15) );
AOI211_X1 g_116_14 (.ZN (n_116_14), .A (n_117_11), .B (n_114_15), .C1 (n_114_13), .C2 (n_109_13) );
AOI211_X1 g_118_15 (.ZN (n_118_15), .A (n_118_13), .B (n_113_13), .C1 (n_112_14), .C2 (n_111_12) );
AOI211_X1 g_117_13 (.ZN (n_117_13), .A (n_116_14), .B (n_115_12), .C1 (n_114_15), .C2 (n_113_11) );
AOI211_X1 g_119_12 (.ZN (n_119_12), .A (n_118_15), .B (n_117_11), .C1 (n_113_13), .C2 (n_114_13) );
AOI211_X1 g_121_11 (.ZN (n_121_11), .A (n_117_13), .B (n_118_13), .C1 (n_115_12), .C2 (n_112_14) );
AOI211_X1 g_122_13 (.ZN (n_122_13), .A (n_119_12), .B (n_116_14), .C1 (n_117_11), .C2 (n_114_15) );
AOI211_X1 g_120_14 (.ZN (n_120_14), .A (n_121_11), .B (n_118_15), .C1 (n_118_13), .C2 (n_113_13) );
AOI211_X1 g_122_15 (.ZN (n_122_15), .A (n_122_13), .B (n_117_13), .C1 (n_116_14), .C2 (n_115_12) );
AOI211_X1 g_121_13 (.ZN (n_121_13), .A (n_120_14), .B (n_119_12), .C1 (n_118_15), .C2 (n_117_11) );
AOI211_X1 g_123_12 (.ZN (n_123_12), .A (n_122_15), .B (n_121_11), .C1 (n_117_13), .C2 (n_118_13) );
AOI211_X1 g_125_11 (.ZN (n_125_11), .A (n_121_13), .B (n_122_13), .C1 (n_119_12), .C2 (n_116_14) );
AOI211_X1 g_126_13 (.ZN (n_126_13), .A (n_123_12), .B (n_120_14), .C1 (n_121_11), .C2 (n_118_15) );
AOI211_X1 g_124_14 (.ZN (n_124_14), .A (n_125_11), .B (n_122_15), .C1 (n_122_13), .C2 (n_117_13) );
AOI211_X1 g_126_15 (.ZN (n_126_15), .A (n_126_13), .B (n_121_13), .C1 (n_120_14), .C2 (n_119_12) );
AOI211_X1 g_125_13 (.ZN (n_125_13), .A (n_124_14), .B (n_123_12), .C1 (n_122_15), .C2 (n_121_11) );
AOI211_X1 g_127_12 (.ZN (n_127_12), .A (n_126_15), .B (n_125_11), .C1 (n_121_13), .C2 (n_122_13) );
AOI211_X1 g_129_11 (.ZN (n_129_11), .A (n_125_13), .B (n_126_13), .C1 (n_123_12), .C2 (n_120_14) );
AOI211_X1 g_130_13 (.ZN (n_130_13), .A (n_127_12), .B (n_124_14), .C1 (n_125_11), .C2 (n_122_15) );
AOI211_X1 g_128_14 (.ZN (n_128_14), .A (n_129_11), .B (n_126_15), .C1 (n_126_13), .C2 (n_121_13) );
AOI211_X1 g_130_15 (.ZN (n_130_15), .A (n_130_13), .B (n_125_13), .C1 (n_124_14), .C2 (n_123_12) );
AOI211_X1 g_132_14 (.ZN (n_132_14), .A (n_128_14), .B (n_127_12), .C1 (n_126_15), .C2 (n_125_11) );
AOI211_X1 g_131_12 (.ZN (n_131_12), .A (n_130_15), .B (n_129_11), .C1 (n_125_13), .C2 (n_126_13) );
AOI211_X1 g_129_13 (.ZN (n_129_13), .A (n_132_14), .B (n_130_13), .C1 (n_127_12), .C2 (n_124_14) );
AOI211_X1 g_127_14 (.ZN (n_127_14), .A (n_131_12), .B (n_128_14), .C1 (n_129_11), .C2 (n_126_15) );
AOI211_X1 g_126_12 (.ZN (n_126_12), .A (n_129_13), .B (n_130_15), .C1 (n_130_13), .C2 (n_125_13) );
AOI211_X1 g_124_13 (.ZN (n_124_13), .A (n_127_14), .B (n_132_14), .C1 (n_128_14), .C2 (n_127_12) );
AOI211_X1 g_122_14 (.ZN (n_122_14), .A (n_126_12), .B (n_131_12), .C1 (n_130_15), .C2 (n_129_11) );
AOI211_X1 g_120_13 (.ZN (n_120_13), .A (n_124_13), .B (n_129_13), .C1 (n_132_14), .C2 (n_130_13) );
AOI211_X1 g_118_12 (.ZN (n_118_12), .A (n_122_14), .B (n_127_14), .C1 (n_131_12), .C2 (n_128_14) );
AOI211_X1 g_117_14 (.ZN (n_117_14), .A (n_120_13), .B (n_126_12), .C1 (n_129_13), .C2 (n_130_15) );
AOI211_X1 g_119_15 (.ZN (n_119_15), .A (n_118_12), .B (n_124_13), .C1 (n_127_14), .C2 (n_132_14) );
AOI211_X1 g_121_16 (.ZN (n_121_16), .A (n_117_14), .B (n_122_14), .C1 (n_126_12), .C2 (n_131_12) );
AOI211_X1 g_123_15 (.ZN (n_123_15), .A (n_119_15), .B (n_120_13), .C1 (n_124_13), .C2 (n_129_13) );
AOI211_X1 g_125_14 (.ZN (n_125_14), .A (n_121_16), .B (n_118_12), .C1 (n_122_14), .C2 (n_127_14) );
AOI211_X1 g_124_16 (.ZN (n_124_16), .A (n_123_15), .B (n_117_14), .C1 (n_120_13), .C2 (n_126_12) );
AOI211_X1 g_123_14 (.ZN (n_123_14), .A (n_125_14), .B (n_119_15), .C1 (n_118_12), .C2 (n_124_13) );
AOI211_X1 g_125_15 (.ZN (n_125_15), .A (n_124_16), .B (n_121_16), .C1 (n_117_14), .C2 (n_122_14) );
AOI211_X1 g_123_16 (.ZN (n_123_16), .A (n_123_14), .B (n_123_15), .C1 (n_119_15), .C2 (n_120_13) );
AOI211_X1 g_121_15 (.ZN (n_121_15), .A (n_125_15), .B (n_125_14), .C1 (n_121_16), .C2 (n_118_12) );
AOI211_X1 g_119_14 (.ZN (n_119_14), .A (n_123_16), .B (n_124_16), .C1 (n_123_15), .C2 (n_117_14) );
AOI211_X1 g_120_16 (.ZN (n_120_16), .A (n_121_15), .B (n_123_14), .C1 (n_125_14), .C2 (n_119_15) );
AOI211_X1 g_122_17 (.ZN (n_122_17), .A (n_119_14), .B (n_125_15), .C1 (n_124_16), .C2 (n_121_16) );
AOI211_X1 g_120_18 (.ZN (n_120_18), .A (n_120_16), .B (n_123_16), .C1 (n_123_14), .C2 (n_123_15) );
AOI211_X1 g_119_16 (.ZN (n_119_16), .A (n_122_17), .B (n_121_15), .C1 (n_125_15), .C2 (n_125_14) );
AOI211_X1 g_118_14 (.ZN (n_118_14), .A (n_120_18), .B (n_119_14), .C1 (n_123_16), .C2 (n_124_16) );
AOI211_X1 g_116_13 (.ZN (n_116_13), .A (n_119_16), .B (n_120_16), .C1 (n_121_15), .C2 (n_123_14) );
AOI211_X1 g_114_12 (.ZN (n_114_12), .A (n_118_14), .B (n_122_17), .C1 (n_119_14), .C2 (n_125_15) );
AOI211_X1 g_112_13 (.ZN (n_112_13), .A (n_116_13), .B (n_120_18), .C1 (n_120_16), .C2 (n_123_16) );
AOI211_X1 g_114_14 (.ZN (n_114_14), .A (n_114_12), .B (n_119_16), .C1 (n_122_17), .C2 (n_121_15) );
AOI211_X1 g_116_15 (.ZN (n_116_15), .A (n_112_13), .B (n_118_14), .C1 (n_120_18), .C2 (n_119_14) );
AOI211_X1 g_117_17 (.ZN (n_117_17), .A (n_114_14), .B (n_116_13), .C1 (n_119_16), .C2 (n_120_16) );
AOI211_X1 g_115_16 (.ZN (n_115_16), .A (n_116_15), .B (n_114_12), .C1 (n_118_14), .C2 (n_122_17) );
AOI211_X1 g_117_15 (.ZN (n_117_15), .A (n_117_17), .B (n_112_13), .C1 (n_116_13), .C2 (n_120_18) );
AOI211_X1 g_115_14 (.ZN (n_115_14), .A (n_115_16), .B (n_114_14), .C1 (n_114_12), .C2 (n_119_16) );
AOI211_X1 g_113_15 (.ZN (n_113_15), .A (n_117_15), .B (n_116_15), .C1 (n_112_13), .C2 (n_118_14) );
AOI211_X1 g_111_14 (.ZN (n_111_14), .A (n_115_14), .B (n_117_17), .C1 (n_114_14), .C2 (n_116_13) );
AOI211_X1 g_112_16 (.ZN (n_112_16), .A (n_113_15), .B (n_115_16), .C1 (n_116_15), .C2 (n_114_12) );
AOI211_X1 g_113_14 (.ZN (n_113_14), .A (n_111_14), .B (n_117_15), .C1 (n_117_17), .C2 (n_112_13) );
AOI211_X1 g_111_15 (.ZN (n_111_15), .A (n_112_16), .B (n_115_14), .C1 (n_115_16), .C2 (n_114_14) );
AOI211_X1 g_113_16 (.ZN (n_113_16), .A (n_113_14), .B (n_113_15), .C1 (n_117_15), .C2 (n_116_15) );
AOI211_X1 g_115_15 (.ZN (n_115_15), .A (n_111_15), .B (n_111_14), .C1 (n_115_14), .C2 (n_117_17) );
AOI211_X1 g_117_16 (.ZN (n_117_16), .A (n_113_16), .B (n_112_16), .C1 (n_113_15), .C2 (n_115_16) );
AOI211_X1 g_115_17 (.ZN (n_115_17), .A (n_115_15), .B (n_113_14), .C1 (n_111_14), .C2 (n_117_15) );
AOI211_X1 g_113_18 (.ZN (n_113_18), .A (n_117_16), .B (n_111_15), .C1 (n_112_16), .C2 (n_115_14) );
AOI211_X1 g_114_16 (.ZN (n_114_16), .A (n_115_17), .B (n_113_16), .C1 (n_113_14), .C2 (n_113_15) );
AOI211_X1 g_112_15 (.ZN (n_112_15), .A (n_113_18), .B (n_115_15), .C1 (n_111_15), .C2 (n_111_14) );
AOI211_X1 g_110_14 (.ZN (n_110_14), .A (n_114_16), .B (n_117_16), .C1 (n_113_16), .C2 (n_112_16) );
AOI211_X1 g_108_13 (.ZN (n_108_13), .A (n_112_15), .B (n_115_17), .C1 (n_115_15), .C2 (n_113_14) );
AOI211_X1 g_106_12 (.ZN (n_106_12), .A (n_110_14), .B (n_113_18), .C1 (n_117_16), .C2 (n_111_15) );
AOI211_X1 g_105_14 (.ZN (n_105_14), .A (n_108_13), .B (n_114_16), .C1 (n_115_17), .C2 (n_113_16) );
AOI211_X1 g_107_15 (.ZN (n_107_15), .A (n_106_12), .B (n_112_15), .C1 (n_113_18), .C2 (n_115_15) );
AOI211_X1 g_109_16 (.ZN (n_109_16), .A (n_105_14), .B (n_110_14), .C1 (n_114_16), .C2 (n_117_16) );
AOI211_X1 g_111_17 (.ZN (n_111_17), .A (n_107_15), .B (n_108_13), .C1 (n_112_15), .C2 (n_115_17) );
AOI211_X1 g_109_18 (.ZN (n_109_18), .A (n_109_16), .B (n_106_12), .C1 (n_110_14), .C2 (n_113_18) );
AOI211_X1 g_110_16 (.ZN (n_110_16), .A (n_111_17), .B (n_105_14), .C1 (n_108_13), .C2 (n_114_16) );
AOI211_X1 g_108_15 (.ZN (n_108_15), .A (n_109_18), .B (n_107_15), .C1 (n_106_12), .C2 (n_112_15) );
AOI211_X1 g_106_14 (.ZN (n_106_14), .A (n_110_16), .B (n_109_16), .C1 (n_105_14), .C2 (n_110_14) );
AOI211_X1 g_104_13 (.ZN (n_104_13), .A (n_108_15), .B (n_111_17), .C1 (n_107_15), .C2 (n_108_13) );
AOI211_X1 g_102_12 (.ZN (n_102_12), .A (n_106_14), .B (n_109_18), .C1 (n_109_16), .C2 (n_106_12) );
AOI211_X1 g_100_13 (.ZN (n_100_13), .A (n_104_13), .B (n_110_16), .C1 (n_111_17), .C2 (n_105_14) );
AOI211_X1 g_102_14 (.ZN (n_102_14), .A (n_102_12), .B (n_108_15), .C1 (n_109_18), .C2 (n_107_15) );
AOI211_X1 g_104_15 (.ZN (n_104_15), .A (n_100_13), .B (n_106_14), .C1 (n_110_16), .C2 (n_109_16) );
AOI211_X1 g_106_16 (.ZN (n_106_16), .A (n_102_14), .B (n_104_13), .C1 (n_108_15), .C2 (n_111_17) );
AOI211_X1 g_107_14 (.ZN (n_107_14), .A (n_104_15), .B (n_102_12), .C1 (n_106_14), .C2 (n_109_18) );
AOI211_X1 g_108_16 (.ZN (n_108_16), .A (n_106_16), .B (n_100_13), .C1 (n_104_13), .C2 (n_110_16) );
AOI211_X1 g_110_17 (.ZN (n_110_17), .A (n_107_14), .B (n_102_14), .C1 (n_102_12), .C2 (n_108_15) );
AOI211_X1 g_109_15 (.ZN (n_109_15), .A (n_108_16), .B (n_104_15), .C1 (n_100_13), .C2 (n_106_14) );
AOI211_X1 g_108_17 (.ZN (n_108_17), .A (n_110_17), .B (n_106_16), .C1 (n_102_14), .C2 (n_104_13) );
AOI211_X1 g_107_19 (.ZN (n_107_19), .A (n_109_15), .B (n_107_14), .C1 (n_104_15), .C2 (n_102_12) );
AOI211_X1 g_106_17 (.ZN (n_106_17), .A (n_108_17), .B (n_108_16), .C1 (n_106_16), .C2 (n_100_13) );
AOI211_X1 g_105_15 (.ZN (n_105_15), .A (n_107_19), .B (n_110_17), .C1 (n_107_14), .C2 (n_102_14) );
AOI211_X1 g_103_14 (.ZN (n_103_14), .A (n_106_17), .B (n_109_15), .C1 (n_108_16), .C2 (n_104_15) );
AOI211_X1 g_104_16 (.ZN (n_104_16), .A (n_105_15), .B (n_108_17), .C1 (n_110_17), .C2 (n_106_16) );
AOI211_X1 g_105_18 (.ZN (n_105_18), .A (n_103_14), .B (n_107_19), .C1 (n_109_15), .C2 (n_107_14) );
AOI211_X1 g_107_17 (.ZN (n_107_17), .A (n_104_16), .B (n_106_17), .C1 (n_108_17), .C2 (n_108_16) );
AOI211_X1 g_105_16 (.ZN (n_105_16), .A (n_105_18), .B (n_105_15), .C1 (n_107_19), .C2 (n_110_17) );
AOI211_X1 g_103_15 (.ZN (n_103_15), .A (n_107_17), .B (n_103_14), .C1 (n_106_17), .C2 (n_109_15) );
AOI211_X1 g_101_14 (.ZN (n_101_14), .A (n_105_16), .B (n_104_16), .C1 (n_105_15), .C2 (n_108_17) );
AOI211_X1 g_99_15 (.ZN (n_99_15), .A (n_103_15), .B (n_105_18), .C1 (n_103_14), .C2 (n_107_19) );
AOI211_X1 g_101_16 (.ZN (n_101_16), .A (n_101_14), .B (n_107_17), .C1 (n_104_16), .C2 (n_106_17) );
AOI211_X1 g_103_17 (.ZN (n_103_17), .A (n_99_15), .B (n_105_16), .C1 (n_105_18), .C2 (n_105_15) );
AOI211_X1 g_101_18 (.ZN (n_101_18), .A (n_101_16), .B (n_103_15), .C1 (n_107_17), .C2 (n_103_14) );
AOI211_X1 g_102_16 (.ZN (n_102_16), .A (n_103_17), .B (n_101_14), .C1 (n_105_16), .C2 (n_104_16) );
AOI211_X1 g_100_15 (.ZN (n_100_15), .A (n_101_18), .B (n_99_15), .C1 (n_103_15), .C2 (n_105_18) );
AOI211_X1 g_98_14 (.ZN (n_98_14), .A (n_102_16), .B (n_101_16), .C1 (n_101_14), .C2 (n_107_17) );
AOI211_X1 g_96_13 (.ZN (n_96_13), .A (n_100_15), .B (n_103_17), .C1 (n_99_15), .C2 (n_105_16) );
AOI211_X1 g_94_12 (.ZN (n_94_12), .A (n_98_14), .B (n_101_18), .C1 (n_101_16), .C2 (n_103_15) );
AOI211_X1 g_93_14 (.ZN (n_93_14), .A (n_96_13), .B (n_102_16), .C1 (n_103_17), .C2 (n_101_14) );
AOI211_X1 g_95_15 (.ZN (n_95_15), .A (n_94_12), .B (n_100_15), .C1 (n_101_18), .C2 (n_99_15) );
AOI211_X1 g_97_16 (.ZN (n_97_16), .A (n_93_14), .B (n_98_14), .C1 (n_102_16), .C2 (n_101_16) );
AOI211_X1 g_99_17 (.ZN (n_99_17), .A (n_95_15), .B (n_96_13), .C1 (n_100_15), .C2 (n_103_17) );
AOI211_X1 g_97_18 (.ZN (n_97_18), .A (n_97_16), .B (n_94_12), .C1 (n_98_14), .C2 (n_101_18) );
AOI211_X1 g_96_16 (.ZN (n_96_16), .A (n_99_17), .B (n_93_14), .C1 (n_96_13), .C2 (n_102_16) );
AOI211_X1 g_95_14 (.ZN (n_95_14), .A (n_97_18), .B (n_95_15), .C1 (n_94_12), .C2 (n_100_15) );
AOI211_X1 g_97_15 (.ZN (n_97_15), .A (n_96_16), .B (n_97_16), .C1 (n_93_14), .C2 (n_98_14) );
AOI211_X1 g_99_14 (.ZN (n_99_14), .A (n_95_14), .B (n_99_17), .C1 (n_95_15), .C2 (n_96_13) );
AOI211_X1 g_100_16 (.ZN (n_100_16), .A (n_97_15), .B (n_97_18), .C1 (n_97_16), .C2 (n_94_12) );
AOI211_X1 g_98_17 (.ZN (n_98_17), .A (n_99_14), .B (n_96_16), .C1 (n_99_17), .C2 (n_93_14) );
AOI211_X1 g_99_19 (.ZN (n_99_19), .A (n_100_16), .B (n_95_14), .C1 (n_97_18), .C2 (n_95_15) );
AOI211_X1 g_100_17 (.ZN (n_100_17), .A (n_98_17), .B (n_97_15), .C1 (n_96_16), .C2 (n_97_16) );
AOI211_X1 g_101_15 (.ZN (n_101_15), .A (n_99_19), .B (n_99_14), .C1 (n_95_14), .C2 (n_99_17) );
AOI211_X1 g_99_16 (.ZN (n_99_16), .A (n_100_17), .B (n_100_16), .C1 (n_97_15), .C2 (n_97_18) );
AOI211_X1 g_98_18 (.ZN (n_98_18), .A (n_101_15), .B (n_98_17), .C1 (n_99_14), .C2 (n_96_16) );
AOI211_X1 g_96_17 (.ZN (n_96_17), .A (n_99_16), .B (n_99_19), .C1 (n_100_16), .C2 (n_95_14) );
AOI211_X1 g_98_16 (.ZN (n_98_16), .A (n_98_18), .B (n_100_17), .C1 (n_98_17), .C2 (n_97_15) );
AOI211_X1 g_96_15 (.ZN (n_96_15), .A (n_96_17), .B (n_101_15), .C1 (n_99_19), .C2 (n_99_14) );
AOI211_X1 g_94_14 (.ZN (n_94_14), .A (n_98_16), .B (n_99_16), .C1 (n_100_17), .C2 (n_100_16) );
AOI211_X1 g_92_13 (.ZN (n_92_13), .A (n_96_15), .B (n_98_18), .C1 (n_101_15), .C2 (n_98_17) );
AOI211_X1 g_90_12 (.ZN (n_90_12), .A (n_94_14), .B (n_96_17), .C1 (n_99_16), .C2 (n_99_19) );
AOI211_X1 g_88_13 (.ZN (n_88_13), .A (n_92_13), .B (n_98_16), .C1 (n_98_18), .C2 (n_100_17) );
AOI211_X1 g_90_14 (.ZN (n_90_14), .A (n_90_12), .B (n_96_15), .C1 (n_96_17), .C2 (n_101_15) );
AOI211_X1 g_92_15 (.ZN (n_92_15), .A (n_88_13), .B (n_94_14), .C1 (n_98_16), .C2 (n_99_16) );
AOI211_X1 g_94_16 (.ZN (n_94_16), .A (n_90_14), .B (n_92_13), .C1 (n_96_15), .C2 (n_98_18) );
AOI211_X1 g_95_18 (.ZN (n_95_18), .A (n_92_15), .B (n_90_12), .C1 (n_94_14), .C2 (n_96_17) );
AOI211_X1 g_97_17 (.ZN (n_97_17), .A (n_94_16), .B (n_88_13), .C1 (n_92_13), .C2 (n_98_16) );
AOI211_X1 g_95_16 (.ZN (n_95_16), .A (n_95_18), .B (n_90_14), .C1 (n_90_12), .C2 (n_96_15) );
AOI211_X1 g_93_15 (.ZN (n_93_15), .A (n_97_17), .B (n_92_15), .C1 (n_88_13), .C2 (n_94_14) );
AOI211_X1 g_91_14 (.ZN (n_91_14), .A (n_95_16), .B (n_94_16), .C1 (n_90_14), .C2 (n_92_13) );
AOI211_X1 g_92_16 (.ZN (n_92_16), .A (n_93_15), .B (n_95_18), .C1 (n_92_15), .C2 (n_90_12) );
AOI211_X1 g_94_17 (.ZN (n_94_17), .A (n_91_14), .B (n_97_17), .C1 (n_94_16), .C2 (n_88_13) );
AOI211_X1 g_96_18 (.ZN (n_96_18), .A (n_92_16), .B (n_95_16), .C1 (n_95_18), .C2 (n_90_14) );
AOI211_X1 g_97_20 (.ZN (n_97_20), .A (n_94_17), .B (n_93_15), .C1 (n_97_17), .C2 (n_92_15) );
AOI211_X1 g_95_19 (.ZN (n_95_19), .A (n_96_18), .B (n_91_14), .C1 (n_95_16), .C2 (n_94_16) );
AOI211_X1 g_93_18 (.ZN (n_93_18), .A (n_97_20), .B (n_92_16), .C1 (n_93_15), .C2 (n_95_18) );
AOI211_X1 g_95_17 (.ZN (n_95_17), .A (n_95_19), .B (n_94_17), .C1 (n_91_14), .C2 (n_97_17) );
AOI211_X1 g_93_16 (.ZN (n_93_16), .A (n_93_18), .B (n_96_18), .C1 (n_92_16), .C2 (n_95_16) );
AOI211_X1 g_91_15 (.ZN (n_91_15), .A (n_95_17), .B (n_97_20), .C1 (n_94_17), .C2 (n_93_15) );
AOI211_X1 g_89_14 (.ZN (n_89_14), .A (n_93_16), .B (n_95_19), .C1 (n_96_18), .C2 (n_91_14) );
AOI211_X1 g_87_15 (.ZN (n_87_15), .A (n_91_15), .B (n_93_18), .C1 (n_97_20), .C2 (n_92_16) );
AOI211_X1 g_89_16 (.ZN (n_89_16), .A (n_89_14), .B (n_95_17), .C1 (n_95_19), .C2 (n_94_17) );
AOI211_X1 g_91_17 (.ZN (n_91_17), .A (n_87_15), .B (n_93_16), .C1 (n_93_18), .C2 (n_96_18) );
AOI211_X1 g_89_18 (.ZN (n_89_18), .A (n_89_16), .B (n_91_15), .C1 (n_95_17), .C2 (n_97_20) );
AOI211_X1 g_90_16 (.ZN (n_90_16), .A (n_91_17), .B (n_89_14), .C1 (n_93_16), .C2 (n_95_19) );
AOI211_X1 g_88_15 (.ZN (n_88_15), .A (n_89_18), .B (n_87_15), .C1 (n_91_15), .C2 (n_93_18) );
AOI211_X1 g_86_14 (.ZN (n_86_14), .A (n_90_16), .B (n_89_16), .C1 (n_89_14), .C2 (n_95_17) );
AOI211_X1 g_84_13 (.ZN (n_84_13), .A (n_88_15), .B (n_91_17), .C1 (n_87_15), .C2 (n_93_16) );
AOI211_X1 g_82_12 (.ZN (n_82_12), .A (n_86_14), .B (n_89_18), .C1 (n_89_16), .C2 (n_91_15) );
AOI211_X1 g_80_13 (.ZN (n_80_13), .A (n_84_13), .B (n_90_16), .C1 (n_91_17), .C2 (n_89_14) );
AOI211_X1 g_78_14 (.ZN (n_78_14), .A (n_82_12), .B (n_88_15), .C1 (n_89_18), .C2 (n_87_15) );
AOI211_X1 g_76_15 (.ZN (n_76_15), .A (n_80_13), .B (n_86_14), .C1 (n_90_16), .C2 (n_89_16) );
AOI211_X1 g_74_16 (.ZN (n_74_16), .A (n_78_14), .B (n_84_13), .C1 (n_88_15), .C2 (n_91_17) );
AOI211_X1 g_72_17 (.ZN (n_72_17), .A (n_76_15), .B (n_82_12), .C1 (n_86_14), .C2 (n_89_18) );
AOI211_X1 g_70_18 (.ZN (n_70_18), .A (n_74_16), .B (n_80_13), .C1 (n_84_13), .C2 (n_90_16) );
AOI211_X1 g_68_19 (.ZN (n_68_19), .A (n_72_17), .B (n_78_14), .C1 (n_82_12), .C2 (n_88_15) );
AOI211_X1 g_66_20 (.ZN (n_66_20), .A (n_70_18), .B (n_76_15), .C1 (n_80_13), .C2 (n_86_14) );
AOI211_X1 g_64_21 (.ZN (n_64_21), .A (n_68_19), .B (n_74_16), .C1 (n_78_14), .C2 (n_84_13) );
AOI211_X1 g_63_23 (.ZN (n_63_23), .A (n_66_20), .B (n_72_17), .C1 (n_76_15), .C2 (n_82_12) );
AOI211_X1 g_62_21 (.ZN (n_62_21), .A (n_64_21), .B (n_70_18), .C1 (n_74_16), .C2 (n_80_13) );
AOI211_X1 g_64_20 (.ZN (n_64_20), .A (n_63_23), .B (n_68_19), .C1 (n_72_17), .C2 (n_78_14) );
AOI211_X1 g_66_19 (.ZN (n_66_19), .A (n_62_21), .B (n_66_20), .C1 (n_70_18), .C2 (n_76_15) );
AOI211_X1 g_68_20 (.ZN (n_68_20), .A (n_64_20), .B (n_64_21), .C1 (n_68_19), .C2 (n_74_16) );
AOI211_X1 g_66_21 (.ZN (n_66_21), .A (n_66_19), .B (n_63_23), .C1 (n_66_20), .C2 (n_72_17) );
AOI211_X1 g_64_22 (.ZN (n_64_22), .A (n_68_20), .B (n_62_21), .C1 (n_64_21), .C2 (n_70_18) );
AOI211_X1 g_62_23 (.ZN (n_62_23), .A (n_66_21), .B (n_64_20), .C1 (n_63_23), .C2 (n_68_19) );
AOI211_X1 g_60_22 (.ZN (n_60_22), .A (n_64_22), .B (n_66_19), .C1 (n_62_21), .C2 (n_66_20) );
AOI211_X1 g_58_23 (.ZN (n_58_23), .A (n_62_23), .B (n_68_20), .C1 (n_64_20), .C2 (n_64_21) );
AOI211_X1 g_56_24 (.ZN (n_56_24), .A (n_60_22), .B (n_66_21), .C1 (n_66_19), .C2 (n_63_23) );
AOI211_X1 g_54_25 (.ZN (n_54_25), .A (n_58_23), .B (n_64_22), .C1 (n_68_20), .C2 (n_62_21) );
AOI211_X1 g_52_26 (.ZN (n_52_26), .A (n_56_24), .B (n_62_23), .C1 (n_66_21), .C2 (n_64_20) );
AOI211_X1 g_50_27 (.ZN (n_50_27), .A (n_54_25), .B (n_60_22), .C1 (n_64_22), .C2 (n_66_19) );
AOI211_X1 g_48_28 (.ZN (n_48_28), .A (n_52_26), .B (n_58_23), .C1 (n_62_23), .C2 (n_68_20) );
AOI211_X1 g_46_29 (.ZN (n_46_29), .A (n_50_27), .B (n_56_24), .C1 (n_60_22), .C2 (n_66_21) );
AOI211_X1 g_44_30 (.ZN (n_44_30), .A (n_48_28), .B (n_54_25), .C1 (n_58_23), .C2 (n_64_22) );
AOI211_X1 g_43_28 (.ZN (n_43_28), .A (n_46_29), .B (n_52_26), .C1 (n_56_24), .C2 (n_62_23) );
AOI211_X1 g_41_29 (.ZN (n_41_29), .A (n_44_30), .B (n_50_27), .C1 (n_54_25), .C2 (n_60_22) );
AOI211_X1 g_39_30 (.ZN (n_39_30), .A (n_43_28), .B (n_48_28), .C1 (n_52_26), .C2 (n_58_23) );
AOI211_X1 g_37_31 (.ZN (n_37_31), .A (n_41_29), .B (n_46_29), .C1 (n_50_27), .C2 (n_56_24) );
AOI211_X1 g_35_32 (.ZN (n_35_32), .A (n_39_30), .B (n_44_30), .C1 (n_48_28), .C2 (n_54_25) );
AOI211_X1 g_34_34 (.ZN (n_34_34), .A (n_37_31), .B (n_43_28), .C1 (n_46_29), .C2 (n_52_26) );
AOI211_X1 g_36_33 (.ZN (n_36_33), .A (n_35_32), .B (n_41_29), .C1 (n_44_30), .C2 (n_50_27) );
AOI211_X1 g_34_32 (.ZN (n_34_32), .A (n_34_34), .B (n_39_30), .C1 (n_43_28), .C2 (n_48_28) );
AOI211_X1 g_36_31 (.ZN (n_36_31), .A (n_36_33), .B (n_37_31), .C1 (n_41_29), .C2 (n_46_29) );
AOI211_X1 g_38_30 (.ZN (n_38_30), .A (n_34_32), .B (n_35_32), .C1 (n_39_30), .C2 (n_44_30) );
AOI211_X1 g_37_32 (.ZN (n_37_32), .A (n_36_31), .B (n_34_34), .C1 (n_37_31), .C2 (n_43_28) );
AOI211_X1 g_39_31 (.ZN (n_39_31), .A (n_38_30), .B (n_36_33), .C1 (n_35_32), .C2 (n_41_29) );
AOI211_X1 g_41_30 (.ZN (n_41_30), .A (n_37_32), .B (n_34_32), .C1 (n_34_34), .C2 (n_39_30) );
AOI211_X1 g_43_31 (.ZN (n_43_31), .A (n_39_31), .B (n_36_31), .C1 (n_36_33), .C2 (n_37_31) );
AOI211_X1 g_45_30 (.ZN (n_45_30), .A (n_41_30), .B (n_38_30), .C1 (n_34_32), .C2 (n_35_32) );
AOI211_X1 g_47_29 (.ZN (n_47_29), .A (n_43_31), .B (n_37_32), .C1 (n_36_31), .C2 (n_34_34) );
AOI211_X1 g_46_31 (.ZN (n_46_31), .A (n_45_30), .B (n_39_31), .C1 (n_38_30), .C2 (n_36_33) );
AOI211_X1 g_45_29 (.ZN (n_45_29), .A (n_47_29), .B (n_41_30), .C1 (n_37_32), .C2 (n_34_32) );
AOI211_X1 g_47_28 (.ZN (n_47_28), .A (n_46_31), .B (n_43_31), .C1 (n_39_31), .C2 (n_36_31) );
AOI211_X1 g_49_27 (.ZN (n_49_27), .A (n_45_29), .B (n_45_30), .C1 (n_41_30), .C2 (n_38_30) );
AOI211_X1 g_51_26 (.ZN (n_51_26), .A (n_47_28), .B (n_47_29), .C1 (n_43_31), .C2 (n_37_32) );
AOI211_X1 g_53_25 (.ZN (n_53_25), .A (n_49_27), .B (n_46_31), .C1 (n_45_30), .C2 (n_39_31) );
AOI211_X1 g_52_27 (.ZN (n_52_27), .A (n_51_26), .B (n_45_29), .C1 (n_47_29), .C2 (n_41_30) );
AOI211_X1 g_54_26 (.ZN (n_54_26), .A (n_53_25), .B (n_47_28), .C1 (n_46_31), .C2 (n_43_31) );
AOI211_X1 g_56_25 (.ZN (n_56_25), .A (n_52_27), .B (n_49_27), .C1 (n_45_29), .C2 (n_45_30) );
AOI211_X1 g_58_24 (.ZN (n_58_24), .A (n_54_26), .B (n_51_26), .C1 (n_47_28), .C2 (n_47_29) );
AOI211_X1 g_60_23 (.ZN (n_60_23), .A (n_56_25), .B (n_53_25), .C1 (n_49_27), .C2 (n_46_31) );
AOI211_X1 g_59_25 (.ZN (n_59_25), .A (n_58_24), .B (n_52_27), .C1 (n_51_26), .C2 (n_45_29) );
AOI211_X1 g_61_24 (.ZN (n_61_24), .A (n_60_23), .B (n_54_26), .C1 (n_53_25), .C2 (n_47_28) );
AOI211_X1 g_63_25 (.ZN (n_63_25), .A (n_59_25), .B (n_56_25), .C1 (n_52_27), .C2 (n_49_27) );
AOI211_X1 g_65_24 (.ZN (n_65_24), .A (n_61_24), .B (n_58_24), .C1 (n_54_26), .C2 (n_51_26) );
AOI211_X1 g_66_22 (.ZN (n_66_22), .A (n_63_25), .B (n_60_23), .C1 (n_56_25), .C2 (n_53_25) );
AOI211_X1 g_67_20 (.ZN (n_67_20), .A (n_65_24), .B (n_59_25), .C1 (n_58_24), .C2 (n_52_27) );
AOI211_X1 g_69_19 (.ZN (n_69_19), .A (n_66_22), .B (n_61_24), .C1 (n_60_23), .C2 (n_54_26) );
AOI211_X1 g_71_18 (.ZN (n_71_18), .A (n_67_20), .B (n_63_25), .C1 (n_59_25), .C2 (n_56_25) );
AOI211_X1 g_73_17 (.ZN (n_73_17), .A (n_69_19), .B (n_65_24), .C1 (n_61_24), .C2 (n_58_24) );
AOI211_X1 g_75_16 (.ZN (n_75_16), .A (n_71_18), .B (n_66_22), .C1 (n_63_25), .C2 (n_60_23) );
AOI211_X1 g_77_15 (.ZN (n_77_15), .A (n_73_17), .B (n_67_20), .C1 (n_65_24), .C2 (n_59_25) );
AOI211_X1 g_79_14 (.ZN (n_79_14), .A (n_75_16), .B (n_69_19), .C1 (n_66_22), .C2 (n_61_24) );
AOI211_X1 g_78_16 (.ZN (n_78_16), .A (n_77_15), .B (n_71_18), .C1 (n_67_20), .C2 (n_63_25) );
AOI211_X1 g_80_15 (.ZN (n_80_15), .A (n_79_14), .B (n_73_17), .C1 (n_69_19), .C2 (n_65_24) );
AOI211_X1 g_82_14 (.ZN (n_82_14), .A (n_78_16), .B (n_75_16), .C1 (n_71_18), .C2 (n_66_22) );
AOI211_X1 g_84_15 (.ZN (n_84_15), .A (n_80_15), .B (n_77_15), .C1 (n_73_17), .C2 (n_67_20) );
AOI211_X1 g_86_16 (.ZN (n_86_16), .A (n_82_14), .B (n_79_14), .C1 (n_75_16), .C2 (n_69_19) );
AOI211_X1 g_87_14 (.ZN (n_87_14), .A (n_84_15), .B (n_78_16), .C1 (n_77_15), .C2 (n_71_18) );
AOI211_X1 g_88_16 (.ZN (n_88_16), .A (n_86_16), .B (n_80_15), .C1 (n_79_14), .C2 (n_73_17) );
AOI211_X1 g_90_17 (.ZN (n_90_17), .A (n_87_14), .B (n_82_14), .C1 (n_78_16), .C2 (n_75_16) );
AOI211_X1 g_89_15 (.ZN (n_89_15), .A (n_88_16), .B (n_84_15), .C1 (n_80_15), .C2 (n_77_15) );
AOI211_X1 g_88_17 (.ZN (n_88_17), .A (n_90_17), .B (n_86_16), .C1 (n_82_14), .C2 (n_79_14) );
AOI211_X1 g_87_19 (.ZN (n_87_19), .A (n_89_15), .B (n_87_14), .C1 (n_84_15), .C2 (n_78_16) );
AOI211_X1 g_86_17 (.ZN (n_86_17), .A (n_88_17), .B (n_88_16), .C1 (n_86_16), .C2 (n_80_15) );
AOI211_X1 g_85_15 (.ZN (n_85_15), .A (n_87_19), .B (n_90_17), .C1 (n_87_14), .C2 (n_82_14) );
AOI211_X1 g_83_14 (.ZN (n_83_14), .A (n_86_17), .B (n_89_15), .C1 (n_88_16), .C2 (n_84_15) );
AOI211_X1 g_84_16 (.ZN (n_84_16), .A (n_85_15), .B (n_88_17), .C1 (n_90_17), .C2 (n_86_16) );
AOI211_X1 g_85_18 (.ZN (n_85_18), .A (n_83_14), .B (n_87_19), .C1 (n_89_15), .C2 (n_87_14) );
AOI211_X1 g_87_17 (.ZN (n_87_17), .A (n_84_16), .B (n_86_17), .C1 (n_88_17), .C2 (n_88_16) );
AOI211_X1 g_85_16 (.ZN (n_85_16), .A (n_85_18), .B (n_85_15), .C1 (n_87_19), .C2 (n_90_17) );
AOI211_X1 g_83_15 (.ZN (n_83_15), .A (n_87_17), .B (n_83_14), .C1 (n_86_17), .C2 (n_89_15) );
AOI211_X1 g_81_14 (.ZN (n_81_14), .A (n_85_16), .B (n_84_16), .C1 (n_85_15), .C2 (n_88_17) );
AOI211_X1 g_79_15 (.ZN (n_79_15), .A (n_83_15), .B (n_85_18), .C1 (n_83_14), .C2 (n_87_19) );
AOI211_X1 g_77_16 (.ZN (n_77_16), .A (n_81_14), .B (n_87_17), .C1 (n_84_16), .C2 (n_86_17) );
AOI211_X1 g_75_17 (.ZN (n_75_17), .A (n_79_15), .B (n_85_16), .C1 (n_85_18), .C2 (n_85_15) );
AOI211_X1 g_73_18 (.ZN (n_73_18), .A (n_77_16), .B (n_83_15), .C1 (n_87_17), .C2 (n_83_14) );
AOI211_X1 g_71_19 (.ZN (n_71_19), .A (n_75_17), .B (n_81_14), .C1 (n_85_16), .C2 (n_84_16) );
AOI211_X1 g_69_20 (.ZN (n_69_20), .A (n_73_18), .B (n_79_15), .C1 (n_83_15), .C2 (n_85_18) );
AOI211_X1 g_67_21 (.ZN (n_67_21), .A (n_71_19), .B (n_77_16), .C1 (n_81_14), .C2 (n_87_17) );
AOI211_X1 g_65_22 (.ZN (n_65_22), .A (n_69_20), .B (n_75_17), .C1 (n_79_15), .C2 (n_85_16) );
AOI211_X1 g_67_23 (.ZN (n_67_23), .A (n_67_21), .B (n_73_18), .C1 (n_77_16), .C2 (n_83_15) );
AOI211_X1 g_68_21 (.ZN (n_68_21), .A (n_65_22), .B (n_71_19), .C1 (n_75_17), .C2 (n_81_14) );
AOI211_X1 g_70_20 (.ZN (n_70_20), .A (n_67_23), .B (n_69_20), .C1 (n_73_18), .C2 (n_79_15) );
AOI211_X1 g_72_19 (.ZN (n_72_19), .A (n_68_21), .B (n_67_21), .C1 (n_71_19), .C2 (n_77_16) );
AOI211_X1 g_74_18 (.ZN (n_74_18), .A (n_70_20), .B (n_65_22), .C1 (n_69_20), .C2 (n_75_17) );
AOI211_X1 g_76_17 (.ZN (n_76_17), .A (n_72_19), .B (n_67_23), .C1 (n_67_21), .C2 (n_73_18) );
AOI211_X1 g_75_19 (.ZN (n_75_19), .A (n_74_18), .B (n_68_21), .C1 (n_65_22), .C2 (n_71_19) );
AOI211_X1 g_77_18 (.ZN (n_77_18), .A (n_76_17), .B (n_70_20), .C1 (n_67_23), .C2 (n_69_20) );
AOI211_X1 g_79_17 (.ZN (n_79_17), .A (n_75_19), .B (n_72_19), .C1 (n_68_21), .C2 (n_67_21) );
AOI211_X1 g_81_16 (.ZN (n_81_16), .A (n_77_18), .B (n_74_18), .C1 (n_70_20), .C2 (n_65_22) );
AOI211_X1 g_83_17 (.ZN (n_83_17), .A (n_79_17), .B (n_76_17), .C1 (n_72_19), .C2 (n_67_23) );
AOI211_X1 g_81_18 (.ZN (n_81_18), .A (n_81_16), .B (n_75_19), .C1 (n_74_18), .C2 (n_68_21) );
AOI211_X1 g_82_16 (.ZN (n_82_16), .A (n_83_17), .B (n_77_18), .C1 (n_76_17), .C2 (n_70_20) );
AOI211_X1 g_84_17 (.ZN (n_84_17), .A (n_81_18), .B (n_79_17), .C1 (n_75_19), .C2 (n_72_19) );
AOI211_X1 g_83_19 (.ZN (n_83_19), .A (n_82_16), .B (n_81_16), .C1 (n_77_18), .C2 (n_74_18) );
AOI211_X1 g_82_17 (.ZN (n_82_17), .A (n_84_17), .B (n_83_17), .C1 (n_79_17), .C2 (n_76_17) );
AOI211_X1 g_80_16 (.ZN (n_80_16), .A (n_83_19), .B (n_81_18), .C1 (n_81_16), .C2 (n_75_19) );
AOI211_X1 g_78_17 (.ZN (n_78_17), .A (n_82_17), .B (n_82_16), .C1 (n_83_17), .C2 (n_77_18) );
AOI211_X1 g_76_18 (.ZN (n_76_18), .A (n_80_16), .B (n_84_17), .C1 (n_81_18), .C2 (n_79_17) );
AOI211_X1 g_74_19 (.ZN (n_74_19), .A (n_78_17), .B (n_83_19), .C1 (n_82_16), .C2 (n_81_16) );
AOI211_X1 g_72_20 (.ZN (n_72_20), .A (n_76_18), .B (n_82_17), .C1 (n_84_17), .C2 (n_83_17) );
AOI211_X1 g_70_21 (.ZN (n_70_21), .A (n_74_19), .B (n_80_16), .C1 (n_83_19), .C2 (n_81_18) );
AOI211_X1 g_68_22 (.ZN (n_68_22), .A (n_72_20), .B (n_78_17), .C1 (n_82_17), .C2 (n_82_16) );
AOI211_X1 g_66_23 (.ZN (n_66_23), .A (n_70_21), .B (n_76_18), .C1 (n_80_16), .C2 (n_84_17) );
AOI211_X1 g_65_21 (.ZN (n_65_21), .A (n_68_22), .B (n_74_19), .C1 (n_78_17), .C2 (n_83_19) );
AOI211_X1 g_64_23 (.ZN (n_64_23), .A (n_66_23), .B (n_72_20), .C1 (n_76_18), .C2 (n_82_17) );
AOI211_X1 g_62_24 (.ZN (n_62_24), .A (n_65_21), .B (n_70_21), .C1 (n_74_19), .C2 (n_80_16) );
AOI211_X1 g_63_22 (.ZN (n_63_22), .A (n_64_23), .B (n_68_22), .C1 (n_72_20), .C2 (n_78_17) );
AOI211_X1 g_61_23 (.ZN (n_61_23), .A (n_62_24), .B (n_66_23), .C1 (n_70_21), .C2 (n_76_18) );
AOI211_X1 g_59_24 (.ZN (n_59_24), .A (n_63_22), .B (n_65_21), .C1 (n_68_22), .C2 (n_74_19) );
AOI211_X1 g_57_25 (.ZN (n_57_25), .A (n_61_23), .B (n_64_23), .C1 (n_66_23), .C2 (n_72_20) );
AOI211_X1 g_55_26 (.ZN (n_55_26), .A (n_59_24), .B (n_62_24), .C1 (n_65_21), .C2 (n_70_21) );
AOI211_X1 g_53_27 (.ZN (n_53_27), .A (n_57_25), .B (n_63_22), .C1 (n_64_23), .C2 (n_68_22) );
AOI211_X1 g_51_28 (.ZN (n_51_28), .A (n_55_26), .B (n_61_23), .C1 (n_62_24), .C2 (n_66_23) );
AOI211_X1 g_49_29 (.ZN (n_49_29), .A (n_53_27), .B (n_59_24), .C1 (n_63_22), .C2 (n_65_21) );
AOI211_X1 g_47_30 (.ZN (n_47_30), .A (n_51_28), .B (n_57_25), .C1 (n_61_23), .C2 (n_64_23) );
AOI211_X1 g_45_31 (.ZN (n_45_31), .A (n_49_29), .B (n_55_26), .C1 (n_59_24), .C2 (n_62_24) );
AOI211_X1 g_43_30 (.ZN (n_43_30), .A (n_47_30), .B (n_53_27), .C1 (n_57_25), .C2 (n_63_22) );
AOI211_X1 g_41_31 (.ZN (n_41_31), .A (n_45_31), .B (n_51_28), .C1 (n_55_26), .C2 (n_61_23) );
AOI211_X1 g_39_32 (.ZN (n_39_32), .A (n_43_30), .B (n_49_29), .C1 (n_53_27), .C2 (n_59_24) );
AOI211_X1 g_37_33 (.ZN (n_37_33), .A (n_41_31), .B (n_47_30), .C1 (n_51_28), .C2 (n_57_25) );
AOI211_X1 g_38_31 (.ZN (n_38_31), .A (n_39_32), .B (n_45_31), .C1 (n_49_29), .C2 (n_55_26) );
AOI211_X1 g_36_32 (.ZN (n_36_32), .A (n_37_33), .B (n_43_30), .C1 (n_47_30), .C2 (n_53_27) );
AOI211_X1 g_34_33 (.ZN (n_34_33), .A (n_38_31), .B (n_41_31), .C1 (n_45_31), .C2 (n_51_28) );
AOI211_X1 g_36_34 (.ZN (n_36_34), .A (n_36_32), .B (n_39_32), .C1 (n_43_30), .C2 (n_49_29) );
AOI211_X1 g_38_33 (.ZN (n_38_33), .A (n_34_33), .B (n_37_33), .C1 (n_41_31), .C2 (n_47_30) );
AOI211_X1 g_40_32 (.ZN (n_40_32), .A (n_36_34), .B (n_38_31), .C1 (n_39_32), .C2 (n_45_31) );
AOI211_X1 g_42_31 (.ZN (n_42_31), .A (n_38_33), .B (n_36_32), .C1 (n_37_33), .C2 (n_43_30) );
AOI211_X1 g_44_32 (.ZN (n_44_32), .A (n_40_32), .B (n_34_33), .C1 (n_38_31), .C2 (n_41_31) );
AOI211_X1 g_42_33 (.ZN (n_42_33), .A (n_42_31), .B (n_36_34), .C1 (n_36_32), .C2 (n_39_32) );
AOI211_X1 g_40_34 (.ZN (n_40_34), .A (n_44_32), .B (n_38_33), .C1 (n_34_33), .C2 (n_37_33) );
AOI211_X1 g_41_32 (.ZN (n_41_32), .A (n_42_33), .B (n_40_32), .C1 (n_36_34), .C2 (n_38_31) );
AOI211_X1 g_42_30 (.ZN (n_42_30), .A (n_40_34), .B (n_42_31), .C1 (n_38_33), .C2 (n_36_32) );
AOI211_X1 g_40_31 (.ZN (n_40_31), .A (n_41_32), .B (n_44_32), .C1 (n_40_32), .C2 (n_34_33) );
AOI211_X1 g_38_32 (.ZN (n_38_32), .A (n_42_30), .B (n_42_33), .C1 (n_42_31), .C2 (n_36_34) );
AOI211_X1 g_39_34 (.ZN (n_39_34), .A (n_40_31), .B (n_40_34), .C1 (n_44_32), .C2 (n_38_33) );
AOI211_X1 g_41_33 (.ZN (n_41_33), .A (n_38_32), .B (n_41_32), .C1 (n_42_33), .C2 (n_40_32) );
AOI211_X1 g_43_32 (.ZN (n_43_32), .A (n_39_34), .B (n_42_30), .C1 (n_40_34), .C2 (n_42_31) );
AOI211_X1 g_42_34 (.ZN (n_42_34), .A (n_41_33), .B (n_40_31), .C1 (n_41_32), .C2 (n_44_32) );
AOI211_X1 g_40_33 (.ZN (n_40_33), .A (n_43_32), .B (n_38_32), .C1 (n_42_30), .C2 (n_42_33) );
AOI211_X1 g_42_32 (.ZN (n_42_32), .A (n_42_34), .B (n_39_34), .C1 (n_40_31), .C2 (n_40_34) );
AOI211_X1 g_44_31 (.ZN (n_44_31), .A (n_40_33), .B (n_41_33), .C1 (n_38_32), .C2 (n_41_32) );
AOI211_X1 g_46_30 (.ZN (n_46_30), .A (n_42_32), .B (n_43_32), .C1 (n_39_34), .C2 (n_42_30) );
AOI211_X1 g_48_29 (.ZN (n_48_29), .A (n_44_31), .B (n_42_34), .C1 (n_41_33), .C2 (n_40_31) );
AOI211_X1 g_50_28 (.ZN (n_50_28), .A (n_46_30), .B (n_40_33), .C1 (n_43_32), .C2 (n_38_32) );
AOI211_X1 g_49_30 (.ZN (n_49_30), .A (n_48_29), .B (n_42_32), .C1 (n_42_34), .C2 (n_39_34) );
AOI211_X1 g_51_29 (.ZN (n_51_29), .A (n_50_28), .B (n_44_31), .C1 (n_40_33), .C2 (n_41_33) );
AOI211_X1 g_53_28 (.ZN (n_53_28), .A (n_49_30), .B (n_46_30), .C1 (n_42_32), .C2 (n_43_32) );
AOI211_X1 g_55_27 (.ZN (n_55_27), .A (n_51_29), .B (n_48_29), .C1 (n_44_31), .C2 (n_42_34) );
AOI211_X1 g_57_26 (.ZN (n_57_26), .A (n_53_28), .B (n_50_28), .C1 (n_46_30), .C2 (n_40_33) );
AOI211_X1 g_56_28 (.ZN (n_56_28), .A (n_55_27), .B (n_49_30), .C1 (n_48_29), .C2 (n_42_32) );
AOI211_X1 g_54_27 (.ZN (n_54_27), .A (n_57_26), .B (n_51_29), .C1 (n_50_28), .C2 (n_44_31) );
AOI211_X1 g_56_26 (.ZN (n_56_26), .A (n_56_28), .B (n_53_28), .C1 (n_49_30), .C2 (n_46_30) );
AOI211_X1 g_58_25 (.ZN (n_58_25), .A (n_54_27), .B (n_55_27), .C1 (n_51_29), .C2 (n_48_29) );
AOI211_X1 g_60_24 (.ZN (n_60_24), .A (n_56_26), .B (n_57_26), .C1 (n_53_28), .C2 (n_50_28) );
AOI211_X1 g_61_26 (.ZN (n_61_26), .A (n_58_25), .B (n_56_28), .C1 (n_55_27), .C2 (n_49_30) );
AOI211_X1 g_59_27 (.ZN (n_59_27), .A (n_60_24), .B (n_54_27), .C1 (n_57_26), .C2 (n_51_29) );
AOI211_X1 g_60_25 (.ZN (n_60_25), .A (n_61_26), .B (n_56_26), .C1 (n_56_28), .C2 (n_53_28) );
AOI211_X1 g_58_26 (.ZN (n_58_26), .A (n_59_27), .B (n_58_25), .C1 (n_54_27), .C2 (n_55_27) );
AOI211_X1 g_56_27 (.ZN (n_56_27), .A (n_60_25), .B (n_60_24), .C1 (n_56_26), .C2 (n_57_26) );
AOI211_X1 g_54_28 (.ZN (n_54_28), .A (n_58_26), .B (n_61_26), .C1 (n_58_25), .C2 (n_56_28) );
AOI211_X1 g_52_29 (.ZN (n_52_29), .A (n_56_27), .B (n_59_27), .C1 (n_60_24), .C2 (n_54_27) );
AOI211_X1 g_50_30 (.ZN (n_50_30), .A (n_54_28), .B (n_60_25), .C1 (n_61_26), .C2 (n_56_26) );
AOI211_X1 g_48_31 (.ZN (n_48_31), .A (n_52_29), .B (n_58_26), .C1 (n_59_27), .C2 (n_58_25) );
AOI211_X1 g_46_32 (.ZN (n_46_32), .A (n_50_30), .B (n_56_27), .C1 (n_60_25), .C2 (n_60_24) );
AOI211_X1 g_44_33 (.ZN (n_44_33), .A (n_48_31), .B (n_54_28), .C1 (n_58_26), .C2 (n_61_26) );
AOI211_X1 g_43_35 (.ZN (n_43_35), .A (n_46_32), .B (n_52_29), .C1 (n_56_27), .C2 (n_59_27) );
AOI211_X1 g_45_34 (.ZN (n_45_34), .A (n_44_33), .B (n_50_30), .C1 (n_54_28), .C2 (n_60_25) );
AOI211_X1 g_43_33 (.ZN (n_43_33), .A (n_43_35), .B (n_48_31), .C1 (n_52_29), .C2 (n_58_26) );
AOI211_X1 g_45_32 (.ZN (n_45_32), .A (n_45_34), .B (n_46_32), .C1 (n_50_30), .C2 (n_56_27) );
AOI211_X1 g_47_31 (.ZN (n_47_31), .A (n_43_33), .B (n_44_33), .C1 (n_48_31), .C2 (n_54_28) );
AOI211_X1 g_46_33 (.ZN (n_46_33), .A (n_45_32), .B (n_43_35), .C1 (n_46_32), .C2 (n_52_29) );
AOI211_X1 g_48_32 (.ZN (n_48_32), .A (n_47_31), .B (n_45_34), .C1 (n_44_33), .C2 (n_50_30) );
AOI211_X1 g_50_31 (.ZN (n_50_31), .A (n_46_33), .B (n_43_33), .C1 (n_43_35), .C2 (n_48_31) );
AOI211_X1 g_48_30 (.ZN (n_48_30), .A (n_48_32), .B (n_45_32), .C1 (n_45_34), .C2 (n_46_32) );
AOI211_X1 g_50_29 (.ZN (n_50_29), .A (n_50_31), .B (n_47_31), .C1 (n_43_33), .C2 (n_44_33) );
AOI211_X1 g_52_28 (.ZN (n_52_28), .A (n_48_30), .B (n_46_33), .C1 (n_45_32), .C2 (n_43_35) );
AOI211_X1 g_54_29 (.ZN (n_54_29), .A (n_50_29), .B (n_48_32), .C1 (n_47_31), .C2 (n_45_34) );
AOI211_X1 g_52_30 (.ZN (n_52_30), .A (n_52_28), .B (n_50_31), .C1 (n_46_33), .C2 (n_43_33) );
AOI211_X1 g_51_32 (.ZN (n_51_32), .A (n_54_29), .B (n_48_30), .C1 (n_48_32), .C2 (n_45_32) );
AOI211_X1 g_49_31 (.ZN (n_49_31), .A (n_52_30), .B (n_50_29), .C1 (n_50_31), .C2 (n_47_31) );
AOI211_X1 g_51_30 (.ZN (n_51_30), .A (n_51_32), .B (n_52_28), .C1 (n_48_30), .C2 (n_46_33) );
AOI211_X1 g_53_29 (.ZN (n_53_29), .A (n_49_31), .B (n_54_29), .C1 (n_50_29), .C2 (n_48_32) );
AOI211_X1 g_55_28 (.ZN (n_55_28), .A (n_51_30), .B (n_52_30), .C1 (n_52_28), .C2 (n_50_31) );
AOI211_X1 g_57_27 (.ZN (n_57_27), .A (n_53_29), .B (n_51_32), .C1 (n_54_29), .C2 (n_48_30) );
AOI211_X1 g_59_26 (.ZN (n_59_26), .A (n_55_28), .B (n_49_31), .C1 (n_52_30), .C2 (n_50_29) );
AOI211_X1 g_61_25 (.ZN (n_61_25), .A (n_57_27), .B (n_51_30), .C1 (n_51_32), .C2 (n_52_28) );
AOI211_X1 g_63_24 (.ZN (n_63_24), .A (n_59_26), .B (n_53_29), .C1 (n_49_31), .C2 (n_54_29) );
AOI211_X1 g_65_23 (.ZN (n_65_23), .A (n_61_25), .B (n_55_28), .C1 (n_51_30), .C2 (n_52_30) );
AOI211_X1 g_67_22 (.ZN (n_67_22), .A (n_63_24), .B (n_57_27), .C1 (n_53_29), .C2 (n_51_32) );
AOI211_X1 g_69_21 (.ZN (n_69_21), .A (n_65_23), .B (n_59_26), .C1 (n_55_28), .C2 (n_49_31) );
AOI211_X1 g_71_20 (.ZN (n_71_20), .A (n_67_22), .B (n_61_25), .C1 (n_57_27), .C2 (n_51_30) );
AOI211_X1 g_73_19 (.ZN (n_73_19), .A (n_69_21), .B (n_63_24), .C1 (n_59_26), .C2 (n_53_29) );
AOI211_X1 g_75_18 (.ZN (n_75_18), .A (n_71_20), .B (n_65_23), .C1 (n_61_25), .C2 (n_55_28) );
AOI211_X1 g_77_17 (.ZN (n_77_17), .A (n_73_19), .B (n_67_22), .C1 (n_63_24), .C2 (n_57_27) );
AOI211_X1 g_79_16 (.ZN (n_79_16), .A (n_75_18), .B (n_69_21), .C1 (n_65_23), .C2 (n_59_26) );
AOI211_X1 g_81_15 (.ZN (n_81_15), .A (n_77_17), .B (n_71_20), .C1 (n_67_22), .C2 (n_61_25) );
AOI211_X1 g_80_17 (.ZN (n_80_17), .A (n_79_16), .B (n_73_19), .C1 (n_69_21), .C2 (n_63_24) );
AOI211_X1 g_78_18 (.ZN (n_78_18), .A (n_81_15), .B (n_75_18), .C1 (n_71_20), .C2 (n_65_23) );
AOI211_X1 g_76_19 (.ZN (n_76_19), .A (n_80_17), .B (n_77_17), .C1 (n_73_19), .C2 (n_67_22) );
AOI211_X1 g_74_20 (.ZN (n_74_20), .A (n_78_18), .B (n_79_16), .C1 (n_75_18), .C2 (n_69_21) );
AOI211_X1 g_72_21 (.ZN (n_72_21), .A (n_76_19), .B (n_81_15), .C1 (n_77_17), .C2 (n_71_20) );
AOI211_X1 g_70_22 (.ZN (n_70_22), .A (n_74_20), .B (n_80_17), .C1 (n_79_16), .C2 (n_73_19) );
AOI211_X1 g_68_23 (.ZN (n_68_23), .A (n_72_21), .B (n_78_18), .C1 (n_81_15), .C2 (n_75_18) );
AOI211_X1 g_66_24 (.ZN (n_66_24), .A (n_70_22), .B (n_76_19), .C1 (n_80_17), .C2 (n_77_17) );
AOI211_X1 g_64_25 (.ZN (n_64_25), .A (n_68_23), .B (n_74_20), .C1 (n_78_18), .C2 (n_79_16) );
AOI211_X1 g_62_26 (.ZN (n_62_26), .A (n_66_24), .B (n_72_21), .C1 (n_76_19), .C2 (n_81_15) );
AOI211_X1 g_60_27 (.ZN (n_60_27), .A (n_64_25), .B (n_70_22), .C1 (n_74_20), .C2 (n_80_17) );
AOI211_X1 g_58_28 (.ZN (n_58_28), .A (n_62_26), .B (n_68_23), .C1 (n_72_21), .C2 (n_78_18) );
AOI211_X1 g_56_29 (.ZN (n_56_29), .A (n_60_27), .B (n_66_24), .C1 (n_70_22), .C2 (n_76_19) );
AOI211_X1 g_54_30 (.ZN (n_54_30), .A (n_58_28), .B (n_64_25), .C1 (n_68_23), .C2 (n_74_20) );
AOI211_X1 g_52_31 (.ZN (n_52_31), .A (n_56_29), .B (n_62_26), .C1 (n_66_24), .C2 (n_72_21) );
AOI211_X1 g_50_32 (.ZN (n_50_32), .A (n_54_30), .B (n_60_27), .C1 (n_64_25), .C2 (n_70_22) );
AOI211_X1 g_48_33 (.ZN (n_48_33), .A (n_52_31), .B (n_58_28), .C1 (n_62_26), .C2 (n_68_23) );
AOI211_X1 g_46_34 (.ZN (n_46_34), .A (n_50_32), .B (n_56_29), .C1 (n_60_27), .C2 (n_66_24) );
AOI211_X1 g_47_32 (.ZN (n_47_32), .A (n_48_33), .B (n_54_30), .C1 (n_58_28), .C2 (n_64_25) );
AOI211_X1 g_45_33 (.ZN (n_45_33), .A (n_46_34), .B (n_52_31), .C1 (n_56_29), .C2 (n_62_26) );
AOI211_X1 g_43_34 (.ZN (n_43_34), .A (n_47_32), .B (n_50_32), .C1 (n_54_30), .C2 (n_60_27) );
AOI211_X1 g_41_35 (.ZN (n_41_35), .A (n_45_33), .B (n_48_33), .C1 (n_52_31), .C2 (n_58_28) );
AOI211_X1 g_39_36 (.ZN (n_39_36), .A (n_43_34), .B (n_46_34), .C1 (n_50_32), .C2 (n_56_29) );
AOI211_X1 g_38_34 (.ZN (n_38_34), .A (n_41_35), .B (n_47_32), .C1 (n_48_33), .C2 (n_54_30) );
AOI211_X1 g_36_35 (.ZN (n_36_35), .A (n_39_36), .B (n_45_33), .C1 (n_46_34), .C2 (n_52_31) );
AOI211_X1 g_35_33 (.ZN (n_35_33), .A (n_38_34), .B (n_43_34), .C1 (n_47_32), .C2 (n_50_32) );
AOI211_X1 g_34_35 (.ZN (n_34_35), .A (n_36_35), .B (n_41_35), .C1 (n_45_33), .C2 (n_48_33) );
AOI211_X1 g_35_37 (.ZN (n_35_37), .A (n_35_33), .B (n_39_36), .C1 (n_43_34), .C2 (n_46_34) );
AOI211_X1 g_37_36 (.ZN (n_37_36), .A (n_34_35), .B (n_38_34), .C1 (n_41_35), .C2 (n_47_32) );
AOI211_X1 g_39_35 (.ZN (n_39_35), .A (n_35_37), .B (n_36_35), .C1 (n_39_36), .C2 (n_45_33) );
AOI211_X1 g_41_34 (.ZN (n_41_34), .A (n_37_36), .B (n_35_33), .C1 (n_38_34), .C2 (n_43_34) );
AOI211_X1 g_39_33 (.ZN (n_39_33), .A (n_39_35), .B (n_34_35), .C1 (n_36_35), .C2 (n_41_35) );
AOI211_X1 g_37_34 (.ZN (n_37_34), .A (n_41_34), .B (n_35_37), .C1 (n_35_33), .C2 (n_39_36) );
AOI211_X1 g_35_35 (.ZN (n_35_35), .A (n_39_33), .B (n_37_36), .C1 (n_34_35), .C2 (n_38_34) );
AOI211_X1 g_33_34 (.ZN (n_33_34), .A (n_37_34), .B (n_39_35), .C1 (n_35_37), .C2 (n_36_35) );
AOI211_X1 g_31_33 (.ZN (n_31_33), .A (n_35_35), .B (n_41_34), .C1 (n_37_36), .C2 (n_35_33) );
AOI211_X1 g_29_34 (.ZN (n_29_34), .A (n_33_34), .B (n_39_33), .C1 (n_39_35), .C2 (n_34_35) );
AOI211_X1 g_30_32 (.ZN (n_30_32), .A (n_31_33), .B (n_37_34), .C1 (n_41_34), .C2 (n_35_37) );
AOI211_X1 g_32_33 (.ZN (n_32_33), .A (n_29_34), .B (n_35_35), .C1 (n_39_33), .C2 (n_37_36) );
AOI211_X1 g_31_35 (.ZN (n_31_35), .A (n_30_32), .B (n_33_34), .C1 (n_37_34), .C2 (n_39_35) );
AOI211_X1 g_33_36 (.ZN (n_33_36), .A (n_32_33), .B (n_31_33), .C1 (n_35_35), .C2 (n_41_34) );
AOI211_X1 g_31_37 (.ZN (n_31_37), .A (n_31_35), .B (n_29_34), .C1 (n_33_34), .C2 (n_39_33) );
AOI211_X1 g_32_35 (.ZN (n_32_35), .A (n_33_36), .B (n_30_32), .C1 (n_31_33), .C2 (n_37_34) );
AOI211_X1 g_30_34 (.ZN (n_30_34), .A (n_31_37), .B (n_32_33), .C1 (n_29_34), .C2 (n_35_35) );
AOI211_X1 g_28_33 (.ZN (n_28_33), .A (n_32_35), .B (n_31_35), .C1 (n_30_32), .C2 (n_33_34) );
AOI211_X1 g_26_34 (.ZN (n_26_34), .A (n_30_34), .B (n_33_36), .C1 (n_32_33), .C2 (n_31_33) );
AOI211_X1 g_24_35 (.ZN (n_24_35), .A (n_28_33), .B (n_31_37), .C1 (n_31_35), .C2 (n_29_34) );
AOI211_X1 g_22_36 (.ZN (n_22_36), .A (n_26_34), .B (n_32_35), .C1 (n_33_36), .C2 (n_30_32) );
AOI211_X1 g_20_37 (.ZN (n_20_37), .A (n_24_35), .B (n_30_34), .C1 (n_31_37), .C2 (n_32_33) );
AOI211_X1 g_18_38 (.ZN (n_18_38), .A (n_22_36), .B (n_28_33), .C1 (n_32_35), .C2 (n_31_35) );
AOI211_X1 g_16_39 (.ZN (n_16_39), .A (n_20_37), .B (n_26_34), .C1 (n_30_34), .C2 (n_33_36) );
AOI211_X1 g_14_40 (.ZN (n_14_40), .A (n_18_38), .B (n_24_35), .C1 (n_28_33), .C2 (n_31_37) );
AOI211_X1 g_12_41 (.ZN (n_12_41), .A (n_16_39), .B (n_22_36), .C1 (n_26_34), .C2 (n_32_35) );
AOI211_X1 g_10_42 (.ZN (n_10_42), .A (n_14_40), .B (n_20_37), .C1 (n_24_35), .C2 (n_30_34) );
AOI211_X1 g_8_41 (.ZN (n_8_41), .A (n_12_41), .B (n_18_38), .C1 (n_22_36), .C2 (n_28_33) );
AOI211_X1 g_6_42 (.ZN (n_6_42), .A (n_10_42), .B (n_16_39), .C1 (n_20_37), .C2 (n_26_34) );
AOI211_X1 g_5_44 (.ZN (n_5_44), .A (n_8_41), .B (n_14_40), .C1 (n_18_38), .C2 (n_24_35) );
AOI211_X1 g_7_43 (.ZN (n_7_43), .A (n_6_42), .B (n_12_41), .C1 (n_16_39), .C2 (n_22_36) );
AOI211_X1 g_9_44 (.ZN (n_9_44), .A (n_5_44), .B (n_10_42), .C1 (n_14_40), .C2 (n_20_37) );
AOI211_X1 g_7_45 (.ZN (n_7_45), .A (n_7_43), .B (n_8_41), .C1 (n_12_41), .C2 (n_18_38) );
AOI211_X1 g_8_43 (.ZN (n_8_43), .A (n_9_44), .B (n_6_42), .C1 (n_10_42), .C2 (n_16_39) );
AOI211_X1 g_9_45 (.ZN (n_9_45), .A (n_7_45), .B (n_5_44), .C1 (n_8_41), .C2 (n_14_40) );
AOI211_X1 g_10_43 (.ZN (n_10_43), .A (n_8_43), .B (n_7_43), .C1 (n_6_42), .C2 (n_12_41) );
AOI211_X1 g_12_42 (.ZN (n_12_42), .A (n_9_45), .B (n_9_44), .C1 (n_5_44), .C2 (n_10_42) );
AOI211_X1 g_10_41 (.ZN (n_10_41), .A (n_10_43), .B (n_7_45), .C1 (n_7_43), .C2 (n_8_41) );
AOI211_X1 g_12_40 (.ZN (n_12_40), .A (n_12_42), .B (n_8_43), .C1 (n_9_44), .C2 (n_6_42) );
AOI211_X1 g_14_41 (.ZN (n_14_41), .A (n_10_41), .B (n_9_45), .C1 (n_7_45), .C2 (n_5_44) );
AOI211_X1 g_16_40 (.ZN (n_16_40), .A (n_12_40), .B (n_10_43), .C1 (n_8_43), .C2 (n_7_43) );
AOI211_X1 g_18_39 (.ZN (n_18_39), .A (n_14_41), .B (n_12_42), .C1 (n_9_45), .C2 (n_9_44) );
AOI211_X1 g_17_41 (.ZN (n_17_41), .A (n_16_40), .B (n_10_41), .C1 (n_10_43), .C2 (n_7_45) );
AOI211_X1 g_19_40 (.ZN (n_19_40), .A (n_18_39), .B (n_12_40), .C1 (n_12_42), .C2 (n_8_43) );
AOI211_X1 g_21_39 (.ZN (n_21_39), .A (n_17_41), .B (n_14_41), .C1 (n_10_41), .C2 (n_9_45) );
AOI211_X1 g_23_38 (.ZN (n_23_38), .A (n_19_40), .B (n_16_40), .C1 (n_12_40), .C2 (n_10_43) );
AOI211_X1 g_25_37 (.ZN (n_25_37), .A (n_21_39), .B (n_18_39), .C1 (n_14_41), .C2 (n_12_42) );
AOI211_X1 g_27_36 (.ZN (n_27_36), .A (n_23_38), .B (n_17_41), .C1 (n_16_40), .C2 (n_10_41) );
AOI211_X1 g_25_35 (.ZN (n_25_35), .A (n_25_37), .B (n_19_40), .C1 (n_18_39), .C2 (n_12_40) );
AOI211_X1 g_27_34 (.ZN (n_27_34), .A (n_27_36), .B (n_21_39), .C1 (n_17_41), .C2 (n_14_41) );
AOI211_X1 g_29_33 (.ZN (n_29_33), .A (n_25_35), .B (n_23_38), .C1 (n_19_40), .C2 (n_16_40) );
AOI211_X1 g_30_35 (.ZN (n_30_35), .A (n_27_34), .B (n_25_37), .C1 (n_21_39), .C2 (n_18_39) );
AOI211_X1 g_28_36 (.ZN (n_28_36), .A (n_29_33), .B (n_27_36), .C1 (n_23_38), .C2 (n_17_41) );
AOI211_X1 g_26_37 (.ZN (n_26_37), .A (n_30_35), .B (n_25_35), .C1 (n_25_37), .C2 (n_19_40) );
AOI211_X1 g_27_35 (.ZN (n_27_35), .A (n_28_36), .B (n_27_34), .C1 (n_27_36), .C2 (n_21_39) );
AOI211_X1 g_29_36 (.ZN (n_29_36), .A (n_26_37), .B (n_29_33), .C1 (n_25_35), .C2 (n_23_38) );
AOI211_X1 g_28_38 (.ZN (n_28_38), .A (n_27_35), .B (n_30_35), .C1 (n_27_34), .C2 (n_25_37) );
AOI211_X1 g_30_37 (.ZN (n_30_37), .A (n_29_36), .B (n_28_36), .C1 (n_29_33), .C2 (n_27_36) );
AOI211_X1 g_29_35 (.ZN (n_29_35), .A (n_28_38), .B (n_26_37), .C1 (n_30_35), .C2 (n_25_35) );
AOI211_X1 g_31_34 (.ZN (n_31_34), .A (n_30_37), .B (n_27_35), .C1 (n_28_36), .C2 (n_27_34) );
AOI211_X1 g_32_36 (.ZN (n_32_36), .A (n_29_35), .B (n_29_36), .C1 (n_26_37), .C2 (n_29_33) );
AOI211_X1 g_33_38 (.ZN (n_33_38), .A (n_31_34), .B (n_28_38), .C1 (n_27_35), .C2 (n_30_35) );
AOI211_X1 g_34_36 (.ZN (n_34_36), .A (n_32_36), .B (n_30_37), .C1 (n_29_36), .C2 (n_28_36) );
AOI211_X1 g_35_34 (.ZN (n_35_34), .A (n_33_38), .B (n_29_35), .C1 (n_28_38), .C2 (n_26_37) );
AOI211_X1 g_37_35 (.ZN (n_37_35), .A (n_34_36), .B (n_31_34), .C1 (n_30_37), .C2 (n_27_35) );
AOI211_X1 g_35_36 (.ZN (n_35_36), .A (n_35_34), .B (n_32_36), .C1 (n_29_35), .C2 (n_29_36) );
AOI211_X1 g_33_35 (.ZN (n_33_35), .A (n_37_35), .B (n_33_38), .C1 (n_31_34), .C2 (n_28_38) );
AOI211_X1 g_31_36 (.ZN (n_31_36), .A (n_35_36), .B (n_34_36), .C1 (n_32_36), .C2 (n_30_37) );
AOI211_X1 g_33_37 (.ZN (n_33_37), .A (n_33_35), .B (n_35_34), .C1 (n_33_38), .C2 (n_29_35) );
AOI211_X1 g_31_38 (.ZN (n_31_38), .A (n_31_36), .B (n_37_35), .C1 (n_34_36), .C2 (n_31_34) );
AOI211_X1 g_30_36 (.ZN (n_30_36), .A (n_33_37), .B (n_35_36), .C1 (n_35_34), .C2 (n_32_36) );
AOI211_X1 g_28_35 (.ZN (n_28_35), .A (n_31_38), .B (n_33_35), .C1 (n_37_35), .C2 (n_33_38) );
AOI211_X1 g_29_37 (.ZN (n_29_37), .A (n_30_36), .B (n_31_36), .C1 (n_35_36), .C2 (n_34_36) );
AOI211_X1 g_27_38 (.ZN (n_27_38), .A (n_28_35), .B (n_33_37), .C1 (n_33_35), .C2 (n_35_34) );
AOI211_X1 g_26_36 (.ZN (n_26_36), .A (n_29_37), .B (n_31_38), .C1 (n_31_36), .C2 (n_37_35) );
AOI211_X1 g_24_37 (.ZN (n_24_37), .A (n_27_38), .B (n_30_36), .C1 (n_33_37), .C2 (n_35_36) );
AOI211_X1 g_22_38 (.ZN (n_22_38), .A (n_26_36), .B (n_28_35), .C1 (n_31_38), .C2 (n_33_35) );
AOI211_X1 g_20_39 (.ZN (n_20_39), .A (n_24_37), .B (n_29_37), .C1 (n_30_36), .C2 (n_31_36) );
AOI211_X1 g_18_40 (.ZN (n_18_40), .A (n_22_38), .B (n_27_38), .C1 (n_28_35), .C2 (n_33_37) );
AOI211_X1 g_16_41 (.ZN (n_16_41), .A (n_20_39), .B (n_26_36), .C1 (n_29_37), .C2 (n_31_38) );
AOI211_X1 g_14_42 (.ZN (n_14_42), .A (n_18_40), .B (n_24_37), .C1 (n_27_38), .C2 (n_30_36) );
AOI211_X1 g_12_43 (.ZN (n_12_43), .A (n_16_41), .B (n_22_38), .C1 (n_26_36), .C2 (n_28_35) );
AOI211_X1 g_13_41 (.ZN (n_13_41), .A (n_14_42), .B (n_20_39), .C1 (n_24_37), .C2 (n_29_37) );
AOI211_X1 g_11_42 (.ZN (n_11_42), .A (n_12_43), .B (n_18_40), .C1 (n_22_38), .C2 (n_27_38) );
AOI211_X1 g_9_43 (.ZN (n_9_43), .A (n_13_41), .B (n_16_41), .C1 (n_20_39), .C2 (n_26_36) );
AOI211_X1 g_7_44 (.ZN (n_7_44), .A (n_11_42), .B (n_14_42), .C1 (n_18_40), .C2 (n_24_37) );
AOI211_X1 g_6_46 (.ZN (n_6_46), .A (n_9_43), .B (n_12_43), .C1 (n_16_41), .C2 (n_22_38) );
AOI211_X1 g_8_45 (.ZN (n_8_45), .A (n_7_44), .B (n_13_41), .C1 (n_14_42), .C2 (n_20_39) );
AOI211_X1 g_10_44 (.ZN (n_10_44), .A (n_6_46), .B (n_11_42), .C1 (n_12_43), .C2 (n_18_40) );
AOI211_X1 g_9_46 (.ZN (n_9_46), .A (n_8_45), .B (n_9_43), .C1 (n_13_41), .C2 (n_16_41) );
AOI211_X1 g_11_45 (.ZN (n_11_45), .A (n_10_44), .B (n_7_44), .C1 (n_11_42), .C2 (n_14_42) );
AOI211_X1 g_13_44 (.ZN (n_13_44), .A (n_9_46), .B (n_6_46), .C1 (n_9_43), .C2 (n_12_43) );
AOI211_X1 g_11_43 (.ZN (n_11_43), .A (n_11_45), .B (n_8_45), .C1 (n_7_44), .C2 (n_13_41) );
AOI211_X1 g_13_42 (.ZN (n_13_42), .A (n_13_44), .B (n_10_44), .C1 (n_6_46), .C2 (n_11_42) );
AOI211_X1 g_15_41 (.ZN (n_15_41), .A (n_11_43), .B (n_9_46), .C1 (n_8_45), .C2 (n_9_43) );
AOI211_X1 g_17_40 (.ZN (n_17_40), .A (n_13_42), .B (n_11_45), .C1 (n_10_44), .C2 (n_7_44) );
AOI211_X1 g_19_39 (.ZN (n_19_39), .A (n_15_41), .B (n_13_44), .C1 (n_9_46), .C2 (n_6_46) );
AOI211_X1 g_21_38 (.ZN (n_21_38), .A (n_17_40), .B (n_11_43), .C1 (n_11_45), .C2 (n_8_45) );
AOI211_X1 g_23_37 (.ZN (n_23_37), .A (n_19_39), .B (n_13_42), .C1 (n_13_44), .C2 (n_10_44) );
AOI211_X1 g_25_36 (.ZN (n_25_36), .A (n_21_38), .B (n_15_41), .C1 (n_11_43), .C2 (n_9_46) );
AOI211_X1 g_24_38 (.ZN (n_24_38), .A (n_23_37), .B (n_17_40), .C1 (n_13_42), .C2 (n_11_45) );
AOI211_X1 g_22_39 (.ZN (n_22_39), .A (n_25_36), .B (n_19_39), .C1 (n_15_41), .C2 (n_13_44) );
AOI211_X1 g_20_40 (.ZN (n_20_40), .A (n_24_38), .B (n_21_38), .C1 (n_17_40), .C2 (n_11_43) );
AOI211_X1 g_18_41 (.ZN (n_18_41), .A (n_22_39), .B (n_23_37), .C1 (n_19_39), .C2 (n_13_42) );
AOI211_X1 g_16_42 (.ZN (n_16_42), .A (n_20_40), .B (n_25_36), .C1 (n_21_38), .C2 (n_15_41) );
AOI211_X1 g_14_43 (.ZN (n_14_43), .A (n_18_41), .B (n_24_38), .C1 (n_23_37), .C2 (n_17_40) );
AOI211_X1 g_12_44 (.ZN (n_12_44), .A (n_16_42), .B (n_22_39), .C1 (n_25_36), .C2 (n_19_39) );
AOI211_X1 g_10_45 (.ZN (n_10_45), .A (n_14_43), .B (n_20_40), .C1 (n_24_38), .C2 (n_21_38) );
AOI211_X1 g_8_46 (.ZN (n_8_46), .A (n_12_44), .B (n_18_41), .C1 (n_22_39), .C2 (n_23_37) );
AOI211_X1 g_6_47 (.ZN (n_6_47), .A (n_10_45), .B (n_16_42), .C1 (n_20_40), .C2 (n_25_36) );
AOI211_X1 g_5_49 (.ZN (n_5_49), .A (n_8_46), .B (n_14_43), .C1 (n_18_41), .C2 (n_24_38) );
AOI211_X1 g_7_48 (.ZN (n_7_48), .A (n_6_47), .B (n_12_44), .C1 (n_16_42), .C2 (n_22_39) );
AOI211_X1 g_9_47 (.ZN (n_9_47), .A (n_5_49), .B (n_10_45), .C1 (n_14_43), .C2 (n_20_40) );
AOI211_X1 g_11_46 (.ZN (n_11_46), .A (n_7_48), .B (n_8_46), .C1 (n_12_44), .C2 (n_18_41) );
AOI211_X1 g_13_45 (.ZN (n_13_45), .A (n_9_47), .B (n_6_47), .C1 (n_10_45), .C2 (n_16_42) );
AOI211_X1 g_11_44 (.ZN (n_11_44), .A (n_11_46), .B (n_5_49), .C1 (n_8_46), .C2 (n_14_43) );
AOI211_X1 g_13_43 (.ZN (n_13_43), .A (n_13_45), .B (n_7_48), .C1 (n_6_47), .C2 (n_12_44) );
AOI211_X1 g_15_42 (.ZN (n_15_42), .A (n_11_44), .B (n_9_47), .C1 (n_5_49), .C2 (n_10_45) );
AOI211_X1 g_14_44 (.ZN (n_14_44), .A (n_13_43), .B (n_11_46), .C1 (n_7_48), .C2 (n_8_46) );
AOI211_X1 g_16_43 (.ZN (n_16_43), .A (n_15_42), .B (n_13_45), .C1 (n_9_47), .C2 (n_6_47) );
AOI211_X1 g_18_42 (.ZN (n_18_42), .A (n_14_44), .B (n_11_44), .C1 (n_11_46), .C2 (n_5_49) );
AOI211_X1 g_20_41 (.ZN (n_20_41), .A (n_16_43), .B (n_13_43), .C1 (n_13_45), .C2 (n_7_48) );
AOI211_X1 g_22_40 (.ZN (n_22_40), .A (n_18_42), .B (n_15_42), .C1 (n_11_44), .C2 (n_9_47) );
AOI211_X1 g_24_39 (.ZN (n_24_39), .A (n_20_41), .B (n_14_44), .C1 (n_13_43), .C2 (n_11_46) );
AOI211_X1 g_26_38 (.ZN (n_26_38), .A (n_22_40), .B (n_16_43), .C1 (n_15_42), .C2 (n_13_45) );
AOI211_X1 g_28_37 (.ZN (n_28_37), .A (n_24_39), .B (n_18_42), .C1 (n_14_44), .C2 (n_11_44) );
AOI211_X1 g_29_39 (.ZN (n_29_39), .A (n_26_38), .B (n_20_41), .C1 (n_16_43), .C2 (n_13_43) );
AOI211_X1 g_27_40 (.ZN (n_27_40), .A (n_28_37), .B (n_22_40), .C1 (n_18_42), .C2 (n_15_42) );
AOI211_X1 g_25_39 (.ZN (n_25_39), .A (n_29_39), .B (n_24_39), .C1 (n_20_41), .C2 (n_14_44) );
AOI211_X1 g_23_40 (.ZN (n_23_40), .A (n_27_40), .B (n_26_38), .C1 (n_22_40), .C2 (n_16_43) );
AOI211_X1 g_21_41 (.ZN (n_21_41), .A (n_25_39), .B (n_28_37), .C1 (n_24_39), .C2 (n_18_42) );
AOI211_X1 g_19_42 (.ZN (n_19_42), .A (n_23_40), .B (n_29_39), .C1 (n_26_38), .C2 (n_20_41) );
AOI211_X1 g_17_43 (.ZN (n_17_43), .A (n_21_41), .B (n_27_40), .C1 (n_28_37), .C2 (n_22_40) );
AOI211_X1 g_15_44 (.ZN (n_15_44), .A (n_19_42), .B (n_25_39), .C1 (n_29_39), .C2 (n_24_39) );
AOI211_X1 g_14_46 (.ZN (n_14_46), .A (n_17_43), .B (n_23_40), .C1 (n_27_40), .C2 (n_26_38) );
AOI211_X1 g_12_45 (.ZN (n_12_45), .A (n_15_44), .B (n_21_41), .C1 (n_25_39), .C2 (n_28_37) );
AOI211_X1 g_10_46 (.ZN (n_10_46), .A (n_14_46), .B (n_19_42), .C1 (n_23_40), .C2 (n_29_39) );
AOI211_X1 g_8_47 (.ZN (n_8_47), .A (n_12_45), .B (n_17_43), .C1 (n_21_41), .C2 (n_27_40) );
AOI211_X1 g_7_49 (.ZN (n_7_49), .A (n_10_46), .B (n_15_44), .C1 (n_19_42), .C2 (n_25_39) );
AOI211_X1 g_5_48 (.ZN (n_5_48), .A (n_8_47), .B (n_14_46), .C1 (n_17_43), .C2 (n_23_40) );
AOI211_X1 g_7_47 (.ZN (n_7_47), .A (n_7_49), .B (n_12_45), .C1 (n_15_44), .C2 (n_21_41) );
AOI211_X1 g_9_48 (.ZN (n_9_48), .A (n_5_48), .B (n_10_46), .C1 (n_14_46), .C2 (n_19_42) );
AOI211_X1 g_11_47 (.ZN (n_11_47), .A (n_7_47), .B (n_8_47), .C1 (n_12_45), .C2 (n_17_43) );
AOI211_X1 g_13_46 (.ZN (n_13_46), .A (n_9_48), .B (n_7_49), .C1 (n_10_46), .C2 (n_15_44) );
AOI211_X1 g_15_45 (.ZN (n_15_45), .A (n_11_47), .B (n_5_48), .C1 (n_8_47), .C2 (n_14_46) );
AOI211_X1 g_17_44 (.ZN (n_17_44), .A (n_13_46), .B (n_7_47), .C1 (n_7_49), .C2 (n_12_45) );
AOI211_X1 g_15_43 (.ZN (n_15_43), .A (n_15_45), .B (n_9_48), .C1 (n_5_48), .C2 (n_10_46) );
AOI211_X1 g_17_42 (.ZN (n_17_42), .A (n_17_44), .B (n_11_47), .C1 (n_7_47), .C2 (n_8_47) );
AOI211_X1 g_19_41 (.ZN (n_19_41), .A (n_15_43), .B (n_13_46), .C1 (n_9_48), .C2 (n_7_49) );
AOI211_X1 g_21_40 (.ZN (n_21_40), .A (n_17_42), .B (n_15_45), .C1 (n_11_47), .C2 (n_5_48) );
AOI211_X1 g_23_39 (.ZN (n_23_39), .A (n_19_41), .B (n_17_44), .C1 (n_13_46), .C2 (n_7_47) );
AOI211_X1 g_25_38 (.ZN (n_25_38), .A (n_21_40), .B (n_15_43), .C1 (n_15_45), .C2 (n_9_48) );
AOI211_X1 g_27_37 (.ZN (n_27_37), .A (n_23_39), .B (n_17_42), .C1 (n_17_44), .C2 (n_11_47) );
AOI211_X1 g_26_39 (.ZN (n_26_39), .A (n_25_38), .B (n_19_41), .C1 (n_15_43), .C2 (n_13_46) );
AOI211_X1 g_24_40 (.ZN (n_24_40), .A (n_27_37), .B (n_21_40), .C1 (n_17_42), .C2 (n_15_45) );
AOI211_X1 g_22_41 (.ZN (n_22_41), .A (n_26_39), .B (n_23_39), .C1 (n_19_41), .C2 (n_17_44) );
AOI211_X1 g_20_42 (.ZN (n_20_42), .A (n_24_40), .B (n_25_38), .C1 (n_21_40), .C2 (n_15_43) );
AOI211_X1 g_18_43 (.ZN (n_18_43), .A (n_22_41), .B (n_27_37), .C1 (n_23_39), .C2 (n_17_42) );
AOI211_X1 g_16_44 (.ZN (n_16_44), .A (n_20_42), .B (n_26_39), .C1 (n_25_38), .C2 (n_19_41) );
AOI211_X1 g_14_45 (.ZN (n_14_45), .A (n_18_43), .B (n_24_40), .C1 (n_27_37), .C2 (n_21_40) );
AOI211_X1 g_12_46 (.ZN (n_12_46), .A (n_16_44), .B (n_22_41), .C1 (n_26_39), .C2 (n_23_39) );
AOI211_X1 g_10_47 (.ZN (n_10_47), .A (n_14_45), .B (n_20_42), .C1 (n_24_40), .C2 (n_25_38) );
AOI211_X1 g_8_48 (.ZN (n_8_48), .A (n_12_46), .B (n_18_43), .C1 (n_22_41), .C2 (n_27_37) );
AOI211_X1 g_6_49 (.ZN (n_6_49), .A (n_10_47), .B (n_16_44), .C1 (n_20_42), .C2 (n_26_39) );
AOI211_X1 g_4_50 (.ZN (n_4_50), .A (n_8_48), .B (n_14_45), .C1 (n_18_43), .C2 (n_24_40) );
AOI211_X1 g_3_52 (.ZN (n_3_52), .A (n_6_49), .B (n_12_46), .C1 (n_16_44), .C2 (n_22_41) );
AOI211_X1 g_5_51 (.ZN (n_5_51), .A (n_4_50), .B (n_10_47), .C1 (n_14_45), .C2 (n_20_42) );
AOI211_X1 g_7_50 (.ZN (n_7_50), .A (n_3_52), .B (n_8_48), .C1 (n_12_46), .C2 (n_18_43) );
AOI211_X1 g_9_49 (.ZN (n_9_49), .A (n_5_51), .B (n_6_49), .C1 (n_10_47), .C2 (n_16_44) );
AOI211_X1 g_11_48 (.ZN (n_11_48), .A (n_7_50), .B (n_4_50), .C1 (n_8_48), .C2 (n_14_45) );
AOI211_X1 g_13_47 (.ZN (n_13_47), .A (n_9_49), .B (n_3_52), .C1 (n_6_49), .C2 (n_12_46) );
AOI211_X1 g_15_46 (.ZN (n_15_46), .A (n_11_48), .B (n_5_51), .C1 (n_4_50), .C2 (n_10_47) );
AOI211_X1 g_17_45 (.ZN (n_17_45), .A (n_13_47), .B (n_7_50), .C1 (n_3_52), .C2 (n_8_48) );
AOI211_X1 g_19_44 (.ZN (n_19_44), .A (n_15_46), .B (n_9_49), .C1 (n_5_51), .C2 (n_6_49) );
AOI211_X1 g_21_43 (.ZN (n_21_43), .A (n_17_45), .B (n_11_48), .C1 (n_7_50), .C2 (n_4_50) );
AOI211_X1 g_23_42 (.ZN (n_23_42), .A (n_19_44), .B (n_13_47), .C1 (n_9_49), .C2 (n_3_52) );
AOI211_X1 g_25_41 (.ZN (n_25_41), .A (n_21_43), .B (n_15_46), .C1 (n_11_48), .C2 (n_5_51) );
AOI211_X1 g_24_43 (.ZN (n_24_43), .A (n_23_42), .B (n_17_45), .C1 (n_13_47), .C2 (n_7_50) );
AOI211_X1 g_23_41 (.ZN (n_23_41), .A (n_25_41), .B (n_19_44), .C1 (n_15_46), .C2 (n_9_49) );
AOI211_X1 g_25_40 (.ZN (n_25_40), .A (n_24_43), .B (n_21_43), .C1 (n_17_45), .C2 (n_11_48) );
AOI211_X1 g_27_39 (.ZN (n_27_39), .A (n_23_41), .B (n_23_42), .C1 (n_19_44), .C2 (n_13_47) );
AOI211_X1 g_29_38 (.ZN (n_29_38), .A (n_25_40), .B (n_25_41), .C1 (n_21_43), .C2 (n_15_46) );
AOI211_X1 g_28_40 (.ZN (n_28_40), .A (n_27_39), .B (n_24_43), .C1 (n_23_42), .C2 (n_17_45) );
AOI211_X1 g_30_39 (.ZN (n_30_39), .A (n_29_38), .B (n_23_41), .C1 (n_25_41), .C2 (n_19_44) );
AOI211_X1 g_32_38 (.ZN (n_32_38), .A (n_28_40), .B (n_25_40), .C1 (n_24_43), .C2 (n_21_43) );
AOI211_X1 g_34_37 (.ZN (n_34_37), .A (n_30_39), .B (n_27_39), .C1 (n_23_41), .C2 (n_23_42) );
AOI211_X1 g_36_36 (.ZN (n_36_36), .A (n_32_38), .B (n_29_38), .C1 (n_25_40), .C2 (n_25_41) );
AOI211_X1 g_38_35 (.ZN (n_38_35), .A (n_34_37), .B (n_28_40), .C1 (n_27_39), .C2 (n_24_43) );
AOI211_X1 g_37_37 (.ZN (n_37_37), .A (n_36_36), .B (n_30_39), .C1 (n_29_38), .C2 (n_23_41) );
AOI211_X1 g_35_38 (.ZN (n_35_38), .A (n_38_35), .B (n_32_38), .C1 (n_28_40), .C2 (n_25_40) );
AOI211_X1 g_33_39 (.ZN (n_33_39), .A (n_37_37), .B (n_34_37), .C1 (n_30_39), .C2 (n_27_39) );
AOI211_X1 g_32_37 (.ZN (n_32_37), .A (n_35_38), .B (n_36_36), .C1 (n_32_38), .C2 (n_29_38) );
AOI211_X1 g_30_38 (.ZN (n_30_38), .A (n_33_39), .B (n_38_35), .C1 (n_34_37), .C2 (n_28_40) );
AOI211_X1 g_28_39 (.ZN (n_28_39), .A (n_32_37), .B (n_37_37), .C1 (n_36_36), .C2 (n_30_39) );
AOI211_X1 g_26_40 (.ZN (n_26_40), .A (n_30_38), .B (n_35_38), .C1 (n_38_35), .C2 (n_32_38) );
AOI211_X1 g_24_41 (.ZN (n_24_41), .A (n_28_39), .B (n_33_39), .C1 (n_37_37), .C2 (n_34_37) );
AOI211_X1 g_22_42 (.ZN (n_22_42), .A (n_26_40), .B (n_32_37), .C1 (n_35_38), .C2 (n_36_36) );
AOI211_X1 g_20_43 (.ZN (n_20_43), .A (n_24_41), .B (n_30_38), .C1 (n_33_39), .C2 (n_38_35) );
AOI211_X1 g_18_44 (.ZN (n_18_44), .A (n_22_42), .B (n_28_39), .C1 (n_32_37), .C2 (n_37_37) );
AOI211_X1 g_16_45 (.ZN (n_16_45), .A (n_20_43), .B (n_26_40), .C1 (n_30_38), .C2 (n_35_38) );
AOI211_X1 g_15_47 (.ZN (n_15_47), .A (n_18_44), .B (n_24_41), .C1 (n_28_39), .C2 (n_33_39) );
AOI211_X1 g_17_46 (.ZN (n_17_46), .A (n_16_45), .B (n_22_42), .C1 (n_26_40), .C2 (n_32_37) );
AOI211_X1 g_19_45 (.ZN (n_19_45), .A (n_15_47), .B (n_20_43), .C1 (n_24_41), .C2 (n_30_38) );
AOI211_X1 g_21_44 (.ZN (n_21_44), .A (n_17_46), .B (n_18_44), .C1 (n_22_42), .C2 (n_28_39) );
AOI211_X1 g_19_43 (.ZN (n_19_43), .A (n_19_45), .B (n_16_45), .C1 (n_20_43), .C2 (n_26_40) );
AOI211_X1 g_21_42 (.ZN (n_21_42), .A (n_21_44), .B (n_15_47), .C1 (n_18_44), .C2 (n_24_41) );
AOI211_X1 g_22_44 (.ZN (n_22_44), .A (n_19_43), .B (n_17_46), .C1 (n_16_45), .C2 (n_22_42) );
AOI211_X1 g_20_45 (.ZN (n_20_45), .A (n_21_42), .B (n_19_45), .C1 (n_15_47), .C2 (n_20_43) );
AOI211_X1 g_18_46 (.ZN (n_18_46), .A (n_22_44), .B (n_21_44), .C1 (n_17_46), .C2 (n_18_44) );
AOI211_X1 g_16_47 (.ZN (n_16_47), .A (n_20_45), .B (n_19_43), .C1 (n_19_45), .C2 (n_16_45) );
AOI211_X1 g_14_48 (.ZN (n_14_48), .A (n_18_46), .B (n_21_42), .C1 (n_21_44), .C2 (n_15_47) );
AOI211_X1 g_12_47 (.ZN (n_12_47), .A (n_16_47), .B (n_22_44), .C1 (n_19_43), .C2 (n_17_46) );
AOI211_X1 g_10_48 (.ZN (n_10_48), .A (n_14_48), .B (n_20_45), .C1 (n_21_42), .C2 (n_19_45) );
AOI211_X1 g_8_49 (.ZN (n_8_49), .A (n_12_47), .B (n_18_46), .C1 (n_22_44), .C2 (n_21_44) );
AOI211_X1 g_6_50 (.ZN (n_6_50), .A (n_10_48), .B (n_16_47), .C1 (n_20_45), .C2 (n_19_43) );
AOI211_X1 g_4_51 (.ZN (n_4_51), .A (n_8_49), .B (n_14_48), .C1 (n_18_46), .C2 (n_21_42) );
AOI211_X1 g_3_53 (.ZN (n_3_53), .A (n_6_50), .B (n_12_47), .C1 (n_16_47), .C2 (n_22_44) );
AOI211_X1 g_5_52 (.ZN (n_5_52), .A (n_4_51), .B (n_10_48), .C1 (n_14_48), .C2 (n_20_45) );
AOI211_X1 g_7_51 (.ZN (n_7_51), .A (n_3_53), .B (n_8_49), .C1 (n_12_47), .C2 (n_18_46) );
AOI211_X1 g_9_50 (.ZN (n_9_50), .A (n_5_52), .B (n_6_50), .C1 (n_10_48), .C2 (n_16_47) );
AOI211_X1 g_11_49 (.ZN (n_11_49), .A (n_7_51), .B (n_4_51), .C1 (n_8_49), .C2 (n_14_48) );
AOI211_X1 g_13_48 (.ZN (n_13_48), .A (n_9_50), .B (n_3_53), .C1 (n_6_50), .C2 (n_12_47) );
AOI211_X1 g_12_50 (.ZN (n_12_50), .A (n_11_49), .B (n_5_52), .C1 (n_4_51), .C2 (n_10_48) );
AOI211_X1 g_10_49 (.ZN (n_10_49), .A (n_13_48), .B (n_7_51), .C1 (n_3_53), .C2 (n_8_49) );
AOI211_X1 g_12_48 (.ZN (n_12_48), .A (n_12_50), .B (n_9_50), .C1 (n_5_52), .C2 (n_6_50) );
AOI211_X1 g_14_47 (.ZN (n_14_47), .A (n_10_49), .B (n_11_49), .C1 (n_7_51), .C2 (n_4_51) );
AOI211_X1 g_16_46 (.ZN (n_16_46), .A (n_12_48), .B (n_13_48), .C1 (n_9_50), .C2 (n_3_53) );
AOI211_X1 g_18_45 (.ZN (n_18_45), .A (n_14_47), .B (n_12_50), .C1 (n_11_49), .C2 (n_5_52) );
AOI211_X1 g_20_44 (.ZN (n_20_44), .A (n_16_46), .B (n_10_49), .C1 (n_13_48), .C2 (n_7_51) );
AOI211_X1 g_22_43 (.ZN (n_22_43), .A (n_18_45), .B (n_12_48), .C1 (n_12_50), .C2 (n_9_50) );
AOI211_X1 g_24_42 (.ZN (n_24_42), .A (n_20_44), .B (n_14_47), .C1 (n_10_49), .C2 (n_11_49) );
AOI211_X1 g_26_41 (.ZN (n_26_41), .A (n_22_43), .B (n_16_46), .C1 (n_12_48), .C2 (n_13_48) );
AOI211_X1 g_25_43 (.ZN (n_25_43), .A (n_24_42), .B (n_18_45), .C1 (n_14_47), .C2 (n_12_50) );
AOI211_X1 g_27_42 (.ZN (n_27_42), .A (n_26_41), .B (n_20_44), .C1 (n_16_46), .C2 (n_10_49) );
AOI211_X1 g_29_41 (.ZN (n_29_41), .A (n_25_43), .B (n_22_43), .C1 (n_18_45), .C2 (n_12_48) );
AOI211_X1 g_31_40 (.ZN (n_31_40), .A (n_27_42), .B (n_24_42), .C1 (n_20_44), .C2 (n_14_47) );
AOI211_X1 g_30_42 (.ZN (n_30_42), .A (n_29_41), .B (n_26_41), .C1 (n_22_43), .C2 (n_16_46) );
AOI211_X1 g_29_40 (.ZN (n_29_40), .A (n_31_40), .B (n_25_43), .C1 (n_24_42), .C2 (n_18_45) );
AOI211_X1 g_31_39 (.ZN (n_31_39), .A (n_30_42), .B (n_27_42), .C1 (n_26_41), .C2 (n_20_44) );
AOI211_X1 g_30_41 (.ZN (n_30_41), .A (n_29_40), .B (n_29_41), .C1 (n_25_43), .C2 (n_22_43) );
AOI211_X1 g_32_40 (.ZN (n_32_40), .A (n_31_39), .B (n_31_40), .C1 (n_27_42), .C2 (n_24_42) );
AOI211_X1 g_34_39 (.ZN (n_34_39), .A (n_30_41), .B (n_30_42), .C1 (n_29_41), .C2 (n_26_41) );
AOI211_X1 g_36_38 (.ZN (n_36_38), .A (n_32_40), .B (n_29_40), .C1 (n_31_40), .C2 (n_25_43) );
AOI211_X1 g_38_37 (.ZN (n_38_37), .A (n_34_39), .B (n_31_39), .C1 (n_30_42), .C2 (n_27_42) );
AOI211_X1 g_40_36 (.ZN (n_40_36), .A (n_36_38), .B (n_30_41), .C1 (n_29_40), .C2 (n_29_41) );
AOI211_X1 g_42_35 (.ZN (n_42_35), .A (n_38_37), .B (n_32_40), .C1 (n_31_39), .C2 (n_31_40) );
AOI211_X1 g_44_34 (.ZN (n_44_34), .A (n_40_36), .B (n_34_39), .C1 (n_30_41), .C2 (n_30_42) );
AOI211_X1 g_43_36 (.ZN (n_43_36), .A (n_42_35), .B (n_36_38), .C1 (n_32_40), .C2 (n_29_40) );
AOI211_X1 g_45_35 (.ZN (n_45_35), .A (n_44_34), .B (n_38_37), .C1 (n_34_39), .C2 (n_31_39) );
AOI211_X1 g_47_34 (.ZN (n_47_34), .A (n_43_36), .B (n_40_36), .C1 (n_36_38), .C2 (n_30_41) );
AOI211_X1 g_49_33 (.ZN (n_49_33), .A (n_45_35), .B (n_42_35), .C1 (n_38_37), .C2 (n_32_40) );
AOI211_X1 g_48_35 (.ZN (n_48_35), .A (n_47_34), .B (n_44_34), .C1 (n_40_36), .C2 (n_34_39) );
AOI211_X1 g_47_33 (.ZN (n_47_33), .A (n_49_33), .B (n_43_36), .C1 (n_42_35), .C2 (n_36_38) );
AOI211_X1 g_49_32 (.ZN (n_49_32), .A (n_48_35), .B (n_45_35), .C1 (n_44_34), .C2 (n_38_37) );
AOI211_X1 g_51_31 (.ZN (n_51_31), .A (n_47_33), .B (n_47_34), .C1 (n_43_36), .C2 (n_40_36) );
AOI211_X1 g_53_30 (.ZN (n_53_30), .A (n_49_32), .B (n_49_33), .C1 (n_45_35), .C2 (n_42_35) );
AOI211_X1 g_55_29 (.ZN (n_55_29), .A (n_51_31), .B (n_48_35), .C1 (n_47_34), .C2 (n_44_34) );
AOI211_X1 g_57_28 (.ZN (n_57_28), .A (n_53_30), .B (n_47_33), .C1 (n_49_33), .C2 (n_43_36) );
AOI211_X1 g_56_30 (.ZN (n_56_30), .A (n_55_29), .B (n_49_32), .C1 (n_48_35), .C2 (n_45_35) );
AOI211_X1 g_58_29 (.ZN (n_58_29), .A (n_57_28), .B (n_51_31), .C1 (n_47_33), .C2 (n_47_34) );
AOI211_X1 g_60_28 (.ZN (n_60_28), .A (n_56_30), .B (n_53_30), .C1 (n_49_32), .C2 (n_49_33) );
AOI211_X1 g_58_27 (.ZN (n_58_27), .A (n_58_29), .B (n_55_29), .C1 (n_51_31), .C2 (n_48_35) );
AOI211_X1 g_60_26 (.ZN (n_60_26), .A (n_60_28), .B (n_57_28), .C1 (n_53_30), .C2 (n_47_33) );
AOI211_X1 g_62_25 (.ZN (n_62_25), .A (n_58_27), .B (n_56_30), .C1 (n_55_29), .C2 (n_49_32) );
AOI211_X1 g_64_24 (.ZN (n_64_24), .A (n_60_26), .B (n_58_29), .C1 (n_57_28), .C2 (n_51_31) );
AOI211_X1 g_63_26 (.ZN (n_63_26), .A (n_62_25), .B (n_60_28), .C1 (n_56_30), .C2 (n_53_30) );
AOI211_X1 g_65_25 (.ZN (n_65_25), .A (n_64_24), .B (n_58_27), .C1 (n_58_29), .C2 (n_55_29) );
AOI211_X1 g_67_24 (.ZN (n_67_24), .A (n_63_26), .B (n_60_26), .C1 (n_60_28), .C2 (n_57_28) );
AOI211_X1 g_69_23 (.ZN (n_69_23), .A (n_65_25), .B (n_62_25), .C1 (n_58_27), .C2 (n_56_30) );
AOI211_X1 g_71_22 (.ZN (n_71_22), .A (n_67_24), .B (n_64_24), .C1 (n_60_26), .C2 (n_58_29) );
AOI211_X1 g_73_21 (.ZN (n_73_21), .A (n_69_23), .B (n_63_26), .C1 (n_62_25), .C2 (n_60_28) );
AOI211_X1 g_75_20 (.ZN (n_75_20), .A (n_71_22), .B (n_65_25), .C1 (n_64_24), .C2 (n_58_27) );
AOI211_X1 g_77_19 (.ZN (n_77_19), .A (n_73_21), .B (n_67_24), .C1 (n_63_26), .C2 (n_60_26) );
AOI211_X1 g_79_18 (.ZN (n_79_18), .A (n_75_20), .B (n_69_23), .C1 (n_65_25), .C2 (n_62_25) );
AOI211_X1 g_81_17 (.ZN (n_81_17), .A (n_77_19), .B (n_71_22), .C1 (n_67_24), .C2 (n_64_24) );
AOI211_X1 g_83_16 (.ZN (n_83_16), .A (n_79_18), .B (n_73_21), .C1 (n_69_23), .C2 (n_63_26) );
AOI211_X1 g_82_18 (.ZN (n_82_18), .A (n_81_17), .B (n_75_20), .C1 (n_71_22), .C2 (n_65_25) );
AOI211_X1 g_80_19 (.ZN (n_80_19), .A (n_83_16), .B (n_77_19), .C1 (n_73_21), .C2 (n_67_24) );
AOI211_X1 g_78_20 (.ZN (n_78_20), .A (n_82_18), .B (n_79_18), .C1 (n_75_20), .C2 (n_69_23) );
AOI211_X1 g_76_21 (.ZN (n_76_21), .A (n_80_19), .B (n_81_17), .C1 (n_77_19), .C2 (n_71_22) );
AOI211_X1 g_74_22 (.ZN (n_74_22), .A (n_78_20), .B (n_83_16), .C1 (n_79_18), .C2 (n_73_21) );
AOI211_X1 g_73_20 (.ZN (n_73_20), .A (n_76_21), .B (n_82_18), .C1 (n_81_17), .C2 (n_75_20) );
AOI211_X1 g_71_21 (.ZN (n_71_21), .A (n_74_22), .B (n_80_19), .C1 (n_83_16), .C2 (n_77_19) );
AOI211_X1 g_69_22 (.ZN (n_69_22), .A (n_73_20), .B (n_78_20), .C1 (n_82_18), .C2 (n_79_18) );
AOI211_X1 g_68_24 (.ZN (n_68_24), .A (n_71_21), .B (n_76_21), .C1 (n_80_19), .C2 (n_81_17) );
AOI211_X1 g_70_23 (.ZN (n_70_23), .A (n_69_22), .B (n_74_22), .C1 (n_78_20), .C2 (n_83_16) );
AOI211_X1 g_72_22 (.ZN (n_72_22), .A (n_68_24), .B (n_73_20), .C1 (n_76_21), .C2 (n_82_18) );
AOI211_X1 g_74_21 (.ZN (n_74_21), .A (n_70_23), .B (n_71_21), .C1 (n_74_22), .C2 (n_80_19) );
AOI211_X1 g_76_20 (.ZN (n_76_20), .A (n_72_22), .B (n_69_22), .C1 (n_73_20), .C2 (n_78_20) );
AOI211_X1 g_78_19 (.ZN (n_78_19), .A (n_74_21), .B (n_68_24), .C1 (n_71_21), .C2 (n_76_21) );
AOI211_X1 g_80_18 (.ZN (n_80_18), .A (n_76_20), .B (n_70_23), .C1 (n_69_22), .C2 (n_74_22) );
AOI211_X1 g_79_20 (.ZN (n_79_20), .A (n_78_19), .B (n_72_22), .C1 (n_68_24), .C2 (n_73_20) );
AOI211_X1 g_81_19 (.ZN (n_81_19), .A (n_80_18), .B (n_74_21), .C1 (n_70_23), .C2 (n_71_21) );
AOI211_X1 g_83_18 (.ZN (n_83_18), .A (n_79_20), .B (n_76_20), .C1 (n_72_22), .C2 (n_69_22) );
AOI211_X1 g_85_17 (.ZN (n_85_17), .A (n_81_19), .B (n_78_19), .C1 (n_74_21), .C2 (n_68_24) );
AOI211_X1 g_87_16 (.ZN (n_87_16), .A (n_83_18), .B (n_80_18), .C1 (n_76_20), .C2 (n_70_23) );
AOI211_X1 g_86_18 (.ZN (n_86_18), .A (n_85_17), .B (n_79_20), .C1 (n_78_19), .C2 (n_72_22) );
AOI211_X1 g_84_19 (.ZN (n_84_19), .A (n_87_16), .B (n_81_19), .C1 (n_80_18), .C2 (n_74_21) );
AOI211_X1 g_82_20 (.ZN (n_82_20), .A (n_86_18), .B (n_83_18), .C1 (n_79_20), .C2 (n_76_20) );
AOI211_X1 g_80_21 (.ZN (n_80_21), .A (n_84_19), .B (n_85_17), .C1 (n_81_19), .C2 (n_78_19) );
AOI211_X1 g_79_19 (.ZN (n_79_19), .A (n_82_20), .B (n_87_16), .C1 (n_83_18), .C2 (n_80_18) );
AOI211_X1 g_77_20 (.ZN (n_77_20), .A (n_80_21), .B (n_86_18), .C1 (n_85_17), .C2 (n_79_20) );
AOI211_X1 g_75_21 (.ZN (n_75_21), .A (n_79_19), .B (n_84_19), .C1 (n_87_16), .C2 (n_81_19) );
AOI211_X1 g_73_22 (.ZN (n_73_22), .A (n_77_20), .B (n_82_20), .C1 (n_86_18), .C2 (n_83_18) );
AOI211_X1 g_71_23 (.ZN (n_71_23), .A (n_75_21), .B (n_80_21), .C1 (n_84_19), .C2 (n_85_17) );
AOI211_X1 g_69_24 (.ZN (n_69_24), .A (n_73_22), .B (n_79_19), .C1 (n_82_20), .C2 (n_87_16) );
AOI211_X1 g_67_25 (.ZN (n_67_25), .A (n_71_23), .B (n_77_20), .C1 (n_80_21), .C2 (n_86_18) );
AOI211_X1 g_65_26 (.ZN (n_65_26), .A (n_69_24), .B (n_75_21), .C1 (n_79_19), .C2 (n_84_19) );
AOI211_X1 g_63_27 (.ZN (n_63_27), .A (n_67_25), .B (n_73_22), .C1 (n_77_20), .C2 (n_82_20) );
AOI211_X1 g_61_28 (.ZN (n_61_28), .A (n_65_26), .B (n_71_23), .C1 (n_75_21), .C2 (n_80_21) );
AOI211_X1 g_59_29 (.ZN (n_59_29), .A (n_63_27), .B (n_69_24), .C1 (n_73_22), .C2 (n_79_19) );
AOI211_X1 g_57_30 (.ZN (n_57_30), .A (n_61_28), .B (n_67_25), .C1 (n_71_23), .C2 (n_77_20) );
AOI211_X1 g_55_31 (.ZN (n_55_31), .A (n_59_29), .B (n_65_26), .C1 (n_69_24), .C2 (n_75_21) );
AOI211_X1 g_53_32 (.ZN (n_53_32), .A (n_57_30), .B (n_63_27), .C1 (n_67_25), .C2 (n_73_22) );
AOI211_X1 g_51_33 (.ZN (n_51_33), .A (n_55_31), .B (n_61_28), .C1 (n_65_26), .C2 (n_71_23) );
AOI211_X1 g_49_34 (.ZN (n_49_34), .A (n_53_32), .B (n_59_29), .C1 (n_63_27), .C2 (n_69_24) );
AOI211_X1 g_47_35 (.ZN (n_47_35), .A (n_51_33), .B (n_57_30), .C1 (n_61_28), .C2 (n_67_25) );
AOI211_X1 g_45_36 (.ZN (n_45_36), .A (n_49_34), .B (n_55_31), .C1 (n_59_29), .C2 (n_65_26) );
AOI211_X1 g_43_37 (.ZN (n_43_37), .A (n_47_35), .B (n_53_32), .C1 (n_57_30), .C2 (n_63_27) );
AOI211_X1 g_44_35 (.ZN (n_44_35), .A (n_45_36), .B (n_51_33), .C1 (n_55_31), .C2 (n_61_28) );
AOI211_X1 g_46_36 (.ZN (n_46_36), .A (n_43_37), .B (n_49_34), .C1 (n_53_32), .C2 (n_59_29) );
AOI211_X1 g_44_37 (.ZN (n_44_37), .A (n_44_35), .B (n_47_35), .C1 (n_51_33), .C2 (n_57_30) );
AOI211_X1 g_42_36 (.ZN (n_42_36), .A (n_46_36), .B (n_45_36), .C1 (n_49_34), .C2 (n_55_31) );
AOI211_X1 g_40_35 (.ZN (n_40_35), .A (n_44_37), .B (n_43_37), .C1 (n_47_35), .C2 (n_53_32) );
AOI211_X1 g_38_36 (.ZN (n_38_36), .A (n_42_36), .B (n_44_35), .C1 (n_45_36), .C2 (n_51_33) );
AOI211_X1 g_36_37 (.ZN (n_36_37), .A (n_40_35), .B (n_46_36), .C1 (n_43_37), .C2 (n_49_34) );
AOI211_X1 g_34_38 (.ZN (n_34_38), .A (n_38_36), .B (n_44_37), .C1 (n_44_35), .C2 (n_47_35) );
AOI211_X1 g_32_39 (.ZN (n_32_39), .A (n_36_37), .B (n_42_36), .C1 (n_46_36), .C2 (n_45_36) );
AOI211_X1 g_30_40 (.ZN (n_30_40), .A (n_34_38), .B (n_40_35), .C1 (n_44_37), .C2 (n_43_37) );
AOI211_X1 g_28_41 (.ZN (n_28_41), .A (n_32_39), .B (n_38_36), .C1 (n_42_36), .C2 (n_44_35) );
AOI211_X1 g_26_42 (.ZN (n_26_42), .A (n_30_40), .B (n_36_37), .C1 (n_40_35), .C2 (n_46_36) );
AOI211_X1 g_28_43 (.ZN (n_28_43), .A (n_28_41), .B (n_34_38), .C1 (n_38_36), .C2 (n_44_37) );
AOI211_X1 g_27_41 (.ZN (n_27_41), .A (n_26_42), .B (n_32_39), .C1 (n_36_37), .C2 (n_42_36) );
AOI211_X1 g_25_42 (.ZN (n_25_42), .A (n_28_43), .B (n_30_40), .C1 (n_34_38), .C2 (n_40_35) );
AOI211_X1 g_23_43 (.ZN (n_23_43), .A (n_27_41), .B (n_28_41), .C1 (n_32_39), .C2 (n_38_36) );
AOI211_X1 g_22_45 (.ZN (n_22_45), .A (n_25_42), .B (n_26_42), .C1 (n_30_40), .C2 (n_36_37) );
AOI211_X1 g_24_44 (.ZN (n_24_44), .A (n_23_43), .B (n_28_43), .C1 (n_28_41), .C2 (n_34_38) );
AOI211_X1 g_26_43 (.ZN (n_26_43), .A (n_22_45), .B (n_27_41), .C1 (n_26_42), .C2 (n_32_39) );
AOI211_X1 g_28_42 (.ZN (n_28_42), .A (n_24_44), .B (n_25_42), .C1 (n_28_43), .C2 (n_30_40) );
AOI211_X1 g_27_44 (.ZN (n_27_44), .A (n_26_43), .B (n_23_43), .C1 (n_27_41), .C2 (n_28_41) );
AOI211_X1 g_29_43 (.ZN (n_29_43), .A (n_28_42), .B (n_22_45), .C1 (n_25_42), .C2 (n_26_42) );
AOI211_X1 g_31_42 (.ZN (n_31_42), .A (n_27_44), .B (n_24_44), .C1 (n_23_43), .C2 (n_28_43) );
AOI211_X1 g_33_41 (.ZN (n_33_41), .A (n_29_43), .B (n_26_43), .C1 (n_22_45), .C2 (n_27_41) );
AOI211_X1 g_35_40 (.ZN (n_35_40), .A (n_31_42), .B (n_28_42), .C1 (n_24_44), .C2 (n_25_42) );
AOI211_X1 g_37_39 (.ZN (n_37_39), .A (n_33_41), .B (n_27_44), .C1 (n_26_43), .C2 (n_23_43) );
AOI211_X1 g_39_38 (.ZN (n_39_38), .A (n_35_40), .B (n_29_43), .C1 (n_28_42), .C2 (n_22_45) );
AOI211_X1 g_41_37 (.ZN (n_41_37), .A (n_37_39), .B (n_31_42), .C1 (n_27_44), .C2 (n_24_44) );
AOI211_X1 g_42_39 (.ZN (n_42_39), .A (n_39_38), .B (n_33_41), .C1 (n_29_43), .C2 (n_26_43) );
AOI211_X1 g_44_38 (.ZN (n_44_38), .A (n_41_37), .B (n_35_40), .C1 (n_31_42), .C2 (n_28_42) );
AOI211_X1 g_42_37 (.ZN (n_42_37), .A (n_42_39), .B (n_37_39), .C1 (n_33_41), .C2 (n_27_44) );
AOI211_X1 g_44_36 (.ZN (n_44_36), .A (n_44_38), .B (n_39_38), .C1 (n_35_40), .C2 (n_29_43) );
AOI211_X1 g_46_35 (.ZN (n_46_35), .A (n_42_37), .B (n_41_37), .C1 (n_37_39), .C2 (n_31_42) );
AOI211_X1 g_48_34 (.ZN (n_48_34), .A (n_44_36), .B (n_42_39), .C1 (n_39_38), .C2 (n_33_41) );
AOI211_X1 g_50_33 (.ZN (n_50_33), .A (n_46_35), .B (n_44_38), .C1 (n_41_37), .C2 (n_35_40) );
AOI211_X1 g_52_32 (.ZN (n_52_32), .A (n_48_34), .B (n_42_37), .C1 (n_42_39), .C2 (n_37_39) );
AOI211_X1 g_54_31 (.ZN (n_54_31), .A (n_50_33), .B (n_44_36), .C1 (n_44_38), .C2 (n_39_38) );
AOI211_X1 g_53_33 (.ZN (n_53_33), .A (n_52_32), .B (n_46_35), .C1 (n_42_37), .C2 (n_41_37) );
AOI211_X1 g_51_34 (.ZN (n_51_34), .A (n_54_31), .B (n_48_34), .C1 (n_44_36), .C2 (n_42_39) );
AOI211_X1 g_49_35 (.ZN (n_49_35), .A (n_53_33), .B (n_50_33), .C1 (n_46_35), .C2 (n_44_38) );
AOI211_X1 g_47_36 (.ZN (n_47_36), .A (n_51_34), .B (n_52_32), .C1 (n_48_34), .C2 (n_42_37) );
AOI211_X1 g_45_37 (.ZN (n_45_37), .A (n_49_35), .B (n_54_31), .C1 (n_50_33), .C2 (n_44_36) );
AOI211_X1 g_43_38 (.ZN (n_43_38), .A (n_47_36), .B (n_53_33), .C1 (n_52_32), .C2 (n_46_35) );
AOI211_X1 g_41_39 (.ZN (n_41_39), .A (n_45_37), .B (n_51_34), .C1 (n_54_31), .C2 (n_48_34) );
AOI211_X1 g_40_37 (.ZN (n_40_37), .A (n_43_38), .B (n_49_35), .C1 (n_53_33), .C2 (n_50_33) );
AOI211_X1 g_38_38 (.ZN (n_38_38), .A (n_41_39), .B (n_47_36), .C1 (n_51_34), .C2 (n_52_32) );
AOI211_X1 g_36_39 (.ZN (n_36_39), .A (n_40_37), .B (n_45_37), .C1 (n_49_35), .C2 (n_54_31) );
AOI211_X1 g_34_40 (.ZN (n_34_40), .A (n_38_38), .B (n_43_38), .C1 (n_47_36), .C2 (n_53_33) );
AOI211_X1 g_32_41 (.ZN (n_32_41), .A (n_36_39), .B (n_41_39), .C1 (n_45_37), .C2 (n_51_34) );
AOI211_X1 g_31_43 (.ZN (n_31_43), .A (n_34_40), .B (n_40_37), .C1 (n_43_38), .C2 (n_49_35) );
AOI211_X1 g_29_42 (.ZN (n_29_42), .A (n_32_41), .B (n_38_38), .C1 (n_41_39), .C2 (n_47_36) );
AOI211_X1 g_31_41 (.ZN (n_31_41), .A (n_31_43), .B (n_36_39), .C1 (n_40_37), .C2 (n_45_37) );
AOI211_X1 g_33_40 (.ZN (n_33_40), .A (n_29_42), .B (n_34_40), .C1 (n_38_38), .C2 (n_43_38) );
AOI211_X1 g_35_39 (.ZN (n_35_39), .A (n_31_41), .B (n_32_41), .C1 (n_36_39), .C2 (n_41_39) );
AOI211_X1 g_37_38 (.ZN (n_37_38), .A (n_33_40), .B (n_31_43), .C1 (n_34_40), .C2 (n_40_37) );
AOI211_X1 g_39_37 (.ZN (n_39_37), .A (n_35_39), .B (n_29_42), .C1 (n_32_41), .C2 (n_38_38) );
AOI211_X1 g_41_36 (.ZN (n_41_36), .A (n_37_38), .B (n_31_41), .C1 (n_31_43), .C2 (n_36_39) );
AOI211_X1 g_40_38 (.ZN (n_40_38), .A (n_39_37), .B (n_33_40), .C1 (n_29_42), .C2 (n_34_40) );
AOI211_X1 g_38_39 (.ZN (n_38_39), .A (n_41_36), .B (n_35_39), .C1 (n_31_41), .C2 (n_32_41) );
AOI211_X1 g_36_40 (.ZN (n_36_40), .A (n_40_38), .B (n_37_38), .C1 (n_33_40), .C2 (n_31_43) );
AOI211_X1 g_34_41 (.ZN (n_34_41), .A (n_38_39), .B (n_39_37), .C1 (n_35_39), .C2 (n_29_42) );
AOI211_X1 g_32_42 (.ZN (n_32_42), .A (n_36_40), .B (n_41_36), .C1 (n_37_38), .C2 (n_31_41) );
AOI211_X1 g_30_43 (.ZN (n_30_43), .A (n_34_41), .B (n_40_38), .C1 (n_39_37), .C2 (n_33_40) );
AOI211_X1 g_28_44 (.ZN (n_28_44), .A (n_32_42), .B (n_38_39), .C1 (n_41_36), .C2 (n_35_39) );
AOI211_X1 g_26_45 (.ZN (n_26_45), .A (n_30_43), .B (n_36_40), .C1 (n_40_38), .C2 (n_37_38) );
AOI211_X1 g_27_43 (.ZN (n_27_43), .A (n_28_44), .B (n_34_41), .C1 (n_38_39), .C2 (n_39_37) );
AOI211_X1 g_25_44 (.ZN (n_25_44), .A (n_26_45), .B (n_32_42), .C1 (n_36_40), .C2 (n_41_36) );
AOI211_X1 g_23_45 (.ZN (n_23_45), .A (n_27_43), .B (n_30_43), .C1 (n_34_41), .C2 (n_40_38) );
AOI211_X1 g_21_46 (.ZN (n_21_46), .A (n_25_44), .B (n_28_44), .C1 (n_32_42), .C2 (n_38_39) );
AOI211_X1 g_19_47 (.ZN (n_19_47), .A (n_23_45), .B (n_26_45), .C1 (n_30_43), .C2 (n_36_40) );
AOI211_X1 g_17_48 (.ZN (n_17_48), .A (n_21_46), .B (n_27_43), .C1 (n_28_44), .C2 (n_34_41) );
AOI211_X1 g_15_49 (.ZN (n_15_49), .A (n_19_47), .B (n_25_44), .C1 (n_26_45), .C2 (n_32_42) );
AOI211_X1 g_13_50 (.ZN (n_13_50), .A (n_17_48), .B (n_23_45), .C1 (n_27_43), .C2 (n_30_43) );
AOI211_X1 g_11_51 (.ZN (n_11_51), .A (n_15_49), .B (n_21_46), .C1 (n_25_44), .C2 (n_28_44) );
AOI211_X1 g_12_49 (.ZN (n_12_49), .A (n_13_50), .B (n_19_47), .C1 (n_23_45), .C2 (n_26_45) );
AOI211_X1 g_10_50 (.ZN (n_10_50), .A (n_11_51), .B (n_17_48), .C1 (n_21_46), .C2 (n_27_43) );
AOI211_X1 g_8_51 (.ZN (n_8_51), .A (n_12_49), .B (n_15_49), .C1 (n_19_47), .C2 (n_25_44) );
AOI211_X1 g_6_52 (.ZN (n_6_52), .A (n_10_50), .B (n_13_50), .C1 (n_17_48), .C2 (n_23_45) );
AOI211_X1 g_4_53 (.ZN (n_4_53), .A (n_8_51), .B (n_11_51), .C1 (n_15_49), .C2 (n_21_46) );
AOI211_X1 g_2_54 (.ZN (n_2_54), .A (n_6_52), .B (n_12_49), .C1 (n_13_50), .C2 (n_19_47) );
AOI211_X1 g_1_56 (.ZN (n_1_56), .A (n_4_53), .B (n_10_50), .C1 (n_11_51), .C2 (n_17_48) );
AOI211_X1 g_3_55 (.ZN (n_3_55), .A (n_2_54), .B (n_8_51), .C1 (n_12_49), .C2 (n_15_49) );
AOI211_X1 g_5_54 (.ZN (n_5_54), .A (n_1_56), .B (n_6_52), .C1 (n_10_50), .C2 (n_13_50) );
AOI211_X1 g_7_53 (.ZN (n_7_53), .A (n_3_55), .B (n_4_53), .C1 (n_8_51), .C2 (n_11_51) );
AOI211_X1 g_6_51 (.ZN (n_6_51), .A (n_5_54), .B (n_2_54), .C1 (n_6_52), .C2 (n_12_49) );
AOI211_X1 g_8_50 (.ZN (n_8_50), .A (n_7_53), .B (n_1_56), .C1 (n_4_53), .C2 (n_10_50) );
AOI211_X1 g_9_52 (.ZN (n_9_52), .A (n_6_51), .B (n_3_55), .C1 (n_2_54), .C2 (n_8_51) );
AOI211_X1 g_8_54 (.ZN (n_8_54), .A (n_8_50), .B (n_5_54), .C1 (n_1_56), .C2 (n_6_52) );
AOI211_X1 g_7_52 (.ZN (n_7_52), .A (n_9_52), .B (n_7_53), .C1 (n_3_55), .C2 (n_4_53) );
AOI211_X1 g_5_53 (.ZN (n_5_53), .A (n_8_54), .B (n_6_51), .C1 (n_5_54), .C2 (n_2_54) );
AOI211_X1 g_4_55 (.ZN (n_4_55), .A (n_7_52), .B (n_8_50), .C1 (n_7_53), .C2 (n_1_56) );
AOI211_X1 g_3_57 (.ZN (n_3_57), .A (n_5_53), .B (n_9_52), .C1 (n_6_51), .C2 (n_3_55) );
AOI211_X1 g_5_58 (.ZN (n_5_58), .A (n_4_55), .B (n_8_54), .C1 (n_8_50), .C2 (n_5_54) );
AOI211_X1 g_3_59 (.ZN (n_3_59), .A (n_3_57), .B (n_7_52), .C1 (n_9_52), .C2 (n_7_53) );
AOI211_X1 g_1_60 (.ZN (n_1_60), .A (n_5_58), .B (n_5_53), .C1 (n_8_54), .C2 (n_6_51) );
AOI211_X1 g_2_58 (.ZN (n_2_58), .A (n_3_59), .B (n_4_55), .C1 (n_7_52), .C2 (n_8_50) );
AOI211_X1 g_4_57 (.ZN (n_4_57), .A (n_1_60), .B (n_3_57), .C1 (n_5_53), .C2 (n_9_52) );
AOI211_X1 g_6_56 (.ZN (n_6_56), .A (n_2_58), .B (n_5_58), .C1 (n_4_55), .C2 (n_8_54) );
AOI211_X1 g_7_54 (.ZN (n_7_54), .A (n_4_57), .B (n_3_59), .C1 (n_3_57), .C2 (n_7_52) );
AOI211_X1 g_8_52 (.ZN (n_8_52), .A (n_6_56), .B (n_1_60), .C1 (n_5_58), .C2 (n_5_53) );
AOI211_X1 g_10_51 (.ZN (n_10_51), .A (n_7_54), .B (n_2_58), .C1 (n_3_59), .C2 (n_4_55) );
AOI211_X1 g_9_53 (.ZN (n_9_53), .A (n_8_52), .B (n_4_57), .C1 (n_1_60), .C2 (n_3_57) );
AOI211_X1 g_11_52 (.ZN (n_11_52), .A (n_10_51), .B (n_6_56), .C1 (n_2_58), .C2 (n_5_58) );
AOI211_X1 g_9_51 (.ZN (n_9_51), .A (n_9_53), .B (n_7_54), .C1 (n_4_57), .C2 (n_3_59) );
AOI211_X1 g_11_50 (.ZN (n_11_50), .A (n_11_52), .B (n_8_52), .C1 (n_6_56), .C2 (n_1_60) );
AOI211_X1 g_13_49 (.ZN (n_13_49), .A (n_9_51), .B (n_10_51), .C1 (n_7_54), .C2 (n_2_58) );
AOI211_X1 g_15_48 (.ZN (n_15_48), .A (n_11_50), .B (n_9_53), .C1 (n_8_52), .C2 (n_4_57) );
AOI211_X1 g_17_47 (.ZN (n_17_47), .A (n_13_49), .B (n_11_52), .C1 (n_10_51), .C2 (n_6_56) );
AOI211_X1 g_19_46 (.ZN (n_19_46), .A (n_15_48), .B (n_9_51), .C1 (n_9_53), .C2 (n_7_54) );
AOI211_X1 g_21_45 (.ZN (n_21_45), .A (n_17_47), .B (n_11_50), .C1 (n_11_52), .C2 (n_8_52) );
AOI211_X1 g_23_44 (.ZN (n_23_44), .A (n_19_46), .B (n_13_49), .C1 (n_9_51), .C2 (n_10_51) );
AOI211_X1 g_24_46 (.ZN (n_24_46), .A (n_21_45), .B (n_15_48), .C1 (n_11_50), .C2 (n_9_53) );
AOI211_X1 g_22_47 (.ZN (n_22_47), .A (n_23_44), .B (n_17_47), .C1 (n_13_49), .C2 (n_11_52) );
AOI211_X1 g_20_46 (.ZN (n_20_46), .A (n_24_46), .B (n_19_46), .C1 (n_15_48), .C2 (n_9_51) );
AOI211_X1 g_18_47 (.ZN (n_18_47), .A (n_22_47), .B (n_21_45), .C1 (n_17_47), .C2 (n_11_50) );
AOI211_X1 g_16_48 (.ZN (n_16_48), .A (n_20_46), .B (n_23_44), .C1 (n_19_46), .C2 (n_13_49) );
AOI211_X1 g_14_49 (.ZN (n_14_49), .A (n_18_47), .B (n_24_46), .C1 (n_21_45), .C2 (n_15_48) );
AOI211_X1 g_13_51 (.ZN (n_13_51), .A (n_16_48), .B (n_22_47), .C1 (n_23_44), .C2 (n_17_47) );
AOI211_X1 g_15_50 (.ZN (n_15_50), .A (n_14_49), .B (n_20_46), .C1 (n_24_46), .C2 (n_19_46) );
AOI211_X1 g_17_49 (.ZN (n_17_49), .A (n_13_51), .B (n_18_47), .C1 (n_22_47), .C2 (n_21_45) );
AOI211_X1 g_19_48 (.ZN (n_19_48), .A (n_15_50), .B (n_16_48), .C1 (n_20_46), .C2 (n_23_44) );
AOI211_X1 g_21_47 (.ZN (n_21_47), .A (n_17_49), .B (n_14_49), .C1 (n_18_47), .C2 (n_24_46) );
AOI211_X1 g_23_46 (.ZN (n_23_46), .A (n_19_48), .B (n_13_51), .C1 (n_16_48), .C2 (n_22_47) );
AOI211_X1 g_25_45 (.ZN (n_25_45), .A (n_21_47), .B (n_15_50), .C1 (n_14_49), .C2 (n_20_46) );
AOI211_X1 g_24_47 (.ZN (n_24_47), .A (n_23_46), .B (n_17_49), .C1 (n_13_51), .C2 (n_18_47) );
AOI211_X1 g_22_46 (.ZN (n_22_46), .A (n_25_45), .B (n_19_48), .C1 (n_15_50), .C2 (n_16_48) );
AOI211_X1 g_24_45 (.ZN (n_24_45), .A (n_24_47), .B (n_21_47), .C1 (n_17_49), .C2 (n_14_49) );
AOI211_X1 g_26_44 (.ZN (n_26_44), .A (n_22_46), .B (n_23_46), .C1 (n_19_48), .C2 (n_13_51) );
AOI211_X1 g_25_46 (.ZN (n_25_46), .A (n_24_45), .B (n_25_45), .C1 (n_21_47), .C2 (n_15_50) );
AOI211_X1 g_27_45 (.ZN (n_27_45), .A (n_26_44), .B (n_24_47), .C1 (n_23_46), .C2 (n_17_49) );
AOI211_X1 g_29_44 (.ZN (n_29_44), .A (n_25_46), .B (n_22_46), .C1 (n_25_45), .C2 (n_19_48) );
AOI211_X1 g_28_46 (.ZN (n_28_46), .A (n_27_45), .B (n_24_45), .C1 (n_24_47), .C2 (n_21_47) );
AOI211_X1 g_30_45 (.ZN (n_30_45), .A (n_29_44), .B (n_26_44), .C1 (n_22_46), .C2 (n_23_46) );
AOI211_X1 g_32_44 (.ZN (n_32_44), .A (n_28_46), .B (n_25_46), .C1 (n_24_45), .C2 (n_25_45) );
AOI211_X1 g_33_42 (.ZN (n_33_42), .A (n_30_45), .B (n_27_45), .C1 (n_26_44), .C2 (n_24_47) );
AOI211_X1 g_35_41 (.ZN (n_35_41), .A (n_32_44), .B (n_29_44), .C1 (n_25_46), .C2 (n_22_46) );
AOI211_X1 g_37_40 (.ZN (n_37_40), .A (n_33_42), .B (n_28_46), .C1 (n_27_45), .C2 (n_24_45) );
AOI211_X1 g_39_39 (.ZN (n_39_39), .A (n_35_41), .B (n_30_45), .C1 (n_29_44), .C2 (n_26_44) );
AOI211_X1 g_41_38 (.ZN (n_41_38), .A (n_37_40), .B (n_32_44), .C1 (n_28_46), .C2 (n_25_46) );
AOI211_X1 g_40_40 (.ZN (n_40_40), .A (n_39_39), .B (n_33_42), .C1 (n_30_45), .C2 (n_27_45) );
AOI211_X1 g_38_41 (.ZN (n_38_41), .A (n_41_38), .B (n_35_41), .C1 (n_32_44), .C2 (n_29_44) );
AOI211_X1 g_36_42 (.ZN (n_36_42), .A (n_40_40), .B (n_37_40), .C1 (n_33_42), .C2 (n_28_46) );
AOI211_X1 g_34_43 (.ZN (n_34_43), .A (n_38_41), .B (n_39_39), .C1 (n_35_41), .C2 (n_30_45) );
AOI211_X1 g_33_45 (.ZN (n_33_45), .A (n_36_42), .B (n_41_38), .C1 (n_37_40), .C2 (n_32_44) );
AOI211_X1 g_32_43 (.ZN (n_32_43), .A (n_34_43), .B (n_40_40), .C1 (n_39_39), .C2 (n_33_42) );
AOI211_X1 g_34_42 (.ZN (n_34_42), .A (n_33_45), .B (n_38_41), .C1 (n_41_38), .C2 (n_35_41) );
AOI211_X1 g_36_41 (.ZN (n_36_41), .A (n_32_43), .B (n_36_42), .C1 (n_40_40), .C2 (n_37_40) );
AOI211_X1 g_38_40 (.ZN (n_38_40), .A (n_34_42), .B (n_34_43), .C1 (n_38_41), .C2 (n_39_39) );
AOI211_X1 g_40_39 (.ZN (n_40_39), .A (n_36_41), .B (n_33_45), .C1 (n_36_42), .C2 (n_41_38) );
AOI211_X1 g_42_38 (.ZN (n_42_38), .A (n_38_40), .B (n_32_43), .C1 (n_34_43), .C2 (n_40_40) );
AOI211_X1 g_41_40 (.ZN (n_41_40), .A (n_40_39), .B (n_34_42), .C1 (n_33_45), .C2 (n_38_41) );
AOI211_X1 g_43_39 (.ZN (n_43_39), .A (n_42_38), .B (n_36_41), .C1 (n_32_43), .C2 (n_36_42) );
AOI211_X1 g_45_38 (.ZN (n_45_38), .A (n_41_40), .B (n_38_40), .C1 (n_34_42), .C2 (n_34_43) );
AOI211_X1 g_47_37 (.ZN (n_47_37), .A (n_43_39), .B (n_40_39), .C1 (n_36_41), .C2 (n_33_45) );
AOI211_X1 g_49_36 (.ZN (n_49_36), .A (n_45_38), .B (n_42_38), .C1 (n_38_40), .C2 (n_32_43) );
AOI211_X1 g_50_34 (.ZN (n_50_34), .A (n_47_37), .B (n_41_40), .C1 (n_40_39), .C2 (n_34_42) );
AOI211_X1 g_52_33 (.ZN (n_52_33), .A (n_49_36), .B (n_43_39), .C1 (n_42_38), .C2 (n_36_41) );
AOI211_X1 g_53_31 (.ZN (n_53_31), .A (n_50_34), .B (n_45_38), .C1 (n_41_40), .C2 (n_38_40) );
AOI211_X1 g_55_30 (.ZN (n_55_30), .A (n_52_33), .B (n_47_37), .C1 (n_43_39), .C2 (n_40_39) );
AOI211_X1 g_57_29 (.ZN (n_57_29), .A (n_53_31), .B (n_49_36), .C1 (n_45_38), .C2 (n_42_38) );
AOI211_X1 g_59_28 (.ZN (n_59_28), .A (n_55_30), .B (n_50_34), .C1 (n_47_37), .C2 (n_41_40) );
AOI211_X1 g_61_27 (.ZN (n_61_27), .A (n_57_29), .B (n_52_33), .C1 (n_49_36), .C2 (n_43_39) );
AOI211_X1 g_60_29 (.ZN (n_60_29), .A (n_59_28), .B (n_53_31), .C1 (n_50_34), .C2 (n_45_38) );
AOI211_X1 g_62_28 (.ZN (n_62_28), .A (n_61_27), .B (n_55_30), .C1 (n_52_33), .C2 (n_47_37) );
AOI211_X1 g_64_27 (.ZN (n_64_27), .A (n_60_29), .B (n_57_29), .C1 (n_53_31), .C2 (n_49_36) );
AOI211_X1 g_66_26 (.ZN (n_66_26), .A (n_62_28), .B (n_59_28), .C1 (n_55_30), .C2 (n_50_34) );
AOI211_X1 g_68_25 (.ZN (n_68_25), .A (n_64_27), .B (n_61_27), .C1 (n_57_29), .C2 (n_52_33) );
AOI211_X1 g_70_24 (.ZN (n_70_24), .A (n_66_26), .B (n_60_29), .C1 (n_59_28), .C2 (n_53_31) );
AOI211_X1 g_72_23 (.ZN (n_72_23), .A (n_68_25), .B (n_62_28), .C1 (n_61_27), .C2 (n_55_30) );
AOI211_X1 g_71_25 (.ZN (n_71_25), .A (n_70_24), .B (n_64_27), .C1 (n_60_29), .C2 (n_57_29) );
AOI211_X1 g_73_24 (.ZN (n_73_24), .A (n_72_23), .B (n_66_26), .C1 (n_62_28), .C2 (n_59_28) );
AOI211_X1 g_75_23 (.ZN (n_75_23), .A (n_71_25), .B (n_68_25), .C1 (n_64_27), .C2 (n_61_27) );
AOI211_X1 g_77_22 (.ZN (n_77_22), .A (n_73_24), .B (n_70_24), .C1 (n_66_26), .C2 (n_60_29) );
AOI211_X1 g_79_21 (.ZN (n_79_21), .A (n_75_23), .B (n_72_23), .C1 (n_68_25), .C2 (n_62_28) );
AOI211_X1 g_81_20 (.ZN (n_81_20), .A (n_77_22), .B (n_71_25), .C1 (n_70_24), .C2 (n_64_27) );
AOI211_X1 g_80_22 (.ZN (n_80_22), .A (n_79_21), .B (n_73_24), .C1 (n_72_23), .C2 (n_66_26) );
AOI211_X1 g_78_21 (.ZN (n_78_21), .A (n_81_20), .B (n_75_23), .C1 (n_71_25), .C2 (n_68_25) );
AOI211_X1 g_80_20 (.ZN (n_80_20), .A (n_80_22), .B (n_77_22), .C1 (n_73_24), .C2 (n_70_24) );
AOI211_X1 g_82_19 (.ZN (n_82_19), .A (n_78_21), .B (n_79_21), .C1 (n_75_23), .C2 (n_72_23) );
AOI211_X1 g_84_18 (.ZN (n_84_18), .A (n_80_20), .B (n_81_20), .C1 (n_77_22), .C2 (n_71_25) );
AOI211_X1 g_85_20 (.ZN (n_85_20), .A (n_82_19), .B (n_80_22), .C1 (n_79_21), .C2 (n_73_24) );
AOI211_X1 g_83_21 (.ZN (n_83_21), .A (n_84_18), .B (n_78_21), .C1 (n_81_20), .C2 (n_75_23) );
AOI211_X1 g_81_22 (.ZN (n_81_22), .A (n_85_20), .B (n_80_20), .C1 (n_80_22), .C2 (n_77_22) );
AOI211_X1 g_79_23 (.ZN (n_79_23), .A (n_83_21), .B (n_82_19), .C1 (n_78_21), .C2 (n_79_21) );
AOI211_X1 g_77_24 (.ZN (n_77_24), .A (n_81_22), .B (n_84_18), .C1 (n_80_20), .C2 (n_81_20) );
AOI211_X1 g_78_22 (.ZN (n_78_22), .A (n_79_23), .B (n_85_20), .C1 (n_82_19), .C2 (n_80_22) );
AOI211_X1 g_76_23 (.ZN (n_76_23), .A (n_77_24), .B (n_83_21), .C1 (n_84_18), .C2 (n_78_21) );
AOI211_X1 g_77_21 (.ZN (n_77_21), .A (n_78_22), .B (n_81_22), .C1 (n_85_20), .C2 (n_80_20) );
AOI211_X1 g_75_22 (.ZN (n_75_22), .A (n_76_23), .B (n_79_23), .C1 (n_83_21), .C2 (n_82_19) );
AOI211_X1 g_73_23 (.ZN (n_73_23), .A (n_77_21), .B (n_77_24), .C1 (n_81_22), .C2 (n_84_18) );
AOI211_X1 g_71_24 (.ZN (n_71_24), .A (n_75_22), .B (n_78_22), .C1 (n_79_23), .C2 (n_85_20) );
AOI211_X1 g_69_25 (.ZN (n_69_25), .A (n_73_23), .B (n_76_23), .C1 (n_77_24), .C2 (n_83_21) );
AOI211_X1 g_67_26 (.ZN (n_67_26), .A (n_71_24), .B (n_77_21), .C1 (n_78_22), .C2 (n_81_22) );
AOI211_X1 g_65_27 (.ZN (n_65_27), .A (n_69_25), .B (n_75_22), .C1 (n_76_23), .C2 (n_79_23) );
AOI211_X1 g_66_25 (.ZN (n_66_25), .A (n_67_26), .B (n_73_23), .C1 (n_77_21), .C2 (n_77_24) );
AOI211_X1 g_64_26 (.ZN (n_64_26), .A (n_65_27), .B (n_71_24), .C1 (n_75_22), .C2 (n_78_22) );
AOI211_X1 g_62_27 (.ZN (n_62_27), .A (n_66_25), .B (n_69_25), .C1 (n_73_23), .C2 (n_76_23) );
AOI211_X1 g_61_29 (.ZN (n_61_29), .A (n_64_26), .B (n_67_26), .C1 (n_71_24), .C2 (n_77_21) );
AOI211_X1 g_63_28 (.ZN (n_63_28), .A (n_62_27), .B (n_65_27), .C1 (n_69_25), .C2 (n_75_22) );
AOI211_X1 g_62_30 (.ZN (n_62_30), .A (n_61_29), .B (n_66_25), .C1 (n_67_26), .C2 (n_73_23) );
AOI211_X1 g_64_29 (.ZN (n_64_29), .A (n_63_28), .B (n_64_26), .C1 (n_65_27), .C2 (n_71_24) );
AOI211_X1 g_66_28 (.ZN (n_66_28), .A (n_62_30), .B (n_62_27), .C1 (n_66_25), .C2 (n_69_25) );
AOI211_X1 g_68_27 (.ZN (n_68_27), .A (n_64_29), .B (n_61_29), .C1 (n_64_26), .C2 (n_67_26) );
AOI211_X1 g_70_26 (.ZN (n_70_26), .A (n_66_28), .B (n_63_28), .C1 (n_62_27), .C2 (n_65_27) );
AOI211_X1 g_72_25 (.ZN (n_72_25), .A (n_68_27), .B (n_62_30), .C1 (n_61_29), .C2 (n_66_25) );
AOI211_X1 g_74_24 (.ZN (n_74_24), .A (n_70_26), .B (n_64_29), .C1 (n_63_28), .C2 (n_64_26) );
AOI211_X1 g_73_26 (.ZN (n_73_26), .A (n_72_25), .B (n_66_28), .C1 (n_62_30), .C2 (n_62_27) );
AOI211_X1 g_75_25 (.ZN (n_75_25), .A (n_74_24), .B (n_68_27), .C1 (n_64_29), .C2 (n_61_29) );
AOI211_X1 g_74_23 (.ZN (n_74_23), .A (n_73_26), .B (n_70_26), .C1 (n_66_28), .C2 (n_63_28) );
AOI211_X1 g_76_22 (.ZN (n_76_22), .A (n_75_25), .B (n_72_25), .C1 (n_68_27), .C2 (n_62_30) );
AOI211_X1 g_78_23 (.ZN (n_78_23), .A (n_74_23), .B (n_74_24), .C1 (n_70_26), .C2 (n_64_29) );
AOI211_X1 g_76_24 (.ZN (n_76_24), .A (n_76_22), .B (n_73_26), .C1 (n_72_25), .C2 (n_66_28) );
AOI211_X1 g_74_25 (.ZN (n_74_25), .A (n_78_23), .B (n_75_25), .C1 (n_74_24), .C2 (n_68_27) );
AOI211_X1 g_72_24 (.ZN (n_72_24), .A (n_76_24), .B (n_74_23), .C1 (n_73_26), .C2 (n_70_26) );
AOI211_X1 g_70_25 (.ZN (n_70_25), .A (n_74_25), .B (n_76_22), .C1 (n_75_25), .C2 (n_72_25) );
AOI211_X1 g_68_26 (.ZN (n_68_26), .A (n_72_24), .B (n_78_23), .C1 (n_74_23), .C2 (n_74_24) );
AOI211_X1 g_66_27 (.ZN (n_66_27), .A (n_70_25), .B (n_76_24), .C1 (n_76_22), .C2 (n_73_26) );
AOI211_X1 g_64_28 (.ZN (n_64_28), .A (n_68_26), .B (n_74_25), .C1 (n_78_23), .C2 (n_75_25) );
AOI211_X1 g_62_29 (.ZN (n_62_29), .A (n_66_27), .B (n_72_24), .C1 (n_76_24), .C2 (n_74_23) );
AOI211_X1 g_60_30 (.ZN (n_60_30), .A (n_64_28), .B (n_70_25), .C1 (n_74_25), .C2 (n_76_22) );
AOI211_X1 g_58_31 (.ZN (n_58_31), .A (n_62_29), .B (n_68_26), .C1 (n_72_24), .C2 (n_78_23) );
AOI211_X1 g_56_32 (.ZN (n_56_32), .A (n_60_30), .B (n_66_27), .C1 (n_70_25), .C2 (n_76_24) );
AOI211_X1 g_54_33 (.ZN (n_54_33), .A (n_58_31), .B (n_64_28), .C1 (n_68_26), .C2 (n_74_25) );
AOI211_X1 g_52_34 (.ZN (n_52_34), .A (n_56_32), .B (n_62_29), .C1 (n_66_27), .C2 (n_72_24) );
AOI211_X1 g_50_35 (.ZN (n_50_35), .A (n_54_33), .B (n_60_30), .C1 (n_64_28), .C2 (n_70_25) );
AOI211_X1 g_48_36 (.ZN (n_48_36), .A (n_52_34), .B (n_58_31), .C1 (n_62_29), .C2 (n_68_26) );
AOI211_X1 g_46_37 (.ZN (n_46_37), .A (n_50_35), .B (n_56_32), .C1 (n_60_30), .C2 (n_66_27) );
AOI211_X1 g_45_39 (.ZN (n_45_39), .A (n_48_36), .B (n_54_33), .C1 (n_58_31), .C2 (n_64_28) );
AOI211_X1 g_47_38 (.ZN (n_47_38), .A (n_46_37), .B (n_52_34), .C1 (n_56_32), .C2 (n_62_29) );
AOI211_X1 g_49_37 (.ZN (n_49_37), .A (n_45_39), .B (n_50_35), .C1 (n_54_33), .C2 (n_60_30) );
AOI211_X1 g_51_36 (.ZN (n_51_36), .A (n_47_38), .B (n_48_36), .C1 (n_52_34), .C2 (n_58_31) );
AOI211_X1 g_53_35 (.ZN (n_53_35), .A (n_49_37), .B (n_46_37), .C1 (n_50_35), .C2 (n_56_32) );
AOI211_X1 g_55_34 (.ZN (n_55_34), .A (n_51_36), .B (n_45_39), .C1 (n_48_36), .C2 (n_54_33) );
AOI211_X1 g_54_32 (.ZN (n_54_32), .A (n_53_35), .B (n_47_38), .C1 (n_46_37), .C2 (n_52_34) );
AOI211_X1 g_56_31 (.ZN (n_56_31), .A (n_55_34), .B (n_49_37), .C1 (n_45_39), .C2 (n_50_35) );
AOI211_X1 g_58_30 (.ZN (n_58_30), .A (n_54_32), .B (n_51_36), .C1 (n_47_38), .C2 (n_48_36) );
AOI211_X1 g_60_31 (.ZN (n_60_31), .A (n_56_31), .B (n_53_35), .C1 (n_49_37), .C2 (n_46_37) );
AOI211_X1 g_58_32 (.ZN (n_58_32), .A (n_58_30), .B (n_55_34), .C1 (n_51_36), .C2 (n_45_39) );
AOI211_X1 g_59_30 (.ZN (n_59_30), .A (n_60_31), .B (n_54_32), .C1 (n_53_35), .C2 (n_47_38) );
AOI211_X1 g_57_31 (.ZN (n_57_31), .A (n_58_32), .B (n_56_31), .C1 (n_55_34), .C2 (n_49_37) );
AOI211_X1 g_55_32 (.ZN (n_55_32), .A (n_59_30), .B (n_58_30), .C1 (n_54_32), .C2 (n_51_36) );
AOI211_X1 g_57_33 (.ZN (n_57_33), .A (n_57_31), .B (n_60_31), .C1 (n_56_31), .C2 (n_53_35) );
AOI211_X1 g_59_32 (.ZN (n_59_32), .A (n_55_32), .B (n_58_32), .C1 (n_58_30), .C2 (n_55_34) );
AOI211_X1 g_61_31 (.ZN (n_61_31), .A (n_57_33), .B (n_59_30), .C1 (n_60_31), .C2 (n_54_32) );
AOI211_X1 g_63_30 (.ZN (n_63_30), .A (n_59_32), .B (n_57_31), .C1 (n_58_32), .C2 (n_56_31) );
AOI211_X1 g_65_29 (.ZN (n_65_29), .A (n_61_31), .B (n_55_32), .C1 (n_59_30), .C2 (n_58_30) );
AOI211_X1 g_67_28 (.ZN (n_67_28), .A (n_63_30), .B (n_57_33), .C1 (n_57_31), .C2 (n_60_31) );
AOI211_X1 g_69_27 (.ZN (n_69_27), .A (n_65_29), .B (n_59_32), .C1 (n_55_32), .C2 (n_58_32) );
AOI211_X1 g_71_26 (.ZN (n_71_26), .A (n_67_28), .B (n_61_31), .C1 (n_57_33), .C2 (n_59_30) );
AOI211_X1 g_73_25 (.ZN (n_73_25), .A (n_69_27), .B (n_63_30), .C1 (n_59_32), .C2 (n_57_31) );
AOI211_X1 g_75_24 (.ZN (n_75_24), .A (n_71_26), .B (n_65_29), .C1 (n_61_31), .C2 (n_55_32) );
AOI211_X1 g_77_23 (.ZN (n_77_23), .A (n_73_25), .B (n_67_28), .C1 (n_63_30), .C2 (n_57_33) );
AOI211_X1 g_79_22 (.ZN (n_79_22), .A (n_75_24), .B (n_69_27), .C1 (n_65_29), .C2 (n_59_32) );
AOI211_X1 g_81_21 (.ZN (n_81_21), .A (n_77_23), .B (n_71_26), .C1 (n_67_28), .C2 (n_61_31) );
AOI211_X1 g_83_20 (.ZN (n_83_20), .A (n_79_22), .B (n_73_25), .C1 (n_69_27), .C2 (n_63_30) );
AOI211_X1 g_85_19 (.ZN (n_85_19), .A (n_81_21), .B (n_75_24), .C1 (n_71_26), .C2 (n_65_29) );
AOI211_X1 g_87_18 (.ZN (n_87_18), .A (n_83_20), .B (n_77_23), .C1 (n_73_25), .C2 (n_67_28) );
AOI211_X1 g_89_17 (.ZN (n_89_17), .A (n_85_19), .B (n_79_22), .C1 (n_75_24), .C2 (n_69_27) );
AOI211_X1 g_91_16 (.ZN (n_91_16), .A (n_87_18), .B (n_81_21), .C1 (n_77_23), .C2 (n_71_26) );
AOI211_X1 g_93_17 (.ZN (n_93_17), .A (n_89_17), .B (n_83_20), .C1 (n_79_22), .C2 (n_73_25) );
AOI211_X1 g_91_18 (.ZN (n_91_18), .A (n_91_16), .B (n_85_19), .C1 (n_81_21), .C2 (n_75_24) );
AOI211_X1 g_89_19 (.ZN (n_89_19), .A (n_93_17), .B (n_87_18), .C1 (n_83_20), .C2 (n_77_23) );
AOI211_X1 g_87_20 (.ZN (n_87_20), .A (n_91_18), .B (n_89_17), .C1 (n_85_19), .C2 (n_79_22) );
AOI211_X1 g_88_18 (.ZN (n_88_18), .A (n_89_19), .B (n_91_16), .C1 (n_87_18), .C2 (n_81_21) );
AOI211_X1 g_86_19 (.ZN (n_86_19), .A (n_87_20), .B (n_93_17), .C1 (n_89_17), .C2 (n_83_20) );
AOI211_X1 g_84_20 (.ZN (n_84_20), .A (n_88_18), .B (n_91_18), .C1 (n_91_16), .C2 (n_85_19) );
AOI211_X1 g_82_21 (.ZN (n_82_21), .A (n_86_19), .B (n_89_19), .C1 (n_93_17), .C2 (n_87_18) );
AOI211_X1 g_81_23 (.ZN (n_81_23), .A (n_84_20), .B (n_87_20), .C1 (n_91_18), .C2 (n_89_17) );
AOI211_X1 g_83_22 (.ZN (n_83_22), .A (n_82_21), .B (n_88_18), .C1 (n_89_19), .C2 (n_91_16) );
AOI211_X1 g_85_21 (.ZN (n_85_21), .A (n_81_23), .B (n_86_19), .C1 (n_87_20), .C2 (n_93_17) );
AOI211_X1 g_84_23 (.ZN (n_84_23), .A (n_83_22), .B (n_84_20), .C1 (n_88_18), .C2 (n_91_18) );
AOI211_X1 g_82_22 (.ZN (n_82_22), .A (n_85_21), .B (n_82_21), .C1 (n_86_19), .C2 (n_89_19) );
AOI211_X1 g_84_21 (.ZN (n_84_21), .A (n_84_23), .B (n_81_23), .C1 (n_84_20), .C2 (n_87_20) );
AOI211_X1 g_86_20 (.ZN (n_86_20), .A (n_82_22), .B (n_83_22), .C1 (n_82_21), .C2 (n_88_18) );
AOI211_X1 g_88_19 (.ZN (n_88_19), .A (n_84_21), .B (n_85_21), .C1 (n_81_23), .C2 (n_86_19) );
AOI211_X1 g_90_18 (.ZN (n_90_18), .A (n_86_20), .B (n_84_23), .C1 (n_83_22), .C2 (n_84_20) );
AOI211_X1 g_92_17 (.ZN (n_92_17), .A (n_88_19), .B (n_82_22), .C1 (n_85_21), .C2 (n_82_21) );
AOI211_X1 g_91_19 (.ZN (n_91_19), .A (n_90_18), .B (n_84_21), .C1 (n_84_23), .C2 (n_81_23) );
AOI211_X1 g_89_20 (.ZN (n_89_20), .A (n_92_17), .B (n_86_20), .C1 (n_82_22), .C2 (n_83_22) );
AOI211_X1 g_87_21 (.ZN (n_87_21), .A (n_91_19), .B (n_88_19), .C1 (n_84_21), .C2 (n_85_21) );
AOI211_X1 g_85_22 (.ZN (n_85_22), .A (n_89_20), .B (n_90_18), .C1 (n_86_20), .C2 (n_84_23) );
AOI211_X1 g_83_23 (.ZN (n_83_23), .A (n_87_21), .B (n_92_17), .C1 (n_88_19), .C2 (n_82_22) );
AOI211_X1 g_81_24 (.ZN (n_81_24), .A (n_85_22), .B (n_91_19), .C1 (n_90_18), .C2 (n_84_21) );
AOI211_X1 g_79_25 (.ZN (n_79_25), .A (n_83_23), .B (n_89_20), .C1 (n_92_17), .C2 (n_86_20) );
AOI211_X1 g_80_23 (.ZN (n_80_23), .A (n_81_24), .B (n_87_21), .C1 (n_91_19), .C2 (n_88_19) );
AOI211_X1 g_78_24 (.ZN (n_78_24), .A (n_79_25), .B (n_85_22), .C1 (n_89_20), .C2 (n_90_18) );
AOI211_X1 g_76_25 (.ZN (n_76_25), .A (n_80_23), .B (n_83_23), .C1 (n_87_21), .C2 (n_92_17) );
AOI211_X1 g_74_26 (.ZN (n_74_26), .A (n_78_24), .B (n_81_24), .C1 (n_85_22), .C2 (n_91_19) );
AOI211_X1 g_72_27 (.ZN (n_72_27), .A (n_76_25), .B (n_79_25), .C1 (n_83_23), .C2 (n_89_20) );
AOI211_X1 g_70_28 (.ZN (n_70_28), .A (n_74_26), .B (n_80_23), .C1 (n_81_24), .C2 (n_87_21) );
AOI211_X1 g_69_26 (.ZN (n_69_26), .A (n_72_27), .B (n_78_24), .C1 (n_79_25), .C2 (n_85_22) );
AOI211_X1 g_67_27 (.ZN (n_67_27), .A (n_70_28), .B (n_76_25), .C1 (n_80_23), .C2 (n_83_23) );
AOI211_X1 g_65_28 (.ZN (n_65_28), .A (n_69_26), .B (n_74_26), .C1 (n_78_24), .C2 (n_81_24) );
AOI211_X1 g_63_29 (.ZN (n_63_29), .A (n_67_27), .B (n_72_27), .C1 (n_76_25), .C2 (n_79_25) );
AOI211_X1 g_61_30 (.ZN (n_61_30), .A (n_65_28), .B (n_70_28), .C1 (n_74_26), .C2 (n_80_23) );
AOI211_X1 g_59_31 (.ZN (n_59_31), .A (n_63_29), .B (n_69_26), .C1 (n_72_27), .C2 (n_78_24) );
AOI211_X1 g_57_32 (.ZN (n_57_32), .A (n_61_30), .B (n_67_27), .C1 (n_70_28), .C2 (n_76_25) );
AOI211_X1 g_55_33 (.ZN (n_55_33), .A (n_59_31), .B (n_65_28), .C1 (n_69_26), .C2 (n_74_26) );
AOI211_X1 g_53_34 (.ZN (n_53_34), .A (n_57_32), .B (n_63_29), .C1 (n_67_27), .C2 (n_72_27) );
AOI211_X1 g_51_35 (.ZN (n_51_35), .A (n_55_33), .B (n_61_30), .C1 (n_65_28), .C2 (n_70_28) );
AOI211_X1 g_50_37 (.ZN (n_50_37), .A (n_53_34), .B (n_59_31), .C1 (n_63_29), .C2 (n_69_26) );
AOI211_X1 g_52_36 (.ZN (n_52_36), .A (n_51_35), .B (n_57_32), .C1 (n_61_30), .C2 (n_67_27) );
AOI211_X1 g_54_35 (.ZN (n_54_35), .A (n_50_37), .B (n_55_33), .C1 (n_59_31), .C2 (n_65_28) );
AOI211_X1 g_56_34 (.ZN (n_56_34), .A (n_52_36), .B (n_53_34), .C1 (n_57_32), .C2 (n_63_29) );
AOI211_X1 g_58_33 (.ZN (n_58_33), .A (n_54_35), .B (n_51_35), .C1 (n_55_33), .C2 (n_61_30) );
AOI211_X1 g_60_32 (.ZN (n_60_32), .A (n_56_34), .B (n_50_37), .C1 (n_53_34), .C2 (n_59_31) );
AOI211_X1 g_62_31 (.ZN (n_62_31), .A (n_58_33), .B (n_52_36), .C1 (n_51_35), .C2 (n_57_32) );
AOI211_X1 g_64_30 (.ZN (n_64_30), .A (n_60_32), .B (n_54_35), .C1 (n_50_37), .C2 (n_55_33) );
AOI211_X1 g_66_29 (.ZN (n_66_29), .A (n_62_31), .B (n_56_34), .C1 (n_52_36), .C2 (n_53_34) );
AOI211_X1 g_68_28 (.ZN (n_68_28), .A (n_64_30), .B (n_58_33), .C1 (n_54_35), .C2 (n_51_35) );
AOI211_X1 g_70_27 (.ZN (n_70_27), .A (n_66_29), .B (n_60_32), .C1 (n_56_34), .C2 (n_50_37) );
AOI211_X1 g_72_26 (.ZN (n_72_26), .A (n_68_28), .B (n_62_31), .C1 (n_58_33), .C2 (n_52_36) );
AOI211_X1 g_71_28 (.ZN (n_71_28), .A (n_70_27), .B (n_64_30), .C1 (n_60_32), .C2 (n_54_35) );
AOI211_X1 g_73_27 (.ZN (n_73_27), .A (n_72_26), .B (n_66_29), .C1 (n_62_31), .C2 (n_56_34) );
AOI211_X1 g_75_26 (.ZN (n_75_26), .A (n_71_28), .B (n_68_28), .C1 (n_64_30), .C2 (n_58_33) );
AOI211_X1 g_77_25 (.ZN (n_77_25), .A (n_73_27), .B (n_70_27), .C1 (n_66_29), .C2 (n_60_32) );
AOI211_X1 g_79_24 (.ZN (n_79_24), .A (n_75_26), .B (n_72_26), .C1 (n_68_28), .C2 (n_62_31) );
AOI211_X1 g_78_26 (.ZN (n_78_26), .A (n_77_25), .B (n_71_28), .C1 (n_70_27), .C2 (n_64_30) );
AOI211_X1 g_80_25 (.ZN (n_80_25), .A (n_79_24), .B (n_73_27), .C1 (n_72_26), .C2 (n_66_29) );
AOI211_X1 g_82_24 (.ZN (n_82_24), .A (n_78_26), .B (n_75_26), .C1 (n_71_28), .C2 (n_68_28) );
AOI211_X1 g_81_26 (.ZN (n_81_26), .A (n_80_25), .B (n_77_25), .C1 (n_73_27), .C2 (n_70_27) );
AOI211_X1 g_80_24 (.ZN (n_80_24), .A (n_82_24), .B (n_79_24), .C1 (n_75_26), .C2 (n_72_26) );
AOI211_X1 g_82_23 (.ZN (n_82_23), .A (n_81_26), .B (n_78_26), .C1 (n_77_25), .C2 (n_71_28) );
AOI211_X1 g_84_22 (.ZN (n_84_22), .A (n_80_24), .B (n_80_25), .C1 (n_79_24), .C2 (n_73_27) );
AOI211_X1 g_86_21 (.ZN (n_86_21), .A (n_82_23), .B (n_82_24), .C1 (n_78_26), .C2 (n_75_26) );
AOI211_X1 g_88_20 (.ZN (n_88_20), .A (n_84_22), .B (n_81_26), .C1 (n_80_25), .C2 (n_77_25) );
AOI211_X1 g_90_19 (.ZN (n_90_19), .A (n_86_21), .B (n_80_24), .C1 (n_82_24), .C2 (n_79_24) );
AOI211_X1 g_92_18 (.ZN (n_92_18), .A (n_88_20), .B (n_82_23), .C1 (n_81_26), .C2 (n_78_26) );
AOI211_X1 g_94_19 (.ZN (n_94_19), .A (n_90_19), .B (n_84_22), .C1 (n_80_24), .C2 (n_80_25) );
AOI211_X1 g_92_20 (.ZN (n_92_20), .A (n_92_18), .B (n_86_21), .C1 (n_82_23), .C2 (n_82_24) );
AOI211_X1 g_90_21 (.ZN (n_90_21), .A (n_94_19), .B (n_88_20), .C1 (n_84_22), .C2 (n_81_26) );
AOI211_X1 g_88_22 (.ZN (n_88_22), .A (n_92_20), .B (n_90_19), .C1 (n_86_21), .C2 (n_80_24) );
AOI211_X1 g_86_23 (.ZN (n_86_23), .A (n_90_21), .B (n_92_18), .C1 (n_88_20), .C2 (n_82_23) );
AOI211_X1 g_84_24 (.ZN (n_84_24), .A (n_88_22), .B (n_94_19), .C1 (n_90_19), .C2 (n_84_22) );
AOI211_X1 g_82_25 (.ZN (n_82_25), .A (n_86_23), .B (n_92_20), .C1 (n_92_18), .C2 (n_86_21) );
AOI211_X1 g_80_26 (.ZN (n_80_26), .A (n_84_24), .B (n_90_21), .C1 (n_94_19), .C2 (n_88_20) );
AOI211_X1 g_78_25 (.ZN (n_78_25), .A (n_82_25), .B (n_88_22), .C1 (n_92_20), .C2 (n_90_19) );
AOI211_X1 g_76_26 (.ZN (n_76_26), .A (n_80_26), .B (n_86_23), .C1 (n_90_21), .C2 (n_92_18) );
AOI211_X1 g_74_27 (.ZN (n_74_27), .A (n_78_25), .B (n_84_24), .C1 (n_88_22), .C2 (n_94_19) );
AOI211_X1 g_72_28 (.ZN (n_72_28), .A (n_76_26), .B (n_82_25), .C1 (n_86_23), .C2 (n_92_20) );
AOI211_X1 g_70_29 (.ZN (n_70_29), .A (n_74_27), .B (n_80_26), .C1 (n_84_24), .C2 (n_90_21) );
AOI211_X1 g_71_27 (.ZN (n_71_27), .A (n_72_28), .B (n_78_25), .C1 (n_82_25), .C2 (n_88_22) );
AOI211_X1 g_69_28 (.ZN (n_69_28), .A (n_70_29), .B (n_76_26), .C1 (n_80_26), .C2 (n_86_23) );
AOI211_X1 g_67_29 (.ZN (n_67_29), .A (n_71_27), .B (n_74_27), .C1 (n_78_25), .C2 (n_84_24) );
AOI211_X1 g_65_30 (.ZN (n_65_30), .A (n_69_28), .B (n_72_28), .C1 (n_76_26), .C2 (n_82_25) );
AOI211_X1 g_63_31 (.ZN (n_63_31), .A (n_67_29), .B (n_70_29), .C1 (n_74_27), .C2 (n_80_26) );
AOI211_X1 g_61_32 (.ZN (n_61_32), .A (n_65_30), .B (n_71_27), .C1 (n_72_28), .C2 (n_78_25) );
AOI211_X1 g_59_33 (.ZN (n_59_33), .A (n_63_31), .B (n_69_28), .C1 (n_70_29), .C2 (n_76_26) );
AOI211_X1 g_57_34 (.ZN (n_57_34), .A (n_61_32), .B (n_67_29), .C1 (n_71_27), .C2 (n_74_27) );
AOI211_X1 g_55_35 (.ZN (n_55_35), .A (n_59_33), .B (n_65_30), .C1 (n_69_28), .C2 (n_72_28) );
AOI211_X1 g_56_33 (.ZN (n_56_33), .A (n_57_34), .B (n_63_31), .C1 (n_67_29), .C2 (n_70_29) );
AOI211_X1 g_54_34 (.ZN (n_54_34), .A (n_55_35), .B (n_61_32), .C1 (n_65_30), .C2 (n_71_27) );
AOI211_X1 g_52_35 (.ZN (n_52_35), .A (n_56_33), .B (n_59_33), .C1 (n_63_31), .C2 (n_69_28) );
AOI211_X1 g_50_36 (.ZN (n_50_36), .A (n_54_34), .B (n_57_34), .C1 (n_61_32), .C2 (n_67_29) );
AOI211_X1 g_48_37 (.ZN (n_48_37), .A (n_52_35), .B (n_55_35), .C1 (n_59_33), .C2 (n_65_30) );
AOI211_X1 g_46_38 (.ZN (n_46_38), .A (n_50_36), .B (n_56_33), .C1 (n_57_34), .C2 (n_63_31) );
AOI211_X1 g_44_39 (.ZN (n_44_39), .A (n_48_37), .B (n_54_34), .C1 (n_55_35), .C2 (n_61_32) );
AOI211_X1 g_42_40 (.ZN (n_42_40), .A (n_46_38), .B (n_52_35), .C1 (n_56_33), .C2 (n_59_33) );
AOI211_X1 g_40_41 (.ZN (n_40_41), .A (n_44_39), .B (n_50_36), .C1 (n_54_34), .C2 (n_57_34) );
AOI211_X1 g_38_42 (.ZN (n_38_42), .A (n_42_40), .B (n_48_37), .C1 (n_52_35), .C2 (n_55_35) );
AOI211_X1 g_39_40 (.ZN (n_39_40), .A (n_40_41), .B (n_46_38), .C1 (n_50_36), .C2 (n_56_33) );
AOI211_X1 g_37_41 (.ZN (n_37_41), .A (n_38_42), .B (n_44_39), .C1 (n_48_37), .C2 (n_54_34) );
AOI211_X1 g_35_42 (.ZN (n_35_42), .A (n_39_40), .B (n_42_40), .C1 (n_46_38), .C2 (n_52_35) );
AOI211_X1 g_33_43 (.ZN (n_33_43), .A (n_37_41), .B (n_40_41), .C1 (n_44_39), .C2 (n_50_36) );
AOI211_X1 g_31_44 (.ZN (n_31_44), .A (n_35_42), .B (n_38_42), .C1 (n_42_40), .C2 (n_48_37) );
AOI211_X1 g_29_45 (.ZN (n_29_45), .A (n_33_43), .B (n_39_40), .C1 (n_40_41), .C2 (n_46_38) );
AOI211_X1 g_27_46 (.ZN (n_27_46), .A (n_31_44), .B (n_37_41), .C1 (n_38_42), .C2 (n_44_39) );
AOI211_X1 g_25_47 (.ZN (n_25_47), .A (n_29_45), .B (n_35_42), .C1 (n_39_40), .C2 (n_42_40) );
AOI211_X1 g_23_48 (.ZN (n_23_48), .A (n_27_46), .B (n_33_43), .C1 (n_37_41), .C2 (n_40_41) );
AOI211_X1 g_21_49 (.ZN (n_21_49), .A (n_25_47), .B (n_31_44), .C1 (n_35_42), .C2 (n_38_42) );
AOI211_X1 g_20_47 (.ZN (n_20_47), .A (n_23_48), .B (n_29_45), .C1 (n_33_43), .C2 (n_39_40) );
AOI211_X1 g_18_48 (.ZN (n_18_48), .A (n_21_49), .B (n_27_46), .C1 (n_31_44), .C2 (n_37_41) );
AOI211_X1 g_16_49 (.ZN (n_16_49), .A (n_20_47), .B (n_25_47), .C1 (n_29_45), .C2 (n_35_42) );
AOI211_X1 g_14_50 (.ZN (n_14_50), .A (n_18_48), .B (n_23_48), .C1 (n_27_46), .C2 (n_33_43) );
AOI211_X1 g_12_51 (.ZN (n_12_51), .A (n_16_49), .B (n_21_49), .C1 (n_25_47), .C2 (n_31_44) );
AOI211_X1 g_10_52 (.ZN (n_10_52), .A (n_14_50), .B (n_20_47), .C1 (n_23_48), .C2 (n_29_45) );
AOI211_X1 g_8_53 (.ZN (n_8_53), .A (n_12_51), .B (n_18_48), .C1 (n_21_49), .C2 (n_27_46) );
AOI211_X1 g_6_54 (.ZN (n_6_54), .A (n_10_52), .B (n_16_49), .C1 (n_20_47), .C2 (n_25_47) );
AOI211_X1 g_8_55 (.ZN (n_8_55), .A (n_8_53), .B (n_14_50), .C1 (n_18_48), .C2 (n_23_48) );
AOI211_X1 g_10_54 (.ZN (n_10_54), .A (n_6_54), .B (n_12_51), .C1 (n_16_49), .C2 (n_21_49) );
AOI211_X1 g_12_53 (.ZN (n_12_53), .A (n_8_55), .B (n_10_52), .C1 (n_14_50), .C2 (n_20_47) );
AOI211_X1 g_14_52 (.ZN (n_14_52), .A (n_10_54), .B (n_8_53), .C1 (n_12_51), .C2 (n_18_48) );
AOI211_X1 g_16_51 (.ZN (n_16_51), .A (n_12_53), .B (n_6_54), .C1 (n_10_52), .C2 (n_16_49) );
AOI211_X1 g_18_50 (.ZN (n_18_50), .A (n_14_52), .B (n_8_55), .C1 (n_8_53), .C2 (n_14_50) );
AOI211_X1 g_20_49 (.ZN (n_20_49), .A (n_16_51), .B (n_10_54), .C1 (n_6_54), .C2 (n_12_51) );
AOI211_X1 g_22_48 (.ZN (n_22_48), .A (n_18_50), .B (n_12_53), .C1 (n_8_55), .C2 (n_10_52) );
AOI211_X1 g_23_50 (.ZN (n_23_50), .A (n_20_49), .B (n_14_52), .C1 (n_10_54), .C2 (n_8_53) );
AOI211_X1 g_24_48 (.ZN (n_24_48), .A (n_22_48), .B (n_16_51), .C1 (n_12_53), .C2 (n_6_54) );
AOI211_X1 g_26_47 (.ZN (n_26_47), .A (n_23_50), .B (n_18_50), .C1 (n_14_52), .C2 (n_8_55) );
AOI211_X1 g_25_49 (.ZN (n_25_49), .A (n_24_48), .B (n_20_49), .C1 (n_16_51), .C2 (n_10_54) );
AOI211_X1 g_27_48 (.ZN (n_27_48), .A (n_26_47), .B (n_22_48), .C1 (n_18_50), .C2 (n_12_53) );
AOI211_X1 g_26_46 (.ZN (n_26_46), .A (n_25_49), .B (n_23_50), .C1 (n_20_49), .C2 (n_14_52) );
AOI211_X1 g_28_45 (.ZN (n_28_45), .A (n_27_48), .B (n_24_48), .C1 (n_22_48), .C2 (n_16_51) );
AOI211_X1 g_30_44 (.ZN (n_30_44), .A (n_26_46), .B (n_26_47), .C1 (n_23_50), .C2 (n_18_50) );
AOI211_X1 g_31_46 (.ZN (n_31_46), .A (n_28_45), .B (n_25_49), .C1 (n_24_48), .C2 (n_20_49) );
AOI211_X1 g_29_47 (.ZN (n_29_47), .A (n_30_44), .B (n_27_48), .C1 (n_26_47), .C2 (n_22_48) );
AOI211_X1 g_28_49 (.ZN (n_28_49), .A (n_31_46), .B (n_26_46), .C1 (n_25_49), .C2 (n_23_50) );
AOI211_X1 g_27_47 (.ZN (n_27_47), .A (n_29_47), .B (n_28_45), .C1 (n_27_48), .C2 (n_24_48) );
AOI211_X1 g_29_46 (.ZN (n_29_46), .A (n_28_49), .B (n_30_44), .C1 (n_26_46), .C2 (n_26_47) );
AOI211_X1 g_31_45 (.ZN (n_31_45), .A (n_27_47), .B (n_31_46), .C1 (n_28_45), .C2 (n_25_49) );
AOI211_X1 g_33_44 (.ZN (n_33_44), .A (n_29_46), .B (n_29_47), .C1 (n_30_44), .C2 (n_27_48) );
AOI211_X1 g_35_43 (.ZN (n_35_43), .A (n_31_45), .B (n_28_49), .C1 (n_31_46), .C2 (n_26_46) );
AOI211_X1 g_37_42 (.ZN (n_37_42), .A (n_33_44), .B (n_27_47), .C1 (n_29_47), .C2 (n_28_45) );
AOI211_X1 g_39_41 (.ZN (n_39_41), .A (n_35_43), .B (n_29_46), .C1 (n_28_49), .C2 (n_30_44) );
AOI211_X1 g_38_43 (.ZN (n_38_43), .A (n_37_42), .B (n_31_45), .C1 (n_27_47), .C2 (n_31_46) );
AOI211_X1 g_40_42 (.ZN (n_40_42), .A (n_39_41), .B (n_33_44), .C1 (n_29_46), .C2 (n_29_47) );
AOI211_X1 g_42_41 (.ZN (n_42_41), .A (n_38_43), .B (n_35_43), .C1 (n_31_45), .C2 (n_28_49) );
AOI211_X1 g_44_40 (.ZN (n_44_40), .A (n_40_42), .B (n_37_42), .C1 (n_33_44), .C2 (n_27_47) );
AOI211_X1 g_46_39 (.ZN (n_46_39), .A (n_42_41), .B (n_39_41), .C1 (n_35_43), .C2 (n_29_46) );
AOI211_X1 g_48_38 (.ZN (n_48_38), .A (n_44_40), .B (n_38_43), .C1 (n_37_42), .C2 (n_31_45) );
AOI211_X1 g_47_40 (.ZN (n_47_40), .A (n_46_39), .B (n_40_42), .C1 (n_39_41), .C2 (n_33_44) );
AOI211_X1 g_49_39 (.ZN (n_49_39), .A (n_48_38), .B (n_42_41), .C1 (n_38_43), .C2 (n_35_43) );
AOI211_X1 g_51_38 (.ZN (n_51_38), .A (n_47_40), .B (n_44_40), .C1 (n_40_42), .C2 (n_37_42) );
AOI211_X1 g_53_37 (.ZN (n_53_37), .A (n_49_39), .B (n_46_39), .C1 (n_42_41), .C2 (n_39_41) );
AOI211_X1 g_55_36 (.ZN (n_55_36), .A (n_51_38), .B (n_48_38), .C1 (n_44_40), .C2 (n_38_43) );
AOI211_X1 g_57_35 (.ZN (n_57_35), .A (n_53_37), .B (n_47_40), .C1 (n_46_39), .C2 (n_40_42) );
AOI211_X1 g_59_34 (.ZN (n_59_34), .A (n_55_36), .B (n_49_39), .C1 (n_48_38), .C2 (n_42_41) );
AOI211_X1 g_61_33 (.ZN (n_61_33), .A (n_57_35), .B (n_51_38), .C1 (n_47_40), .C2 (n_44_40) );
AOI211_X1 g_63_32 (.ZN (n_63_32), .A (n_59_34), .B (n_53_37), .C1 (n_49_39), .C2 (n_46_39) );
AOI211_X1 g_65_31 (.ZN (n_65_31), .A (n_61_33), .B (n_55_36), .C1 (n_51_38), .C2 (n_48_38) );
AOI211_X1 g_67_30 (.ZN (n_67_30), .A (n_63_32), .B (n_57_35), .C1 (n_53_37), .C2 (n_47_40) );
AOI211_X1 g_69_29 (.ZN (n_69_29), .A (n_65_31), .B (n_59_34), .C1 (n_55_36), .C2 (n_49_39) );
AOI211_X1 g_71_30 (.ZN (n_71_30), .A (n_67_30), .B (n_61_33), .C1 (n_57_35), .C2 (n_51_38) );
AOI211_X1 g_73_29 (.ZN (n_73_29), .A (n_69_29), .B (n_63_32), .C1 (n_59_34), .C2 (n_53_37) );
AOI211_X1 g_75_28 (.ZN (n_75_28), .A (n_71_30), .B (n_65_31), .C1 (n_61_33), .C2 (n_55_36) );
AOI211_X1 g_77_27 (.ZN (n_77_27), .A (n_73_29), .B (n_67_30), .C1 (n_63_32), .C2 (n_57_35) );
AOI211_X1 g_79_26 (.ZN (n_79_26), .A (n_75_28), .B (n_69_29), .C1 (n_65_31), .C2 (n_59_34) );
AOI211_X1 g_81_25 (.ZN (n_81_25), .A (n_77_27), .B (n_71_30), .C1 (n_67_30), .C2 (n_61_33) );
AOI211_X1 g_83_24 (.ZN (n_83_24), .A (n_79_26), .B (n_73_29), .C1 (n_69_29), .C2 (n_63_32) );
AOI211_X1 g_85_23 (.ZN (n_85_23), .A (n_81_25), .B (n_75_28), .C1 (n_71_30), .C2 (n_65_31) );
AOI211_X1 g_87_22 (.ZN (n_87_22), .A (n_83_24), .B (n_77_27), .C1 (n_73_29), .C2 (n_67_30) );
AOI211_X1 g_89_21 (.ZN (n_89_21), .A (n_85_23), .B (n_79_26), .C1 (n_75_28), .C2 (n_69_29) );
AOI211_X1 g_91_20 (.ZN (n_91_20), .A (n_87_22), .B (n_81_25), .C1 (n_77_27), .C2 (n_71_30) );
AOI211_X1 g_93_19 (.ZN (n_93_19), .A (n_89_21), .B (n_83_24), .C1 (n_79_26), .C2 (n_73_29) );
AOI211_X1 g_94_21 (.ZN (n_94_21), .A (n_91_20), .B (n_85_23), .C1 (n_81_25), .C2 (n_75_28) );
AOI211_X1 g_96_20 (.ZN (n_96_20), .A (n_93_19), .B (n_87_22), .C1 (n_83_24), .C2 (n_77_27) );
AOI211_X1 g_98_19 (.ZN (n_98_19), .A (n_94_21), .B (n_89_21), .C1 (n_85_23), .C2 (n_79_26) );
AOI211_X1 g_100_18 (.ZN (n_100_18), .A (n_96_20), .B (n_91_20), .C1 (n_87_22), .C2 (n_81_25) );
AOI211_X1 g_102_17 (.ZN (n_102_17), .A (n_98_19), .B (n_93_19), .C1 (n_89_21), .C2 (n_83_24) );
AOI211_X1 g_103_19 (.ZN (n_103_19), .A (n_100_18), .B (n_94_21), .C1 (n_91_20), .C2 (n_85_23) );
AOI211_X1 g_104_17 (.ZN (n_104_17), .A (n_102_17), .B (n_96_20), .C1 (n_93_19), .C2 (n_87_22) );
AOI211_X1 g_102_18 (.ZN (n_102_18), .A (n_103_19), .B (n_98_19), .C1 (n_94_21), .C2 (n_89_21) );
AOI211_X1 g_103_16 (.ZN (n_103_16), .A (n_104_17), .B (n_100_18), .C1 (n_96_20), .C2 (n_91_20) );
AOI211_X1 g_101_17 (.ZN (n_101_17), .A (n_102_18), .B (n_102_17), .C1 (n_98_19), .C2 (n_93_19) );
AOI211_X1 g_99_18 (.ZN (n_99_18), .A (n_103_16), .B (n_103_19), .C1 (n_100_18), .C2 (n_94_21) );
AOI211_X1 g_97_19 (.ZN (n_97_19), .A (n_101_17), .B (n_104_17), .C1 (n_102_17), .C2 (n_96_20) );
AOI211_X1 g_95_20 (.ZN (n_95_20), .A (n_99_18), .B (n_102_18), .C1 (n_103_19), .C2 (n_98_19) );
AOI211_X1 g_94_18 (.ZN (n_94_18), .A (n_97_19), .B (n_103_16), .C1 (n_104_17), .C2 (n_100_18) );
AOI211_X1 g_92_19 (.ZN (n_92_19), .A (n_95_20), .B (n_101_17), .C1 (n_102_18), .C2 (n_102_17) );
AOI211_X1 g_90_20 (.ZN (n_90_20), .A (n_94_18), .B (n_99_18), .C1 (n_103_16), .C2 (n_103_19) );
AOI211_X1 g_88_21 (.ZN (n_88_21), .A (n_92_19), .B (n_97_19), .C1 (n_101_17), .C2 (n_104_17) );
AOI211_X1 g_86_22 (.ZN (n_86_22), .A (n_90_20), .B (n_95_20), .C1 (n_99_18), .C2 (n_102_18) );
AOI211_X1 g_85_24 (.ZN (n_85_24), .A (n_88_21), .B (n_94_18), .C1 (n_97_19), .C2 (n_103_16) );
AOI211_X1 g_83_25 (.ZN (n_83_25), .A (n_86_22), .B (n_92_19), .C1 (n_95_20), .C2 (n_101_17) );
AOI211_X1 g_82_27 (.ZN (n_82_27), .A (n_85_24), .B (n_90_20), .C1 (n_94_18), .C2 (n_99_18) );
AOI211_X1 g_84_26 (.ZN (n_84_26), .A (n_83_25), .B (n_88_21), .C1 (n_92_19), .C2 (n_97_19) );
AOI211_X1 g_86_25 (.ZN (n_86_25), .A (n_82_27), .B (n_86_22), .C1 (n_90_20), .C2 (n_95_20) );
AOI211_X1 g_87_23 (.ZN (n_87_23), .A (n_84_26), .B (n_85_24), .C1 (n_88_21), .C2 (n_94_18) );
AOI211_X1 g_89_22 (.ZN (n_89_22), .A (n_86_25), .B (n_83_25), .C1 (n_86_22), .C2 (n_92_19) );
AOI211_X1 g_91_21 (.ZN (n_91_21), .A (n_87_23), .B (n_82_27), .C1 (n_85_24), .C2 (n_90_20) );
AOI211_X1 g_93_20 (.ZN (n_93_20), .A (n_89_22), .B (n_84_26), .C1 (n_83_25), .C2 (n_88_21) );
AOI211_X1 g_92_22 (.ZN (n_92_22), .A (n_91_21), .B (n_86_25), .C1 (n_82_27), .C2 (n_86_22) );
AOI211_X1 g_90_23 (.ZN (n_90_23), .A (n_93_20), .B (n_87_23), .C1 (n_84_26), .C2 (n_85_24) );
AOI211_X1 g_88_24 (.ZN (n_88_24), .A (n_92_22), .B (n_89_22), .C1 (n_86_25), .C2 (n_83_25) );
AOI211_X1 g_87_26 (.ZN (n_87_26), .A (n_90_23), .B (n_91_21), .C1 (n_87_23), .C2 (n_82_27) );
AOI211_X1 g_86_24 (.ZN (n_86_24), .A (n_88_24), .B (n_93_20), .C1 (n_89_22), .C2 (n_84_26) );
AOI211_X1 g_88_23 (.ZN (n_88_23), .A (n_87_26), .B (n_92_22), .C1 (n_91_21), .C2 (n_86_25) );
AOI211_X1 g_90_22 (.ZN (n_90_22), .A (n_86_24), .B (n_90_23), .C1 (n_93_20), .C2 (n_87_23) );
AOI211_X1 g_92_21 (.ZN (n_92_21), .A (n_88_23), .B (n_88_24), .C1 (n_92_22), .C2 (n_89_22) );
AOI211_X1 g_94_20 (.ZN (n_94_20), .A (n_90_22), .B (n_87_26), .C1 (n_90_23), .C2 (n_91_21) );
AOI211_X1 g_96_19 (.ZN (n_96_19), .A (n_92_21), .B (n_86_24), .C1 (n_88_24), .C2 (n_93_20) );
AOI211_X1 g_95_21 (.ZN (n_95_21), .A (n_94_20), .B (n_88_23), .C1 (n_87_26), .C2 (n_92_22) );
AOI211_X1 g_93_22 (.ZN (n_93_22), .A (n_96_19), .B (n_90_22), .C1 (n_86_24), .C2 (n_90_23) );
AOI211_X1 g_91_23 (.ZN (n_91_23), .A (n_95_21), .B (n_92_21), .C1 (n_88_23), .C2 (n_88_24) );
AOI211_X1 g_89_24 (.ZN (n_89_24), .A (n_93_22), .B (n_94_20), .C1 (n_90_22), .C2 (n_87_26) );
AOI211_X1 g_87_25 (.ZN (n_87_25), .A (n_91_23), .B (n_96_19), .C1 (n_92_21), .C2 (n_86_24) );
AOI211_X1 g_85_26 (.ZN (n_85_26), .A (n_89_24), .B (n_95_21), .C1 (n_94_20), .C2 (n_88_23) );
AOI211_X1 g_83_27 (.ZN (n_83_27), .A (n_87_25), .B (n_93_22), .C1 (n_96_19), .C2 (n_90_22) );
AOI211_X1 g_84_25 (.ZN (n_84_25), .A (n_85_26), .B (n_91_23), .C1 (n_95_21), .C2 (n_92_21) );
AOI211_X1 g_82_26 (.ZN (n_82_26), .A (n_83_27), .B (n_89_24), .C1 (n_93_22), .C2 (n_94_20) );
AOI211_X1 g_80_27 (.ZN (n_80_27), .A (n_84_25), .B (n_87_25), .C1 (n_91_23), .C2 (n_96_19) );
AOI211_X1 g_78_28 (.ZN (n_78_28), .A (n_82_26), .B (n_85_26), .C1 (n_89_24), .C2 (n_95_21) );
AOI211_X1 g_77_26 (.ZN (n_77_26), .A (n_80_27), .B (n_83_27), .C1 (n_87_25), .C2 (n_93_22) );
AOI211_X1 g_75_27 (.ZN (n_75_27), .A (n_78_28), .B (n_84_25), .C1 (n_85_26), .C2 (n_91_23) );
AOI211_X1 g_73_28 (.ZN (n_73_28), .A (n_77_26), .B (n_82_26), .C1 (n_83_27), .C2 (n_89_24) );
AOI211_X1 g_71_29 (.ZN (n_71_29), .A (n_75_27), .B (n_80_27), .C1 (n_84_25), .C2 (n_87_25) );
AOI211_X1 g_69_30 (.ZN (n_69_30), .A (n_73_28), .B (n_78_28), .C1 (n_82_26), .C2 (n_85_26) );
AOI211_X1 g_67_31 (.ZN (n_67_31), .A (n_71_29), .B (n_77_26), .C1 (n_80_27), .C2 (n_83_27) );
AOI211_X1 g_68_29 (.ZN (n_68_29), .A (n_69_30), .B (n_75_27), .C1 (n_78_28), .C2 (n_84_25) );
AOI211_X1 g_66_30 (.ZN (n_66_30), .A (n_67_31), .B (n_73_28), .C1 (n_77_26), .C2 (n_82_26) );
AOI211_X1 g_64_31 (.ZN (n_64_31), .A (n_68_29), .B (n_71_29), .C1 (n_75_27), .C2 (n_80_27) );
AOI211_X1 g_62_32 (.ZN (n_62_32), .A (n_66_30), .B (n_69_30), .C1 (n_73_28), .C2 (n_78_28) );
AOI211_X1 g_60_33 (.ZN (n_60_33), .A (n_64_31), .B (n_67_31), .C1 (n_71_29), .C2 (n_77_26) );
AOI211_X1 g_58_34 (.ZN (n_58_34), .A (n_62_32), .B (n_68_29), .C1 (n_69_30), .C2 (n_75_27) );
AOI211_X1 g_56_35 (.ZN (n_56_35), .A (n_60_33), .B (n_66_30), .C1 (n_67_31), .C2 (n_73_28) );
AOI211_X1 g_54_36 (.ZN (n_54_36), .A (n_58_34), .B (n_64_31), .C1 (n_68_29), .C2 (n_71_29) );
AOI211_X1 g_52_37 (.ZN (n_52_37), .A (n_56_35), .B (n_62_32), .C1 (n_66_30), .C2 (n_69_30) );
AOI211_X1 g_50_38 (.ZN (n_50_38), .A (n_54_36), .B (n_60_33), .C1 (n_64_31), .C2 (n_67_31) );
AOI211_X1 g_48_39 (.ZN (n_48_39), .A (n_52_37), .B (n_58_34), .C1 (n_62_32), .C2 (n_68_29) );
AOI211_X1 g_46_40 (.ZN (n_46_40), .A (n_50_38), .B (n_56_35), .C1 (n_60_33), .C2 (n_66_30) );
AOI211_X1 g_44_41 (.ZN (n_44_41), .A (n_48_39), .B (n_54_36), .C1 (n_58_34), .C2 (n_64_31) );
AOI211_X1 g_42_42 (.ZN (n_42_42), .A (n_46_40), .B (n_52_37), .C1 (n_56_35), .C2 (n_62_32) );
AOI211_X1 g_43_40 (.ZN (n_43_40), .A (n_44_41), .B (n_50_38), .C1 (n_54_36), .C2 (n_60_33) );
AOI211_X1 g_41_41 (.ZN (n_41_41), .A (n_42_42), .B (n_48_39), .C1 (n_52_37), .C2 (n_58_34) );
AOI211_X1 g_39_42 (.ZN (n_39_42), .A (n_43_40), .B (n_46_40), .C1 (n_50_38), .C2 (n_56_35) );
AOI211_X1 g_37_43 (.ZN (n_37_43), .A (n_41_41), .B (n_44_41), .C1 (n_48_39), .C2 (n_54_36) );
AOI211_X1 g_35_44 (.ZN (n_35_44), .A (n_39_42), .B (n_42_42), .C1 (n_46_40), .C2 (n_52_37) );
AOI211_X1 g_34_46 (.ZN (n_34_46), .A (n_37_43), .B (n_43_40), .C1 (n_44_41), .C2 (n_50_38) );
AOI211_X1 g_32_45 (.ZN (n_32_45), .A (n_35_44), .B (n_41_41), .C1 (n_42_42), .C2 (n_48_39) );
AOI211_X1 g_34_44 (.ZN (n_34_44), .A (n_34_46), .B (n_39_42), .C1 (n_43_40), .C2 (n_46_40) );
AOI211_X1 g_36_43 (.ZN (n_36_43), .A (n_32_45), .B (n_37_43), .C1 (n_41_41), .C2 (n_44_41) );
AOI211_X1 g_35_45 (.ZN (n_35_45), .A (n_34_44), .B (n_35_44), .C1 (n_39_42), .C2 (n_42_42) );
AOI211_X1 g_37_44 (.ZN (n_37_44), .A (n_36_43), .B (n_34_46), .C1 (n_37_43), .C2 (n_43_40) );
AOI211_X1 g_39_43 (.ZN (n_39_43), .A (n_35_45), .B (n_32_45), .C1 (n_35_44), .C2 (n_41_41) );
AOI211_X1 g_41_42 (.ZN (n_41_42), .A (n_37_44), .B (n_34_44), .C1 (n_34_46), .C2 (n_39_42) );
AOI211_X1 g_43_41 (.ZN (n_43_41), .A (n_39_43), .B (n_36_43), .C1 (n_32_45), .C2 (n_37_43) );
AOI211_X1 g_45_40 (.ZN (n_45_40), .A (n_41_42), .B (n_35_45), .C1 (n_34_44), .C2 (n_35_44) );
AOI211_X1 g_47_39 (.ZN (n_47_39), .A (n_43_41), .B (n_37_44), .C1 (n_36_43), .C2 (n_34_46) );
AOI211_X1 g_49_38 (.ZN (n_49_38), .A (n_45_40), .B (n_39_43), .C1 (n_35_45), .C2 (n_32_45) );
AOI211_X1 g_51_37 (.ZN (n_51_37), .A (n_47_39), .B (n_41_42), .C1 (n_37_44), .C2 (n_34_44) );
AOI211_X1 g_53_36 (.ZN (n_53_36), .A (n_49_38), .B (n_43_41), .C1 (n_39_43), .C2 (n_36_43) );
AOI211_X1 g_52_38 (.ZN (n_52_38), .A (n_51_37), .B (n_45_40), .C1 (n_41_42), .C2 (n_35_45) );
AOI211_X1 g_54_37 (.ZN (n_54_37), .A (n_53_36), .B (n_47_39), .C1 (n_43_41), .C2 (n_37_44) );
AOI211_X1 g_56_36 (.ZN (n_56_36), .A (n_52_38), .B (n_49_38), .C1 (n_45_40), .C2 (n_39_43) );
AOI211_X1 g_58_35 (.ZN (n_58_35), .A (n_54_37), .B (n_51_37), .C1 (n_47_39), .C2 (n_41_42) );
AOI211_X1 g_60_34 (.ZN (n_60_34), .A (n_56_36), .B (n_53_36), .C1 (n_49_38), .C2 (n_43_41) );
AOI211_X1 g_62_33 (.ZN (n_62_33), .A (n_58_35), .B (n_52_38), .C1 (n_51_37), .C2 (n_45_40) );
AOI211_X1 g_64_32 (.ZN (n_64_32), .A (n_60_34), .B (n_54_37), .C1 (n_53_36), .C2 (n_47_39) );
AOI211_X1 g_66_31 (.ZN (n_66_31), .A (n_62_33), .B (n_56_36), .C1 (n_52_38), .C2 (n_49_38) );
AOI211_X1 g_68_30 (.ZN (n_68_30), .A (n_64_32), .B (n_58_35), .C1 (n_54_37), .C2 (n_51_37) );
AOI211_X1 g_67_32 (.ZN (n_67_32), .A (n_66_31), .B (n_60_34), .C1 (n_56_36), .C2 (n_53_36) );
AOI211_X1 g_69_31 (.ZN (n_69_31), .A (n_68_30), .B (n_62_33), .C1 (n_58_35), .C2 (n_52_38) );
AOI211_X1 g_68_33 (.ZN (n_68_33), .A (n_67_32), .B (n_64_32), .C1 (n_60_34), .C2 (n_54_37) );
AOI211_X1 g_66_32 (.ZN (n_66_32), .A (n_69_31), .B (n_66_31), .C1 (n_62_33), .C2 (n_56_36) );
AOI211_X1 g_68_31 (.ZN (n_68_31), .A (n_68_33), .B (n_68_30), .C1 (n_64_32), .C2 (n_58_35) );
AOI211_X1 g_70_30 (.ZN (n_70_30), .A (n_66_32), .B (n_67_32), .C1 (n_66_31), .C2 (n_60_34) );
AOI211_X1 g_72_29 (.ZN (n_72_29), .A (n_68_31), .B (n_69_31), .C1 (n_68_30), .C2 (n_62_33) );
AOI211_X1 g_74_28 (.ZN (n_74_28), .A (n_70_30), .B (n_68_33), .C1 (n_67_32), .C2 (n_64_32) );
AOI211_X1 g_76_27 (.ZN (n_76_27), .A (n_72_29), .B (n_66_32), .C1 (n_69_31), .C2 (n_66_31) );
AOI211_X1 g_75_29 (.ZN (n_75_29), .A (n_74_28), .B (n_68_31), .C1 (n_68_33), .C2 (n_68_30) );
AOI211_X1 g_77_28 (.ZN (n_77_28), .A (n_76_27), .B (n_70_30), .C1 (n_66_32), .C2 (n_67_32) );
AOI211_X1 g_79_27 (.ZN (n_79_27), .A (n_75_29), .B (n_72_29), .C1 (n_68_31), .C2 (n_69_31) );
AOI211_X1 g_81_28 (.ZN (n_81_28), .A (n_77_28), .B (n_74_28), .C1 (n_70_30), .C2 (n_68_33) );
AOI211_X1 g_79_29 (.ZN (n_79_29), .A (n_79_27), .B (n_76_27), .C1 (n_72_29), .C2 (n_66_32) );
AOI211_X1 g_78_27 (.ZN (n_78_27), .A (n_81_28), .B (n_75_29), .C1 (n_74_28), .C2 (n_68_31) );
AOI211_X1 g_76_28 (.ZN (n_76_28), .A (n_79_29), .B (n_77_28), .C1 (n_76_27), .C2 (n_70_30) );
AOI211_X1 g_74_29 (.ZN (n_74_29), .A (n_78_27), .B (n_79_27), .C1 (n_75_29), .C2 (n_72_29) );
AOI211_X1 g_72_30 (.ZN (n_72_30), .A (n_76_28), .B (n_81_28), .C1 (n_77_28), .C2 (n_74_28) );
AOI211_X1 g_70_31 (.ZN (n_70_31), .A (n_74_29), .B (n_79_29), .C1 (n_79_27), .C2 (n_76_27) );
AOI211_X1 g_68_32 (.ZN (n_68_32), .A (n_72_30), .B (n_78_27), .C1 (n_81_28), .C2 (n_75_29) );
AOI211_X1 g_66_33 (.ZN (n_66_33), .A (n_70_31), .B (n_76_28), .C1 (n_79_29), .C2 (n_77_28) );
AOI211_X1 g_64_34 (.ZN (n_64_34), .A (n_68_32), .B (n_74_29), .C1 (n_78_27), .C2 (n_79_27) );
AOI211_X1 g_65_32 (.ZN (n_65_32), .A (n_66_33), .B (n_72_30), .C1 (n_76_28), .C2 (n_81_28) );
AOI211_X1 g_63_33 (.ZN (n_63_33), .A (n_64_34), .B (n_70_31), .C1 (n_74_29), .C2 (n_79_29) );
AOI211_X1 g_61_34 (.ZN (n_61_34), .A (n_65_32), .B (n_68_32), .C1 (n_72_30), .C2 (n_78_27) );
AOI211_X1 g_59_35 (.ZN (n_59_35), .A (n_63_33), .B (n_66_33), .C1 (n_70_31), .C2 (n_76_28) );
AOI211_X1 g_57_36 (.ZN (n_57_36), .A (n_61_34), .B (n_64_34), .C1 (n_68_32), .C2 (n_74_29) );
AOI211_X1 g_55_37 (.ZN (n_55_37), .A (n_59_35), .B (n_65_32), .C1 (n_66_33), .C2 (n_72_30) );
AOI211_X1 g_53_38 (.ZN (n_53_38), .A (n_57_36), .B (n_63_33), .C1 (n_64_34), .C2 (n_70_31) );
AOI211_X1 g_51_39 (.ZN (n_51_39), .A (n_55_37), .B (n_61_34), .C1 (n_65_32), .C2 (n_68_32) );
AOI211_X1 g_49_40 (.ZN (n_49_40), .A (n_53_38), .B (n_59_35), .C1 (n_63_33), .C2 (n_66_33) );
AOI211_X1 g_47_41 (.ZN (n_47_41), .A (n_51_39), .B (n_57_36), .C1 (n_61_34), .C2 (n_64_34) );
AOI211_X1 g_45_42 (.ZN (n_45_42), .A (n_49_40), .B (n_55_37), .C1 (n_59_35), .C2 (n_65_32) );
AOI211_X1 g_43_43 (.ZN (n_43_43), .A (n_47_41), .B (n_53_38), .C1 (n_57_36), .C2 (n_63_33) );
AOI211_X1 g_41_44 (.ZN (n_41_44), .A (n_45_42), .B (n_51_39), .C1 (n_55_37), .C2 (n_61_34) );
AOI211_X1 g_39_45 (.ZN (n_39_45), .A (n_43_43), .B (n_49_40), .C1 (n_53_38), .C2 (n_59_35) );
AOI211_X1 g_40_43 (.ZN (n_40_43), .A (n_41_44), .B (n_47_41), .C1 (n_51_39), .C2 (n_57_36) );
AOI211_X1 g_38_44 (.ZN (n_38_44), .A (n_39_45), .B (n_45_42), .C1 (n_49_40), .C2 (n_55_37) );
AOI211_X1 g_36_45 (.ZN (n_36_45), .A (n_40_43), .B (n_43_43), .C1 (n_47_41), .C2 (n_53_38) );
AOI211_X1 g_38_46 (.ZN (n_38_46), .A (n_38_44), .B (n_41_44), .C1 (n_45_42), .C2 (n_51_39) );
AOI211_X1 g_39_44 (.ZN (n_39_44), .A (n_36_45), .B (n_39_45), .C1 (n_43_43), .C2 (n_49_40) );
AOI211_X1 g_41_43 (.ZN (n_41_43), .A (n_38_46), .B (n_40_43), .C1 (n_41_44), .C2 (n_47_41) );
AOI211_X1 g_43_42 (.ZN (n_43_42), .A (n_39_44), .B (n_38_44), .C1 (n_39_45), .C2 (n_45_42) );
AOI211_X1 g_45_41 (.ZN (n_45_41), .A (n_41_43), .B (n_36_45), .C1 (n_40_43), .C2 (n_43_43) );
AOI211_X1 g_44_43 (.ZN (n_44_43), .A (n_43_42), .B (n_38_46), .C1 (n_38_44), .C2 (n_41_44) );
AOI211_X1 g_46_42 (.ZN (n_46_42), .A (n_45_41), .B (n_39_44), .C1 (n_36_45), .C2 (n_39_45) );
AOI211_X1 g_48_41 (.ZN (n_48_41), .A (n_44_43), .B (n_41_43), .C1 (n_38_46), .C2 (n_40_43) );
AOI211_X1 g_50_40 (.ZN (n_50_40), .A (n_46_42), .B (n_43_42), .C1 (n_39_44), .C2 (n_38_44) );
AOI211_X1 g_52_39 (.ZN (n_52_39), .A (n_48_41), .B (n_45_41), .C1 (n_41_43), .C2 (n_36_45) );
AOI211_X1 g_54_38 (.ZN (n_54_38), .A (n_50_40), .B (n_44_43), .C1 (n_43_42), .C2 (n_38_46) );
AOI211_X1 g_56_37 (.ZN (n_56_37), .A (n_52_39), .B (n_46_42), .C1 (n_45_41), .C2 (n_39_44) );
AOI211_X1 g_58_36 (.ZN (n_58_36), .A (n_54_38), .B (n_48_41), .C1 (n_44_43), .C2 (n_41_43) );
AOI211_X1 g_60_35 (.ZN (n_60_35), .A (n_56_37), .B (n_50_40), .C1 (n_46_42), .C2 (n_43_42) );
AOI211_X1 g_62_34 (.ZN (n_62_34), .A (n_58_36), .B (n_52_39), .C1 (n_48_41), .C2 (n_45_41) );
AOI211_X1 g_64_33 (.ZN (n_64_33), .A (n_60_35), .B (n_54_38), .C1 (n_50_40), .C2 (n_44_43) );
AOI211_X1 g_66_34 (.ZN (n_66_34), .A (n_62_34), .B (n_56_37), .C1 (n_52_39), .C2 (n_46_42) );
AOI211_X1 g_64_35 (.ZN (n_64_35), .A (n_64_33), .B (n_58_36), .C1 (n_54_38), .C2 (n_48_41) );
AOI211_X1 g_65_33 (.ZN (n_65_33), .A (n_66_34), .B (n_60_35), .C1 (n_56_37), .C2 (n_50_40) );
AOI211_X1 g_63_34 (.ZN (n_63_34), .A (n_64_35), .B (n_62_34), .C1 (n_58_36), .C2 (n_52_39) );
AOI211_X1 g_61_35 (.ZN (n_61_35), .A (n_65_33), .B (n_64_33), .C1 (n_60_35), .C2 (n_54_38) );
AOI211_X1 g_59_36 (.ZN (n_59_36), .A (n_63_34), .B (n_66_34), .C1 (n_62_34), .C2 (n_56_37) );
AOI211_X1 g_57_37 (.ZN (n_57_37), .A (n_61_35), .B (n_64_35), .C1 (n_64_33), .C2 (n_58_36) );
AOI211_X1 g_55_38 (.ZN (n_55_38), .A (n_59_36), .B (n_65_33), .C1 (n_66_34), .C2 (n_60_35) );
AOI211_X1 g_53_39 (.ZN (n_53_39), .A (n_57_37), .B (n_63_34), .C1 (n_64_35), .C2 (n_62_34) );
AOI211_X1 g_51_40 (.ZN (n_51_40), .A (n_55_38), .B (n_61_35), .C1 (n_65_33), .C2 (n_64_33) );
AOI211_X1 g_49_41 (.ZN (n_49_41), .A (n_53_39), .B (n_59_36), .C1 (n_63_34), .C2 (n_66_34) );
AOI211_X1 g_50_39 (.ZN (n_50_39), .A (n_51_40), .B (n_57_37), .C1 (n_61_35), .C2 (n_64_35) );
AOI211_X1 g_48_40 (.ZN (n_48_40), .A (n_49_41), .B (n_55_38), .C1 (n_59_36), .C2 (n_65_33) );
AOI211_X1 g_46_41 (.ZN (n_46_41), .A (n_50_39), .B (n_53_39), .C1 (n_57_37), .C2 (n_63_34) );
AOI211_X1 g_44_42 (.ZN (n_44_42), .A (n_48_40), .B (n_51_40), .C1 (n_55_38), .C2 (n_61_35) );
AOI211_X1 g_42_43 (.ZN (n_42_43), .A (n_46_41), .B (n_49_41), .C1 (n_53_39), .C2 (n_59_36) );
AOI211_X1 g_40_44 (.ZN (n_40_44), .A (n_44_42), .B (n_50_39), .C1 (n_51_40), .C2 (n_57_37) );
AOI211_X1 g_38_45 (.ZN (n_38_45), .A (n_42_43), .B (n_48_40), .C1 (n_49_41), .C2 (n_55_38) );
AOI211_X1 g_36_44 (.ZN (n_36_44), .A (n_40_44), .B (n_46_41), .C1 (n_50_39), .C2 (n_53_39) );
AOI211_X1 g_34_45 (.ZN (n_34_45), .A (n_38_45), .B (n_44_42), .C1 (n_48_40), .C2 (n_51_40) );
AOI211_X1 g_32_46 (.ZN (n_32_46), .A (n_36_44), .B (n_42_43), .C1 (n_46_41), .C2 (n_49_41) );
AOI211_X1 g_30_47 (.ZN (n_30_47), .A (n_34_45), .B (n_40_44), .C1 (n_44_42), .C2 (n_50_39) );
AOI211_X1 g_28_48 (.ZN (n_28_48), .A (n_32_46), .B (n_38_45), .C1 (n_42_43), .C2 (n_48_40) );
AOI211_X1 g_26_49 (.ZN (n_26_49), .A (n_30_47), .B (n_36_44), .C1 (n_40_44), .C2 (n_46_41) );
AOI211_X1 g_24_50 (.ZN (n_24_50), .A (n_28_48), .B (n_34_45), .C1 (n_38_45), .C2 (n_44_42) );
AOI211_X1 g_25_48 (.ZN (n_25_48), .A (n_26_49), .B (n_32_46), .C1 (n_36_44), .C2 (n_42_43) );
AOI211_X1 g_23_47 (.ZN (n_23_47), .A (n_24_50), .B (n_30_47), .C1 (n_34_45), .C2 (n_40_44) );
AOI211_X1 g_21_48 (.ZN (n_21_48), .A (n_25_48), .B (n_28_48), .C1 (n_32_46), .C2 (n_38_45) );
AOI211_X1 g_19_49 (.ZN (n_19_49), .A (n_23_47), .B (n_26_49), .C1 (n_30_47), .C2 (n_36_44) );
AOI211_X1 g_17_50 (.ZN (n_17_50), .A (n_21_48), .B (n_24_50), .C1 (n_28_48), .C2 (n_34_45) );
AOI211_X1 g_15_51 (.ZN (n_15_51), .A (n_19_49), .B (n_25_48), .C1 (n_26_49), .C2 (n_32_46) );
AOI211_X1 g_13_52 (.ZN (n_13_52), .A (n_17_50), .B (n_23_47), .C1 (n_24_50), .C2 (n_30_47) );
AOI211_X1 g_11_53 (.ZN (n_11_53), .A (n_15_51), .B (n_21_48), .C1 (n_25_48), .C2 (n_28_48) );
AOI211_X1 g_9_54 (.ZN (n_9_54), .A (n_13_52), .B (n_19_49), .C1 (n_23_47), .C2 (n_26_49) );
AOI211_X1 g_7_55 (.ZN (n_7_55), .A (n_11_53), .B (n_17_50), .C1 (n_21_48), .C2 (n_24_50) );
AOI211_X1 g_6_53 (.ZN (n_6_53), .A (n_9_54), .B (n_15_51), .C1 (n_19_49), .C2 (n_25_48) );
AOI211_X1 g_4_54 (.ZN (n_4_54), .A (n_7_55), .B (n_13_52), .C1 (n_17_50), .C2 (n_23_47) );
AOI211_X1 g_3_56 (.ZN (n_3_56), .A (n_6_53), .B (n_11_53), .C1 (n_15_51), .C2 (n_21_48) );
AOI211_X1 g_5_55 (.ZN (n_5_55), .A (n_4_54), .B (n_9_54), .C1 (n_13_52), .C2 (n_19_49) );
AOI211_X1 g_6_57 (.ZN (n_6_57), .A (n_3_56), .B (n_7_55), .C1 (n_11_53), .C2 (n_17_50) );
AOI211_X1 g_4_58 (.ZN (n_4_58), .A (n_5_55), .B (n_6_53), .C1 (n_9_54), .C2 (n_15_51) );
AOI211_X1 g_5_56 (.ZN (n_5_56), .A (n_6_57), .B (n_4_54), .C1 (n_7_55), .C2 (n_13_52) );
AOI211_X1 g_7_57 (.ZN (n_7_57), .A (n_4_58), .B (n_3_56), .C1 (n_6_53), .C2 (n_11_53) );
AOI211_X1 g_6_55 (.ZN (n_6_55), .A (n_5_56), .B (n_5_55), .C1 (n_4_54), .C2 (n_9_54) );
AOI211_X1 g_5_57 (.ZN (n_5_57), .A (n_7_57), .B (n_6_57), .C1 (n_3_56), .C2 (n_7_55) );
AOI211_X1 g_7_56 (.ZN (n_7_56), .A (n_6_55), .B (n_4_58), .C1 (n_5_55), .C2 (n_6_53) );
AOI211_X1 g_9_55 (.ZN (n_9_55), .A (n_5_57), .B (n_5_56), .C1 (n_6_57), .C2 (n_4_54) );
AOI211_X1 g_10_53 (.ZN (n_10_53), .A (n_7_56), .B (n_7_57), .C1 (n_4_58), .C2 (n_3_56) );
AOI211_X1 g_12_52 (.ZN (n_12_52), .A (n_9_55), .B (n_6_55), .C1 (n_5_56), .C2 (n_5_55) );
AOI211_X1 g_14_51 (.ZN (n_14_51), .A (n_10_53), .B (n_5_57), .C1 (n_7_57), .C2 (n_6_57) );
AOI211_X1 g_16_50 (.ZN (n_16_50), .A (n_12_52), .B (n_7_56), .C1 (n_6_55), .C2 (n_4_58) );
AOI211_X1 g_18_49 (.ZN (n_18_49), .A (n_14_51), .B (n_9_55), .C1 (n_5_57), .C2 (n_5_56) );
AOI211_X1 g_20_48 (.ZN (n_20_48), .A (n_16_50), .B (n_10_53), .C1 (n_7_56), .C2 (n_7_57) );
AOI211_X1 g_22_49 (.ZN (n_22_49), .A (n_18_49), .B (n_12_52), .C1 (n_9_55), .C2 (n_6_55) );
AOI211_X1 g_20_50 (.ZN (n_20_50), .A (n_20_48), .B (n_14_51), .C1 (n_10_53), .C2 (n_5_57) );
AOI211_X1 g_18_51 (.ZN (n_18_51), .A (n_22_49), .B (n_16_50), .C1 (n_12_52), .C2 (n_7_56) );
AOI211_X1 g_16_52 (.ZN (n_16_52), .A (n_20_50), .B (n_18_49), .C1 (n_14_51), .C2 (n_9_55) );
AOI211_X1 g_14_53 (.ZN (n_14_53), .A (n_18_51), .B (n_20_48), .C1 (n_16_50), .C2 (n_10_53) );
AOI211_X1 g_12_54 (.ZN (n_12_54), .A (n_16_52), .B (n_22_49), .C1 (n_18_49), .C2 (n_12_52) );
AOI211_X1 g_10_55 (.ZN (n_10_55), .A (n_14_53), .B (n_20_50), .C1 (n_20_48), .C2 (n_14_51) );
AOI211_X1 g_8_56 (.ZN (n_8_56), .A (n_12_54), .B (n_18_51), .C1 (n_22_49), .C2 (n_16_50) );
AOI211_X1 g_7_58 (.ZN (n_7_58), .A (n_10_55), .B (n_16_52), .C1 (n_20_50), .C2 (n_18_49) );
AOI211_X1 g_9_57 (.ZN (n_9_57), .A (n_8_56), .B (n_14_53), .C1 (n_18_51), .C2 (n_20_48) );
AOI211_X1 g_11_56 (.ZN (n_11_56), .A (n_7_58), .B (n_12_54), .C1 (n_16_52), .C2 (n_22_49) );
AOI211_X1 g_13_55 (.ZN (n_13_55), .A (n_9_57), .B (n_10_55), .C1 (n_14_53), .C2 (n_20_50) );
AOI211_X1 g_11_54 (.ZN (n_11_54), .A (n_11_56), .B (n_8_56), .C1 (n_12_54), .C2 (n_18_51) );
AOI211_X1 g_13_53 (.ZN (n_13_53), .A (n_13_55), .B (n_7_58), .C1 (n_10_55), .C2 (n_16_52) );
AOI211_X1 g_15_52 (.ZN (n_15_52), .A (n_11_54), .B (n_9_57), .C1 (n_8_56), .C2 (n_14_53) );
AOI211_X1 g_17_51 (.ZN (n_17_51), .A (n_13_53), .B (n_11_56), .C1 (n_7_58), .C2 (n_12_54) );
AOI211_X1 g_19_50 (.ZN (n_19_50), .A (n_15_52), .B (n_13_55), .C1 (n_9_57), .C2 (n_10_55) );
AOI211_X1 g_21_51 (.ZN (n_21_51), .A (n_17_51), .B (n_11_54), .C1 (n_11_56), .C2 (n_8_56) );
AOI211_X1 g_19_52 (.ZN (n_19_52), .A (n_19_50), .B (n_13_53), .C1 (n_13_55), .C2 (n_7_58) );
AOI211_X1 g_17_53 (.ZN (n_17_53), .A (n_21_51), .B (n_15_52), .C1 (n_11_54), .C2 (n_9_57) );
AOI211_X1 g_15_54 (.ZN (n_15_54), .A (n_19_52), .B (n_17_51), .C1 (n_13_53), .C2 (n_11_56) );
AOI211_X1 g_14_56 (.ZN (n_14_56), .A (n_17_53), .B (n_19_50), .C1 (n_15_52), .C2 (n_13_55) );
AOI211_X1 g_13_54 (.ZN (n_13_54), .A (n_15_54), .B (n_21_51), .C1 (n_17_51), .C2 (n_11_54) );
AOI211_X1 g_15_53 (.ZN (n_15_53), .A (n_14_56), .B (n_19_52), .C1 (n_19_50), .C2 (n_13_53) );
AOI211_X1 g_17_52 (.ZN (n_17_52), .A (n_13_54), .B (n_17_53), .C1 (n_21_51), .C2 (n_15_52) );
AOI211_X1 g_19_51 (.ZN (n_19_51), .A (n_15_53), .B (n_15_54), .C1 (n_19_52), .C2 (n_17_51) );
AOI211_X1 g_21_50 (.ZN (n_21_50), .A (n_17_52), .B (n_14_56), .C1 (n_17_53), .C2 (n_19_50) );
AOI211_X1 g_23_49 (.ZN (n_23_49), .A (n_19_51), .B (n_13_54), .C1 (n_15_54), .C2 (n_21_51) );
AOI211_X1 g_22_51 (.ZN (n_22_51), .A (n_21_50), .B (n_15_53), .C1 (n_14_56), .C2 (n_19_52) );
AOI211_X1 g_20_52 (.ZN (n_20_52), .A (n_23_49), .B (n_17_52), .C1 (n_13_54), .C2 (n_17_53) );
AOI211_X1 g_18_53 (.ZN (n_18_53), .A (n_22_51), .B (n_19_51), .C1 (n_15_53), .C2 (n_15_54) );
AOI211_X1 g_16_54 (.ZN (n_16_54), .A (n_20_52), .B (n_21_50), .C1 (n_17_52), .C2 (n_14_56) );
AOI211_X1 g_14_55 (.ZN (n_14_55), .A (n_18_53), .B (n_23_49), .C1 (n_19_51), .C2 (n_13_54) );
AOI211_X1 g_12_56 (.ZN (n_12_56), .A (n_16_54), .B (n_22_51), .C1 (n_21_50), .C2 (n_15_53) );
AOI211_X1 g_10_57 (.ZN (n_10_57), .A (n_14_55), .B (n_20_52), .C1 (n_23_49), .C2 (n_17_52) );
AOI211_X1 g_11_55 (.ZN (n_11_55), .A (n_12_56), .B (n_18_53), .C1 (n_22_51), .C2 (n_19_51) );
AOI211_X1 g_9_56 (.ZN (n_9_56), .A (n_10_57), .B (n_16_54), .C1 (n_20_52), .C2 (n_21_50) );
AOI211_X1 g_8_58 (.ZN (n_8_58), .A (n_11_55), .B (n_14_55), .C1 (n_18_53), .C2 (n_23_49) );
AOI211_X1 g_6_59 (.ZN (n_6_59), .A (n_9_56), .B (n_12_56), .C1 (n_16_54), .C2 (n_22_51) );
AOI211_X1 g_5_61 (.ZN (n_5_61), .A (n_8_58), .B (n_10_57), .C1 (n_14_55), .C2 (n_20_52) );
AOI211_X1 g_4_59 (.ZN (n_4_59), .A (n_6_59), .B (n_11_55), .C1 (n_12_56), .C2 (n_18_53) );
AOI211_X1 g_3_61 (.ZN (n_3_61), .A (n_5_61), .B (n_9_56), .C1 (n_10_57), .C2 (n_16_54) );
AOI211_X1 g_5_60 (.ZN (n_5_60), .A (n_4_59), .B (n_8_58), .C1 (n_11_55), .C2 (n_14_55) );
AOI211_X1 g_6_58 (.ZN (n_6_58), .A (n_3_61), .B (n_6_59), .C1 (n_9_56), .C2 (n_12_56) );
AOI211_X1 g_8_57 (.ZN (n_8_57), .A (n_5_60), .B (n_5_61), .C1 (n_8_58), .C2 (n_10_57) );
AOI211_X1 g_10_56 (.ZN (n_10_56), .A (n_6_58), .B (n_4_59), .C1 (n_6_59), .C2 (n_11_55) );
AOI211_X1 g_12_55 (.ZN (n_12_55), .A (n_8_57), .B (n_3_61), .C1 (n_5_61), .C2 (n_9_56) );
AOI211_X1 g_14_54 (.ZN (n_14_54), .A (n_10_56), .B (n_5_60), .C1 (n_4_59), .C2 (n_8_58) );
AOI211_X1 g_16_53 (.ZN (n_16_53), .A (n_12_55), .B (n_6_58), .C1 (n_3_61), .C2 (n_6_59) );
AOI211_X1 g_18_52 (.ZN (n_18_52), .A (n_14_54), .B (n_8_57), .C1 (n_5_60), .C2 (n_5_61) );
AOI211_X1 g_20_51 (.ZN (n_20_51), .A (n_16_53), .B (n_10_56), .C1 (n_6_58), .C2 (n_4_59) );
AOI211_X1 g_22_50 (.ZN (n_22_50), .A (n_18_52), .B (n_12_55), .C1 (n_8_57), .C2 (n_3_61) );
AOI211_X1 g_24_49 (.ZN (n_24_49), .A (n_20_51), .B (n_14_54), .C1 (n_10_56), .C2 (n_5_60) );
AOI211_X1 g_26_48 (.ZN (n_26_48), .A (n_22_50), .B (n_16_53), .C1 (n_12_55), .C2 (n_6_58) );
AOI211_X1 g_28_47 (.ZN (n_28_47), .A (n_24_49), .B (n_18_52), .C1 (n_14_54), .C2 (n_8_57) );
AOI211_X1 g_30_46 (.ZN (n_30_46), .A (n_26_48), .B (n_20_51), .C1 (n_16_53), .C2 (n_10_56) );
AOI211_X1 g_32_47 (.ZN (n_32_47), .A (n_28_47), .B (n_22_50), .C1 (n_18_52), .C2 (n_12_55) );
AOI211_X1 g_30_48 (.ZN (n_30_48), .A (n_30_46), .B (n_24_49), .C1 (n_20_51), .C2 (n_14_54) );
AOI211_X1 g_29_50 (.ZN (n_29_50), .A (n_32_47), .B (n_26_48), .C1 (n_22_50), .C2 (n_16_53) );
AOI211_X1 g_27_49 (.ZN (n_27_49), .A (n_30_48), .B (n_28_47), .C1 (n_24_49), .C2 (n_18_52) );
AOI211_X1 g_29_48 (.ZN (n_29_48), .A (n_29_50), .B (n_30_46), .C1 (n_26_48), .C2 (n_20_51) );
AOI211_X1 g_31_47 (.ZN (n_31_47), .A (n_27_49), .B (n_32_47), .C1 (n_28_47), .C2 (n_22_50) );
AOI211_X1 g_33_46 (.ZN (n_33_46), .A (n_29_48), .B (n_30_48), .C1 (n_30_46), .C2 (n_24_49) );
AOI211_X1 g_32_48 (.ZN (n_32_48), .A (n_31_47), .B (n_29_50), .C1 (n_32_47), .C2 (n_26_48) );
AOI211_X1 g_34_47 (.ZN (n_34_47), .A (n_33_46), .B (n_27_49), .C1 (n_30_48), .C2 (n_28_47) );
AOI211_X1 g_36_46 (.ZN (n_36_46), .A (n_32_48), .B (n_29_48), .C1 (n_29_50), .C2 (n_30_46) );
AOI211_X1 g_35_48 (.ZN (n_35_48), .A (n_34_47), .B (n_31_47), .C1 (n_27_49), .C2 (n_32_47) );
AOI211_X1 g_33_47 (.ZN (n_33_47), .A (n_36_46), .B (n_33_46), .C1 (n_29_48), .C2 (n_30_48) );
AOI211_X1 g_35_46 (.ZN (n_35_46), .A (n_35_48), .B (n_32_48), .C1 (n_31_47), .C2 (n_29_50) );
AOI211_X1 g_37_45 (.ZN (n_37_45), .A (n_33_47), .B (n_34_47), .C1 (n_33_46), .C2 (n_27_49) );
AOI211_X1 g_36_47 (.ZN (n_36_47), .A (n_35_46), .B (n_36_46), .C1 (n_32_48), .C2 (n_29_48) );
AOI211_X1 g_34_48 (.ZN (n_34_48), .A (n_37_45), .B (n_35_48), .C1 (n_34_47), .C2 (n_31_47) );
AOI211_X1 g_32_49 (.ZN (n_32_49), .A (n_36_47), .B (n_33_47), .C1 (n_36_46), .C2 (n_33_46) );
AOI211_X1 g_30_50 (.ZN (n_30_50), .A (n_34_48), .B (n_35_46), .C1 (n_35_48), .C2 (n_32_48) );
AOI211_X1 g_31_48 (.ZN (n_31_48), .A (n_32_49), .B (n_37_45), .C1 (n_33_47), .C2 (n_34_47) );
AOI211_X1 g_29_49 (.ZN (n_29_49), .A (n_30_50), .B (n_36_47), .C1 (n_35_46), .C2 (n_36_46) );
AOI211_X1 g_27_50 (.ZN (n_27_50), .A (n_31_48), .B (n_34_48), .C1 (n_37_45), .C2 (n_35_48) );
AOI211_X1 g_25_51 (.ZN (n_25_51), .A (n_29_49), .B (n_32_49), .C1 (n_36_47), .C2 (n_33_47) );
AOI211_X1 g_23_52 (.ZN (n_23_52), .A (n_27_50), .B (n_30_50), .C1 (n_34_48), .C2 (n_35_46) );
AOI211_X1 g_21_53 (.ZN (n_21_53), .A (n_25_51), .B (n_31_48), .C1 (n_32_49), .C2 (n_37_45) );
AOI211_X1 g_19_54 (.ZN (n_19_54), .A (n_23_52), .B (n_29_49), .C1 (n_30_50), .C2 (n_36_47) );
AOI211_X1 g_17_55 (.ZN (n_17_55), .A (n_21_53), .B (n_27_50), .C1 (n_31_48), .C2 (n_34_48) );
AOI211_X1 g_15_56 (.ZN (n_15_56), .A (n_19_54), .B (n_25_51), .C1 (n_29_49), .C2 (n_32_49) );
AOI211_X1 g_13_57 (.ZN (n_13_57), .A (n_17_55), .B (n_23_52), .C1 (n_27_50), .C2 (n_30_50) );
AOI211_X1 g_11_58 (.ZN (n_11_58), .A (n_15_56), .B (n_21_53), .C1 (n_25_51), .C2 (n_31_48) );
AOI211_X1 g_9_59 (.ZN (n_9_59), .A (n_13_57), .B (n_19_54), .C1 (n_23_52), .C2 (n_29_49) );
AOI211_X1 g_7_60 (.ZN (n_7_60), .A (n_11_58), .B (n_17_55), .C1 (n_21_53), .C2 (n_27_50) );
AOI211_X1 g_5_59 (.ZN (n_5_59), .A (n_9_59), .B (n_15_56), .C1 (n_19_54), .C2 (n_25_51) );
AOI211_X1 g_3_60 (.ZN (n_3_60), .A (n_7_60), .B (n_13_57), .C1 (n_17_55), .C2 (n_23_52) );
AOI211_X1 g_2_62 (.ZN (n_2_62), .A (n_5_59), .B (n_11_58), .C1 (n_15_56), .C2 (n_21_53) );
AOI211_X1 g_1_64 (.ZN (n_1_64), .A (n_3_60), .B (n_9_59), .C1 (n_13_57), .C2 (n_19_54) );
AOI211_X1 g_3_63 (.ZN (n_3_63), .A (n_2_62), .B (n_7_60), .C1 (n_11_58), .C2 (n_17_55) );
AOI211_X1 g_4_61 (.ZN (n_4_61), .A (n_1_64), .B (n_5_59), .C1 (n_9_59), .C2 (n_15_56) );
AOI211_X1 g_6_60 (.ZN (n_6_60), .A (n_3_63), .B (n_3_60), .C1 (n_7_60), .C2 (n_13_57) );
AOI211_X1 g_5_62 (.ZN (n_5_62), .A (n_4_61), .B (n_2_62), .C1 (n_5_59), .C2 (n_11_58) );
AOI211_X1 g_7_61 (.ZN (n_7_61), .A (n_6_60), .B (n_1_64), .C1 (n_3_60), .C2 (n_9_59) );
AOI211_X1 g_8_59 (.ZN (n_8_59), .A (n_5_62), .B (n_3_63), .C1 (n_2_62), .C2 (n_7_60) );
AOI211_X1 g_10_58 (.ZN (n_10_58), .A (n_7_61), .B (n_4_61), .C1 (n_1_64), .C2 (n_5_59) );
AOI211_X1 g_12_57 (.ZN (n_12_57), .A (n_8_59), .B (n_6_60), .C1 (n_3_63), .C2 (n_3_60) );
AOI211_X1 g_11_59 (.ZN (n_11_59), .A (n_10_58), .B (n_5_62), .C1 (n_4_61), .C2 (n_2_62) );
AOI211_X1 g_9_58 (.ZN (n_9_58), .A (n_12_57), .B (n_7_61), .C1 (n_6_60), .C2 (n_1_64) );
AOI211_X1 g_7_59 (.ZN (n_7_59), .A (n_11_59), .B (n_8_59), .C1 (n_5_62), .C2 (n_3_63) );
AOI211_X1 g_9_60 (.ZN (n_9_60), .A (n_9_58), .B (n_10_58), .C1 (n_7_61), .C2 (n_4_61) );
AOI211_X1 g_8_62 (.ZN (n_8_62), .A (n_7_59), .B (n_12_57), .C1 (n_8_59), .C2 (n_6_60) );
AOI211_X1 g_6_61 (.ZN (n_6_61), .A (n_9_60), .B (n_11_59), .C1 (n_10_58), .C2 (n_5_62) );
AOI211_X1 g_4_62 (.ZN (n_4_62), .A (n_8_62), .B (n_9_58), .C1 (n_12_57), .C2 (n_7_61) );
AOI211_X1 g_6_63 (.ZN (n_6_63), .A (n_6_61), .B (n_7_59), .C1 (n_11_59), .C2 (n_8_59) );
AOI211_X1 g_5_65 (.ZN (n_5_65), .A (n_4_62), .B (n_9_60), .C1 (n_9_58), .C2 (n_10_58) );
AOI211_X1 g_4_63 (.ZN (n_4_63), .A (n_6_63), .B (n_8_62), .C1 (n_7_59), .C2 (n_12_57) );
AOI211_X1 g_3_65 (.ZN (n_3_65), .A (n_5_65), .B (n_6_61), .C1 (n_9_60), .C2 (n_11_59) );
AOI211_X1 g_5_64 (.ZN (n_5_64), .A (n_4_63), .B (n_4_62), .C1 (n_8_62), .C2 (n_9_58) );
AOI211_X1 g_6_62 (.ZN (n_6_62), .A (n_3_65), .B (n_6_63), .C1 (n_6_61), .C2 (n_7_59) );
AOI211_X1 g_8_61 (.ZN (n_8_61), .A (n_5_64), .B (n_5_65), .C1 (n_4_62), .C2 (n_9_60) );
AOI211_X1 g_10_60 (.ZN (n_10_60), .A (n_6_62), .B (n_4_63), .C1 (n_6_63), .C2 (n_8_62) );
AOI211_X1 g_12_59 (.ZN (n_12_59), .A (n_8_61), .B (n_3_65), .C1 (n_5_65), .C2 (n_6_61) );
AOI211_X1 g_11_57 (.ZN (n_11_57), .A (n_10_60), .B (n_5_64), .C1 (n_4_63), .C2 (n_4_62) );
AOI211_X1 g_13_56 (.ZN (n_13_56), .A (n_12_59), .B (n_6_62), .C1 (n_3_65), .C2 (n_6_63) );
AOI211_X1 g_15_55 (.ZN (n_15_55), .A (n_11_57), .B (n_8_61), .C1 (n_5_64), .C2 (n_5_65) );
AOI211_X1 g_17_54 (.ZN (n_17_54), .A (n_13_56), .B (n_10_60), .C1 (n_6_62), .C2 (n_4_63) );
AOI211_X1 g_19_53 (.ZN (n_19_53), .A (n_15_55), .B (n_12_59), .C1 (n_8_61), .C2 (n_3_65) );
AOI211_X1 g_21_52 (.ZN (n_21_52), .A (n_17_54), .B (n_11_57), .C1 (n_10_60), .C2 (n_5_64) );
AOI211_X1 g_23_51 (.ZN (n_23_51), .A (n_19_53), .B (n_13_56), .C1 (n_12_59), .C2 (n_6_62) );
AOI211_X1 g_25_50 (.ZN (n_25_50), .A (n_21_52), .B (n_15_55), .C1 (n_11_57), .C2 (n_8_61) );
AOI211_X1 g_27_51 (.ZN (n_27_51), .A (n_23_51), .B (n_17_54), .C1 (n_13_56), .C2 (n_10_60) );
AOI211_X1 g_25_52 (.ZN (n_25_52), .A (n_25_50), .B (n_19_53), .C1 (n_15_55), .C2 (n_12_59) );
AOI211_X1 g_26_50 (.ZN (n_26_50), .A (n_27_51), .B (n_21_52), .C1 (n_17_54), .C2 (n_11_57) );
AOI211_X1 g_24_51 (.ZN (n_24_51), .A (n_25_52), .B (n_23_51), .C1 (n_19_53), .C2 (n_13_56) );
AOI211_X1 g_22_52 (.ZN (n_22_52), .A (n_26_50), .B (n_25_50), .C1 (n_21_52), .C2 (n_15_55) );
AOI211_X1 g_20_53 (.ZN (n_20_53), .A (n_24_51), .B (n_27_51), .C1 (n_23_51), .C2 (n_17_54) );
AOI211_X1 g_18_54 (.ZN (n_18_54), .A (n_22_52), .B (n_25_52), .C1 (n_25_50), .C2 (n_19_53) );
AOI211_X1 g_16_55 (.ZN (n_16_55), .A (n_20_53), .B (n_26_50), .C1 (n_27_51), .C2 (n_21_52) );
AOI211_X1 g_15_57 (.ZN (n_15_57), .A (n_18_54), .B (n_24_51), .C1 (n_25_52), .C2 (n_23_51) );
AOI211_X1 g_13_58 (.ZN (n_13_58), .A (n_16_55), .B (n_22_52), .C1 (n_26_50), .C2 (n_25_50) );
AOI211_X1 g_12_60 (.ZN (n_12_60), .A (n_15_57), .B (n_20_53), .C1 (n_24_51), .C2 (n_27_51) );
AOI211_X1 g_10_59 (.ZN (n_10_59), .A (n_13_58), .B (n_18_54), .C1 (n_22_52), .C2 (n_25_52) );
AOI211_X1 g_8_60 (.ZN (n_8_60), .A (n_12_60), .B (n_16_55), .C1 (n_20_53), .C2 (n_26_50) );
AOI211_X1 g_10_61 (.ZN (n_10_61), .A (n_10_59), .B (n_15_57), .C1 (n_18_54), .C2 (n_24_51) );
AOI211_X1 g_9_63 (.ZN (n_9_63), .A (n_8_60), .B (n_13_58), .C1 (n_16_55), .C2 (n_22_52) );
AOI211_X1 g_7_62 (.ZN (n_7_62), .A (n_10_61), .B (n_12_60), .C1 (n_15_57), .C2 (n_20_53) );
AOI211_X1 g_9_61 (.ZN (n_9_61), .A (n_9_63), .B (n_10_59), .C1 (n_13_58), .C2 (n_18_54) );
AOI211_X1 g_11_62 (.ZN (n_11_62), .A (n_7_62), .B (n_8_60), .C1 (n_12_60), .C2 (n_16_55) );
AOI211_X1 g_13_61 (.ZN (n_13_61), .A (n_9_61), .B (n_10_61), .C1 (n_10_59), .C2 (n_15_57) );
AOI211_X1 g_14_59 (.ZN (n_14_59), .A (n_11_62), .B (n_9_63), .C1 (n_8_60), .C2 (n_13_58) );
AOI211_X1 g_12_58 (.ZN (n_12_58), .A (n_13_61), .B (n_7_62), .C1 (n_10_61), .C2 (n_12_60) );
AOI211_X1 g_11_60 (.ZN (n_11_60), .A (n_14_59), .B (n_9_61), .C1 (n_9_63), .C2 (n_10_59) );
AOI211_X1 g_13_59 (.ZN (n_13_59), .A (n_12_58), .B (n_11_62), .C1 (n_7_62), .C2 (n_8_60) );
AOI211_X1 g_14_57 (.ZN (n_14_57), .A (n_11_60), .B (n_13_61), .C1 (n_9_61), .C2 (n_10_61) );
AOI211_X1 g_16_56 (.ZN (n_16_56), .A (n_13_59), .B (n_14_59), .C1 (n_11_62), .C2 (n_9_63) );
AOI211_X1 g_18_55 (.ZN (n_18_55), .A (n_14_57), .B (n_12_58), .C1 (n_13_61), .C2 (n_7_62) );
AOI211_X1 g_20_54 (.ZN (n_20_54), .A (n_16_56), .B (n_11_60), .C1 (n_14_59), .C2 (n_9_61) );
AOI211_X1 g_22_53 (.ZN (n_22_53), .A (n_18_55), .B (n_13_59), .C1 (n_12_58), .C2 (n_11_62) );
AOI211_X1 g_24_52 (.ZN (n_24_52), .A (n_20_54), .B (n_14_57), .C1 (n_11_60), .C2 (n_13_61) );
AOI211_X1 g_26_51 (.ZN (n_26_51), .A (n_22_53), .B (n_16_56), .C1 (n_13_59), .C2 (n_14_59) );
AOI211_X1 g_28_50 (.ZN (n_28_50), .A (n_24_52), .B (n_18_55), .C1 (n_14_57), .C2 (n_12_58) );
AOI211_X1 g_30_49 (.ZN (n_30_49), .A (n_26_51), .B (n_20_54), .C1 (n_16_56), .C2 (n_11_60) );
AOI211_X1 g_29_51 (.ZN (n_29_51), .A (n_28_50), .B (n_22_53), .C1 (n_18_55), .C2 (n_13_59) );
AOI211_X1 g_31_50 (.ZN (n_31_50), .A (n_30_49), .B (n_24_52), .C1 (n_20_54), .C2 (n_14_57) );
AOI211_X1 g_33_49 (.ZN (n_33_49), .A (n_29_51), .B (n_26_51), .C1 (n_22_53), .C2 (n_16_56) );
AOI211_X1 g_32_51 (.ZN (n_32_51), .A (n_31_50), .B (n_28_50), .C1 (n_24_52), .C2 (n_18_55) );
AOI211_X1 g_31_49 (.ZN (n_31_49), .A (n_33_49), .B (n_30_49), .C1 (n_26_51), .C2 (n_20_54) );
AOI211_X1 g_33_48 (.ZN (n_33_48), .A (n_32_51), .B (n_29_51), .C1 (n_28_50), .C2 (n_22_53) );
AOI211_X1 g_35_47 (.ZN (n_35_47), .A (n_31_49), .B (n_31_50), .C1 (n_30_49), .C2 (n_24_52) );
AOI211_X1 g_37_46 (.ZN (n_37_46), .A (n_33_48), .B (n_33_49), .C1 (n_29_51), .C2 (n_26_51) );
AOI211_X1 g_36_48 (.ZN (n_36_48), .A (n_35_47), .B (n_32_51), .C1 (n_31_50), .C2 (n_28_50) );
AOI211_X1 g_38_47 (.ZN (n_38_47), .A (n_37_46), .B (n_31_49), .C1 (n_33_49), .C2 (n_30_49) );
AOI211_X1 g_40_46 (.ZN (n_40_46), .A (n_36_48), .B (n_33_48), .C1 (n_32_51), .C2 (n_29_51) );
AOI211_X1 g_42_45 (.ZN (n_42_45), .A (n_38_47), .B (n_35_47), .C1 (n_31_49), .C2 (n_31_50) );
AOI211_X1 g_44_44 (.ZN (n_44_44), .A (n_40_46), .B (n_37_46), .C1 (n_33_48), .C2 (n_33_49) );
AOI211_X1 g_46_43 (.ZN (n_46_43), .A (n_42_45), .B (n_36_48), .C1 (n_35_47), .C2 (n_32_51) );
AOI211_X1 g_48_42 (.ZN (n_48_42), .A (n_44_44), .B (n_38_47), .C1 (n_37_46), .C2 (n_31_49) );
AOI211_X1 g_50_41 (.ZN (n_50_41), .A (n_46_43), .B (n_40_46), .C1 (n_36_48), .C2 (n_33_48) );
AOI211_X1 g_52_40 (.ZN (n_52_40), .A (n_48_42), .B (n_42_45), .C1 (n_38_47), .C2 (n_35_47) );
AOI211_X1 g_54_39 (.ZN (n_54_39), .A (n_50_41), .B (n_44_44), .C1 (n_40_46), .C2 (n_37_46) );
AOI211_X1 g_56_38 (.ZN (n_56_38), .A (n_52_40), .B (n_46_43), .C1 (n_42_45), .C2 (n_36_48) );
AOI211_X1 g_58_37 (.ZN (n_58_37), .A (n_54_39), .B (n_48_42), .C1 (n_44_44), .C2 (n_38_47) );
AOI211_X1 g_60_36 (.ZN (n_60_36), .A (n_56_38), .B (n_50_41), .C1 (n_46_43), .C2 (n_40_46) );
AOI211_X1 g_62_35 (.ZN (n_62_35), .A (n_58_37), .B (n_52_40), .C1 (n_48_42), .C2 (n_42_45) );
AOI211_X1 g_61_37 (.ZN (n_61_37), .A (n_60_36), .B (n_54_39), .C1 (n_50_41), .C2 (n_44_44) );
AOI211_X1 g_63_36 (.ZN (n_63_36), .A (n_62_35), .B (n_56_38), .C1 (n_52_40), .C2 (n_46_43) );
AOI211_X1 g_65_35 (.ZN (n_65_35), .A (n_61_37), .B (n_58_37), .C1 (n_54_39), .C2 (n_48_42) );
AOI211_X1 g_67_34 (.ZN (n_67_34), .A (n_63_36), .B (n_60_36), .C1 (n_56_38), .C2 (n_50_41) );
AOI211_X1 g_69_33 (.ZN (n_69_33), .A (n_65_35), .B (n_62_35), .C1 (n_58_37), .C2 (n_52_40) );
AOI211_X1 g_71_32 (.ZN (n_71_32), .A (n_67_34), .B (n_61_37), .C1 (n_60_36), .C2 (n_54_39) );
AOI211_X1 g_73_31 (.ZN (n_73_31), .A (n_69_33), .B (n_63_36), .C1 (n_62_35), .C2 (n_56_38) );
AOI211_X1 g_75_30 (.ZN (n_75_30), .A (n_71_32), .B (n_65_35), .C1 (n_61_37), .C2 (n_58_37) );
AOI211_X1 g_77_29 (.ZN (n_77_29), .A (n_73_31), .B (n_67_34), .C1 (n_63_36), .C2 (n_60_36) );
AOI211_X1 g_79_28 (.ZN (n_79_28), .A (n_75_30), .B (n_69_33), .C1 (n_65_35), .C2 (n_62_35) );
AOI211_X1 g_81_27 (.ZN (n_81_27), .A (n_77_29), .B (n_71_32), .C1 (n_67_34), .C2 (n_61_37) );
AOI211_X1 g_83_26 (.ZN (n_83_26), .A (n_79_28), .B (n_73_31), .C1 (n_69_33), .C2 (n_63_36) );
AOI211_X1 g_85_25 (.ZN (n_85_25), .A (n_81_27), .B (n_75_30), .C1 (n_71_32), .C2 (n_65_35) );
AOI211_X1 g_87_24 (.ZN (n_87_24), .A (n_83_26), .B (n_77_29), .C1 (n_73_31), .C2 (n_67_34) );
AOI211_X1 g_89_23 (.ZN (n_89_23), .A (n_85_25), .B (n_79_28), .C1 (n_75_30), .C2 (n_69_33) );
AOI211_X1 g_91_22 (.ZN (n_91_22), .A (n_87_24), .B (n_81_27), .C1 (n_77_29), .C2 (n_71_32) );
AOI211_X1 g_93_21 (.ZN (n_93_21), .A (n_89_23), .B (n_83_26), .C1 (n_79_28), .C2 (n_73_31) );
AOI211_X1 g_92_23 (.ZN (n_92_23), .A (n_91_22), .B (n_85_25), .C1 (n_81_27), .C2 (n_75_30) );
AOI211_X1 g_94_22 (.ZN (n_94_22), .A (n_93_21), .B (n_87_24), .C1 (n_83_26), .C2 (n_77_29) );
AOI211_X1 g_96_21 (.ZN (n_96_21), .A (n_92_23), .B (n_89_23), .C1 (n_85_25), .C2 (n_79_28) );
AOI211_X1 g_98_20 (.ZN (n_98_20), .A (n_94_22), .B (n_91_22), .C1 (n_87_24), .C2 (n_81_27) );
AOI211_X1 g_100_19 (.ZN (n_100_19), .A (n_96_21), .B (n_93_21), .C1 (n_89_23), .C2 (n_83_26) );
AOI211_X1 g_99_21 (.ZN (n_99_21), .A (n_98_20), .B (n_92_23), .C1 (n_91_22), .C2 (n_85_25) );
AOI211_X1 g_101_20 (.ZN (n_101_20), .A (n_100_19), .B (n_94_22), .C1 (n_93_21), .C2 (n_87_24) );
AOI211_X1 g_100_22 (.ZN (n_100_22), .A (n_99_21), .B (n_96_21), .C1 (n_92_23), .C2 (n_89_23) );
AOI211_X1 g_99_20 (.ZN (n_99_20), .A (n_101_20), .B (n_98_20), .C1 (n_94_22), .C2 (n_91_22) );
AOI211_X1 g_101_19 (.ZN (n_101_19), .A (n_100_22), .B (n_100_19), .C1 (n_96_21), .C2 (n_93_21) );
AOI211_X1 g_103_18 (.ZN (n_103_18), .A (n_99_20), .B (n_99_21), .C1 (n_98_20), .C2 (n_92_23) );
AOI211_X1 g_105_17 (.ZN (n_105_17), .A (n_101_19), .B (n_101_20), .C1 (n_100_19), .C2 (n_94_22) );
AOI211_X1 g_107_16 (.ZN (n_107_16), .A (n_103_18), .B (n_100_22), .C1 (n_99_21), .C2 (n_96_21) );
AOI211_X1 g_106_18 (.ZN (n_106_18), .A (n_105_17), .B (n_99_20), .C1 (n_101_20), .C2 (n_98_20) );
AOI211_X1 g_104_19 (.ZN (n_104_19), .A (n_107_16), .B (n_101_19), .C1 (n_100_22), .C2 (n_100_19) );
AOI211_X1 g_102_20 (.ZN (n_102_20), .A (n_106_18), .B (n_103_18), .C1 (n_99_20), .C2 (n_99_21) );
AOI211_X1 g_100_21 (.ZN (n_100_21), .A (n_104_19), .B (n_105_17), .C1 (n_101_19), .C2 (n_101_20) );
AOI211_X1 g_98_22 (.ZN (n_98_22), .A (n_102_20), .B (n_107_16), .C1 (n_103_18), .C2 (n_100_22) );
AOI211_X1 g_96_23 (.ZN (n_96_23), .A (n_100_21), .B (n_106_18), .C1 (n_105_17), .C2 (n_99_20) );
AOI211_X1 g_97_21 (.ZN (n_97_21), .A (n_98_22), .B (n_104_19), .C1 (n_107_16), .C2 (n_101_19) );
AOI211_X1 g_95_22 (.ZN (n_95_22), .A (n_96_23), .B (n_102_20), .C1 (n_106_18), .C2 (n_103_18) );
AOI211_X1 g_93_23 (.ZN (n_93_23), .A (n_97_21), .B (n_100_21), .C1 (n_104_19), .C2 (n_105_17) );
AOI211_X1 g_91_24 (.ZN (n_91_24), .A (n_95_22), .B (n_98_22), .C1 (n_102_20), .C2 (n_107_16) );
AOI211_X1 g_89_25 (.ZN (n_89_25), .A (n_93_23), .B (n_96_23), .C1 (n_100_21), .C2 (n_106_18) );
AOI211_X1 g_88_27 (.ZN (n_88_27), .A (n_91_24), .B (n_97_21), .C1 (n_98_22), .C2 (n_104_19) );
AOI211_X1 g_86_26 (.ZN (n_86_26), .A (n_89_25), .B (n_95_22), .C1 (n_96_23), .C2 (n_102_20) );
AOI211_X1 g_88_25 (.ZN (n_88_25), .A (n_88_27), .B (n_93_23), .C1 (n_97_21), .C2 (n_100_21) );
AOI211_X1 g_90_24 (.ZN (n_90_24), .A (n_86_26), .B (n_91_24), .C1 (n_95_22), .C2 (n_98_22) );
AOI211_X1 g_89_26 (.ZN (n_89_26), .A (n_88_25), .B (n_89_25), .C1 (n_93_23), .C2 (n_96_23) );
AOI211_X1 g_91_25 (.ZN (n_91_25), .A (n_90_24), .B (n_88_27), .C1 (n_91_24), .C2 (n_97_21) );
AOI211_X1 g_93_24 (.ZN (n_93_24), .A (n_89_26), .B (n_86_26), .C1 (n_89_25), .C2 (n_95_22) );
AOI211_X1 g_95_23 (.ZN (n_95_23), .A (n_91_25), .B (n_88_25), .C1 (n_88_27), .C2 (n_93_23) );
AOI211_X1 g_97_22 (.ZN (n_97_22), .A (n_93_24), .B (n_90_24), .C1 (n_86_26), .C2 (n_91_24) );
AOI211_X1 g_96_24 (.ZN (n_96_24), .A (n_95_23), .B (n_89_26), .C1 (n_88_25), .C2 (n_89_25) );
AOI211_X1 g_98_23 (.ZN (n_98_23), .A (n_97_22), .B (n_91_25), .C1 (n_90_24), .C2 (n_88_27) );
AOI211_X1 g_96_22 (.ZN (n_96_22), .A (n_96_24), .B (n_93_24), .C1 (n_89_26), .C2 (n_86_26) );
AOI211_X1 g_98_21 (.ZN (n_98_21), .A (n_98_23), .B (n_95_23), .C1 (n_91_25), .C2 (n_88_25) );
AOI211_X1 g_100_20 (.ZN (n_100_20), .A (n_96_22), .B (n_97_22), .C1 (n_93_24), .C2 (n_90_24) );
AOI211_X1 g_102_19 (.ZN (n_102_19), .A (n_98_21), .B (n_96_24), .C1 (n_95_23), .C2 (n_89_26) );
AOI211_X1 g_104_18 (.ZN (n_104_18), .A (n_100_20), .B (n_98_23), .C1 (n_97_22), .C2 (n_91_25) );
AOI211_X1 g_105_20 (.ZN (n_105_20), .A (n_102_19), .B (n_96_22), .C1 (n_96_24), .C2 (n_93_24) );
AOI211_X1 g_103_21 (.ZN (n_103_21), .A (n_104_18), .B (n_98_21), .C1 (n_98_23), .C2 (n_95_23) );
AOI211_X1 g_101_22 (.ZN (n_101_22), .A (n_105_20), .B (n_100_20), .C1 (n_96_22), .C2 (n_97_22) );
AOI211_X1 g_99_23 (.ZN (n_99_23), .A (n_103_21), .B (n_102_19), .C1 (n_98_21), .C2 (n_96_24) );
AOI211_X1 g_97_24 (.ZN (n_97_24), .A (n_101_22), .B (n_104_18), .C1 (n_100_20), .C2 (n_98_23) );
AOI211_X1 g_95_25 (.ZN (n_95_25), .A (n_99_23), .B (n_105_20), .C1 (n_102_19), .C2 (n_96_22) );
AOI211_X1 g_94_23 (.ZN (n_94_23), .A (n_97_24), .B (n_103_21), .C1 (n_104_18), .C2 (n_98_21) );
AOI211_X1 g_92_24 (.ZN (n_92_24), .A (n_95_25), .B (n_101_22), .C1 (n_105_20), .C2 (n_100_20) );
AOI211_X1 g_90_25 (.ZN (n_90_25), .A (n_94_23), .B (n_99_23), .C1 (n_103_21), .C2 (n_102_19) );
AOI211_X1 g_88_26 (.ZN (n_88_26), .A (n_92_24), .B (n_97_24), .C1 (n_101_22), .C2 (n_104_18) );
AOI211_X1 g_86_27 (.ZN (n_86_27), .A (n_90_25), .B (n_95_25), .C1 (n_99_23), .C2 (n_105_20) );
AOI211_X1 g_84_28 (.ZN (n_84_28), .A (n_88_26), .B (n_94_23), .C1 (n_97_24), .C2 (n_103_21) );
AOI211_X1 g_82_29 (.ZN (n_82_29), .A (n_86_27), .B (n_92_24), .C1 (n_95_25), .C2 (n_101_22) );
AOI211_X1 g_80_28 (.ZN (n_80_28), .A (n_84_28), .B (n_90_25), .C1 (n_94_23), .C2 (n_99_23) );
AOI211_X1 g_78_29 (.ZN (n_78_29), .A (n_82_29), .B (n_88_26), .C1 (n_92_24), .C2 (n_97_24) );
AOI211_X1 g_76_30 (.ZN (n_76_30), .A (n_80_28), .B (n_86_27), .C1 (n_90_25), .C2 (n_95_25) );
AOI211_X1 g_74_31 (.ZN (n_74_31), .A (n_78_29), .B (n_84_28), .C1 (n_88_26), .C2 (n_94_23) );
AOI211_X1 g_72_32 (.ZN (n_72_32), .A (n_76_30), .B (n_82_29), .C1 (n_86_27), .C2 (n_92_24) );
AOI211_X1 g_73_30 (.ZN (n_73_30), .A (n_74_31), .B (n_80_28), .C1 (n_84_28), .C2 (n_90_25) );
AOI211_X1 g_71_31 (.ZN (n_71_31), .A (n_72_32), .B (n_78_29), .C1 (n_82_29), .C2 (n_88_26) );
AOI211_X1 g_69_32 (.ZN (n_69_32), .A (n_73_30), .B (n_76_30), .C1 (n_80_28), .C2 (n_86_27) );
AOI211_X1 g_67_33 (.ZN (n_67_33), .A (n_71_31), .B (n_74_31), .C1 (n_78_29), .C2 (n_84_28) );
AOI211_X1 g_65_34 (.ZN (n_65_34), .A (n_69_32), .B (n_72_32), .C1 (n_76_30), .C2 (n_82_29) );
AOI211_X1 g_63_35 (.ZN (n_63_35), .A (n_67_33), .B (n_73_30), .C1 (n_74_31), .C2 (n_80_28) );
AOI211_X1 g_61_36 (.ZN (n_61_36), .A (n_65_34), .B (n_71_31), .C1 (n_72_32), .C2 (n_78_29) );
AOI211_X1 g_59_37 (.ZN (n_59_37), .A (n_63_35), .B (n_69_32), .C1 (n_73_30), .C2 (n_76_30) );
AOI211_X1 g_57_38 (.ZN (n_57_38), .A (n_61_36), .B (n_67_33), .C1 (n_71_31), .C2 (n_74_31) );
AOI211_X1 g_55_39 (.ZN (n_55_39), .A (n_59_37), .B (n_65_34), .C1 (n_69_32), .C2 (n_72_32) );
AOI211_X1 g_53_40 (.ZN (n_53_40), .A (n_57_38), .B (n_63_35), .C1 (n_67_33), .C2 (n_73_30) );
AOI211_X1 g_51_41 (.ZN (n_51_41), .A (n_55_39), .B (n_61_36), .C1 (n_65_34), .C2 (n_71_31) );
AOI211_X1 g_49_42 (.ZN (n_49_42), .A (n_53_40), .B (n_59_37), .C1 (n_63_35), .C2 (n_69_32) );
AOI211_X1 g_47_43 (.ZN (n_47_43), .A (n_51_41), .B (n_57_38), .C1 (n_61_36), .C2 (n_67_33) );
AOI211_X1 g_45_44 (.ZN (n_45_44), .A (n_49_42), .B (n_55_39), .C1 (n_59_37), .C2 (n_65_34) );
AOI211_X1 g_43_45 (.ZN (n_43_45), .A (n_47_43), .B (n_53_40), .C1 (n_57_38), .C2 (n_63_35) );
AOI211_X1 g_41_46 (.ZN (n_41_46), .A (n_45_44), .B (n_51_41), .C1 (n_55_39), .C2 (n_61_36) );
AOI211_X1 g_42_44 (.ZN (n_42_44), .A (n_43_45), .B (n_49_42), .C1 (n_53_40), .C2 (n_59_37) );
AOI211_X1 g_40_45 (.ZN (n_40_45), .A (n_41_46), .B (n_47_43), .C1 (n_51_41), .C2 (n_57_38) );
AOI211_X1 g_39_47 (.ZN (n_39_47), .A (n_42_44), .B (n_45_44), .C1 (n_49_42), .C2 (n_55_39) );
AOI211_X1 g_37_48 (.ZN (n_37_48), .A (n_40_45), .B (n_43_45), .C1 (n_47_43), .C2 (n_53_40) );
AOI211_X1 g_35_49 (.ZN (n_35_49), .A (n_39_47), .B (n_41_46), .C1 (n_45_44), .C2 (n_51_41) );
AOI211_X1 g_33_50 (.ZN (n_33_50), .A (n_37_48), .B (n_42_44), .C1 (n_43_45), .C2 (n_49_42) );
AOI211_X1 g_31_51 (.ZN (n_31_51), .A (n_35_49), .B (n_40_45), .C1 (n_41_46), .C2 (n_47_43) );
AOI211_X1 g_29_52 (.ZN (n_29_52), .A (n_33_50), .B (n_39_47), .C1 (n_42_44), .C2 (n_45_44) );
AOI211_X1 g_27_53 (.ZN (n_27_53), .A (n_31_51), .B (n_37_48), .C1 (n_40_45), .C2 (n_43_45) );
AOI211_X1 g_28_51 (.ZN (n_28_51), .A (n_29_52), .B (n_35_49), .C1 (n_39_47), .C2 (n_41_46) );
AOI211_X1 g_26_52 (.ZN (n_26_52), .A (n_27_53), .B (n_33_50), .C1 (n_37_48), .C2 (n_42_44) );
AOI211_X1 g_24_53 (.ZN (n_24_53), .A (n_28_51), .B (n_31_51), .C1 (n_35_49), .C2 (n_40_45) );
AOI211_X1 g_22_54 (.ZN (n_22_54), .A (n_26_52), .B (n_29_52), .C1 (n_33_50), .C2 (n_39_47) );
AOI211_X1 g_20_55 (.ZN (n_20_55), .A (n_24_53), .B (n_27_53), .C1 (n_31_51), .C2 (n_37_48) );
AOI211_X1 g_18_56 (.ZN (n_18_56), .A (n_22_54), .B (n_28_51), .C1 (n_29_52), .C2 (n_35_49) );
AOI211_X1 g_16_57 (.ZN (n_16_57), .A (n_20_55), .B (n_26_52), .C1 (n_27_53), .C2 (n_33_50) );
AOI211_X1 g_14_58 (.ZN (n_14_58), .A (n_18_56), .B (n_24_53), .C1 (n_28_51), .C2 (n_31_51) );
AOI211_X1 g_13_60 (.ZN (n_13_60), .A (n_16_57), .B (n_22_54), .C1 (n_26_52), .C2 (n_29_52) );
AOI211_X1 g_15_59 (.ZN (n_15_59), .A (n_14_58), .B (n_20_55), .C1 (n_24_53), .C2 (n_27_53) );
AOI211_X1 g_17_58 (.ZN (n_17_58), .A (n_13_60), .B (n_18_56), .C1 (n_22_54), .C2 (n_28_51) );
AOI211_X1 g_19_57 (.ZN (n_19_57), .A (n_15_59), .B (n_16_57), .C1 (n_20_55), .C2 (n_26_52) );
AOI211_X1 g_17_56 (.ZN (n_17_56), .A (n_17_58), .B (n_14_58), .C1 (n_18_56), .C2 (n_24_53) );
AOI211_X1 g_19_55 (.ZN (n_19_55), .A (n_19_57), .B (n_13_60), .C1 (n_16_57), .C2 (n_22_54) );
AOI211_X1 g_21_54 (.ZN (n_21_54), .A (n_17_56), .B (n_15_59), .C1 (n_14_58), .C2 (n_20_55) );
AOI211_X1 g_23_53 (.ZN (n_23_53), .A (n_19_55), .B (n_17_58), .C1 (n_13_60), .C2 (n_18_56) );
AOI211_X1 g_25_54 (.ZN (n_25_54), .A (n_21_54), .B (n_19_57), .C1 (n_15_59), .C2 (n_16_57) );
AOI211_X1 g_23_55 (.ZN (n_23_55), .A (n_23_53), .B (n_17_56), .C1 (n_17_58), .C2 (n_14_58) );
AOI211_X1 g_21_56 (.ZN (n_21_56), .A (n_25_54), .B (n_19_55), .C1 (n_19_57), .C2 (n_13_60) );
AOI211_X1 g_20_58 (.ZN (n_20_58), .A (n_23_55), .B (n_21_54), .C1 (n_17_56), .C2 (n_15_59) );
AOI211_X1 g_19_56 (.ZN (n_19_56), .A (n_21_56), .B (n_23_53), .C1 (n_19_55), .C2 (n_17_58) );
AOI211_X1 g_21_55 (.ZN (n_21_55), .A (n_20_58), .B (n_25_54), .C1 (n_21_54), .C2 (n_19_57) );
AOI211_X1 g_23_54 (.ZN (n_23_54), .A (n_19_56), .B (n_23_55), .C1 (n_23_53), .C2 (n_17_56) );
AOI211_X1 g_25_53 (.ZN (n_25_53), .A (n_21_55), .B (n_21_56), .C1 (n_25_54), .C2 (n_19_55) );
AOI211_X1 g_27_52 (.ZN (n_27_52), .A (n_23_54), .B (n_20_58), .C1 (n_23_55), .C2 (n_21_54) );
AOI211_X1 g_26_54 (.ZN (n_26_54), .A (n_25_53), .B (n_19_56), .C1 (n_21_56), .C2 (n_23_53) );
AOI211_X1 g_28_53 (.ZN (n_28_53), .A (n_27_52), .B (n_21_55), .C1 (n_20_58), .C2 (n_25_54) );
AOI211_X1 g_30_52 (.ZN (n_30_52), .A (n_26_54), .B (n_23_54), .C1 (n_19_56), .C2 (n_23_55) );
AOI211_X1 g_29_54 (.ZN (n_29_54), .A (n_28_53), .B (n_25_53), .C1 (n_21_55), .C2 (n_21_56) );
AOI211_X1 g_28_52 (.ZN (n_28_52), .A (n_30_52), .B (n_27_52), .C1 (n_23_54), .C2 (n_20_58) );
AOI211_X1 g_30_51 (.ZN (n_30_51), .A (n_29_54), .B (n_26_54), .C1 (n_25_53), .C2 (n_19_56) );
AOI211_X1 g_32_50 (.ZN (n_32_50), .A (n_28_52), .B (n_28_53), .C1 (n_27_52), .C2 (n_21_55) );
AOI211_X1 g_34_49 (.ZN (n_34_49), .A (n_30_51), .B (n_30_52), .C1 (n_26_54), .C2 (n_23_54) );
AOI211_X1 g_33_51 (.ZN (n_33_51), .A (n_32_50), .B (n_29_54), .C1 (n_28_53), .C2 (n_25_53) );
AOI211_X1 g_35_50 (.ZN (n_35_50), .A (n_34_49), .B (n_28_52), .C1 (n_30_52), .C2 (n_27_52) );
AOI211_X1 g_37_49 (.ZN (n_37_49), .A (n_33_51), .B (n_30_51), .C1 (n_29_54), .C2 (n_26_54) );
AOI211_X1 g_39_48 (.ZN (n_39_48), .A (n_35_50), .B (n_32_50), .C1 (n_28_52), .C2 (n_28_53) );
AOI211_X1 g_37_47 (.ZN (n_37_47), .A (n_37_49), .B (n_34_49), .C1 (n_30_51), .C2 (n_30_52) );
AOI211_X1 g_39_46 (.ZN (n_39_46), .A (n_39_48), .B (n_33_51), .C1 (n_32_50), .C2 (n_29_54) );
AOI211_X1 g_41_45 (.ZN (n_41_45), .A (n_37_47), .B (n_35_50), .C1 (n_34_49), .C2 (n_28_52) );
AOI211_X1 g_43_44 (.ZN (n_43_44), .A (n_39_46), .B (n_37_49), .C1 (n_33_51), .C2 (n_30_51) );
AOI211_X1 g_45_43 (.ZN (n_45_43), .A (n_41_45), .B (n_39_48), .C1 (n_35_50), .C2 (n_32_50) );
AOI211_X1 g_47_42 (.ZN (n_47_42), .A (n_43_44), .B (n_37_47), .C1 (n_37_49), .C2 (n_34_49) );
AOI211_X1 g_46_44 (.ZN (n_46_44), .A (n_45_43), .B (n_39_46), .C1 (n_39_48), .C2 (n_33_51) );
AOI211_X1 g_48_43 (.ZN (n_48_43), .A (n_47_42), .B (n_41_45), .C1 (n_37_47), .C2 (n_35_50) );
AOI211_X1 g_50_42 (.ZN (n_50_42), .A (n_46_44), .B (n_43_44), .C1 (n_39_46), .C2 (n_37_49) );
AOI211_X1 g_52_41 (.ZN (n_52_41), .A (n_48_43), .B (n_45_43), .C1 (n_41_45), .C2 (n_39_48) );
AOI211_X1 g_54_40 (.ZN (n_54_40), .A (n_50_42), .B (n_47_42), .C1 (n_43_44), .C2 (n_37_47) );
AOI211_X1 g_56_39 (.ZN (n_56_39), .A (n_52_41), .B (n_46_44), .C1 (n_45_43), .C2 (n_39_46) );
AOI211_X1 g_58_38 (.ZN (n_58_38), .A (n_54_40), .B (n_48_43), .C1 (n_47_42), .C2 (n_41_45) );
AOI211_X1 g_60_37 (.ZN (n_60_37), .A (n_56_39), .B (n_50_42), .C1 (n_46_44), .C2 (n_43_44) );
AOI211_X1 g_62_36 (.ZN (n_62_36), .A (n_58_38), .B (n_52_41), .C1 (n_48_43), .C2 (n_45_43) );
AOI211_X1 g_61_38 (.ZN (n_61_38), .A (n_60_37), .B (n_54_40), .C1 (n_50_42), .C2 (n_47_42) );
AOI211_X1 g_63_37 (.ZN (n_63_37), .A (n_62_36), .B (n_56_39), .C1 (n_52_41), .C2 (n_46_44) );
AOI211_X1 g_65_36 (.ZN (n_65_36), .A (n_61_38), .B (n_58_38), .C1 (n_54_40), .C2 (n_48_43) );
AOI211_X1 g_67_35 (.ZN (n_67_35), .A (n_63_37), .B (n_60_37), .C1 (n_56_39), .C2 (n_50_42) );
AOI211_X1 g_69_34 (.ZN (n_69_34), .A (n_65_36), .B (n_62_36), .C1 (n_58_38), .C2 (n_52_41) );
AOI211_X1 g_70_32 (.ZN (n_70_32), .A (n_67_35), .B (n_61_38), .C1 (n_60_37), .C2 (n_54_40) );
AOI211_X1 g_72_31 (.ZN (n_72_31), .A (n_69_34), .B (n_63_37), .C1 (n_62_36), .C2 (n_56_39) );
AOI211_X1 g_74_30 (.ZN (n_74_30), .A (n_70_32), .B (n_65_36), .C1 (n_61_38), .C2 (n_58_38) );
AOI211_X1 g_76_29 (.ZN (n_76_29), .A (n_72_31), .B (n_67_35), .C1 (n_63_37), .C2 (n_60_37) );
AOI211_X1 g_75_31 (.ZN (n_75_31), .A (n_74_30), .B (n_69_34), .C1 (n_65_36), .C2 (n_62_36) );
AOI211_X1 g_77_30 (.ZN (n_77_30), .A (n_76_29), .B (n_70_32), .C1 (n_67_35), .C2 (n_61_38) );
AOI211_X1 g_76_32 (.ZN (n_76_32), .A (n_75_31), .B (n_72_31), .C1 (n_69_34), .C2 (n_63_37) );
AOI211_X1 g_78_31 (.ZN (n_78_31), .A (n_77_30), .B (n_74_30), .C1 (n_70_32), .C2 (n_65_36) );
AOI211_X1 g_80_30 (.ZN (n_80_30), .A (n_76_32), .B (n_76_29), .C1 (n_72_31), .C2 (n_67_35) );
AOI211_X1 g_79_32 (.ZN (n_79_32), .A (n_78_31), .B (n_75_31), .C1 (n_74_30), .C2 (n_69_34) );
AOI211_X1 g_78_30 (.ZN (n_78_30), .A (n_80_30), .B (n_77_30), .C1 (n_76_29), .C2 (n_70_32) );
AOI211_X1 g_80_29 (.ZN (n_80_29), .A (n_79_32), .B (n_76_32), .C1 (n_75_31), .C2 (n_72_31) );
AOI211_X1 g_82_28 (.ZN (n_82_28), .A (n_78_30), .B (n_78_31), .C1 (n_77_30), .C2 (n_74_30) );
AOI211_X1 g_84_27 (.ZN (n_84_27), .A (n_80_29), .B (n_80_30), .C1 (n_76_32), .C2 (n_76_29) );
AOI211_X1 g_86_28 (.ZN (n_86_28), .A (n_82_28), .B (n_79_32), .C1 (n_78_31), .C2 (n_75_31) );
AOI211_X1 g_84_29 (.ZN (n_84_29), .A (n_84_27), .B (n_78_30), .C1 (n_80_30), .C2 (n_77_30) );
AOI211_X1 g_85_27 (.ZN (n_85_27), .A (n_86_28), .B (n_80_29), .C1 (n_79_32), .C2 (n_76_32) );
AOI211_X1 g_83_28 (.ZN (n_83_28), .A (n_84_29), .B (n_82_28), .C1 (n_78_30), .C2 (n_78_31) );
AOI211_X1 g_81_29 (.ZN (n_81_29), .A (n_85_27), .B (n_84_27), .C1 (n_80_29), .C2 (n_80_30) );
AOI211_X1 g_79_30 (.ZN (n_79_30), .A (n_83_28), .B (n_86_28), .C1 (n_82_28), .C2 (n_79_32) );
AOI211_X1 g_77_31 (.ZN (n_77_31), .A (n_81_29), .B (n_84_29), .C1 (n_84_27), .C2 (n_78_30) );
AOI211_X1 g_75_32 (.ZN (n_75_32), .A (n_79_30), .B (n_85_27), .C1 (n_86_28), .C2 (n_80_29) );
AOI211_X1 g_73_33 (.ZN (n_73_33), .A (n_77_31), .B (n_83_28), .C1 (n_84_29), .C2 (n_82_28) );
AOI211_X1 g_71_34 (.ZN (n_71_34), .A (n_75_32), .B (n_81_29), .C1 (n_85_27), .C2 (n_84_27) );
AOI211_X1 g_69_35 (.ZN (n_69_35), .A (n_73_33), .B (n_79_30), .C1 (n_83_28), .C2 (n_86_28) );
AOI211_X1 g_70_33 (.ZN (n_70_33), .A (n_71_34), .B (n_77_31), .C1 (n_81_29), .C2 (n_84_29) );
AOI211_X1 g_68_34 (.ZN (n_68_34), .A (n_69_35), .B (n_75_32), .C1 (n_79_30), .C2 (n_85_27) );
AOI211_X1 g_66_35 (.ZN (n_66_35), .A (n_70_33), .B (n_73_33), .C1 (n_77_31), .C2 (n_83_28) );
AOI211_X1 g_64_36 (.ZN (n_64_36), .A (n_68_34), .B (n_71_34), .C1 (n_75_32), .C2 (n_81_29) );
AOI211_X1 g_62_37 (.ZN (n_62_37), .A (n_66_35), .B (n_69_35), .C1 (n_73_33), .C2 (n_79_30) );
AOI211_X1 g_60_38 (.ZN (n_60_38), .A (n_64_36), .B (n_70_33), .C1 (n_71_34), .C2 (n_77_31) );
AOI211_X1 g_58_39 (.ZN (n_58_39), .A (n_62_37), .B (n_68_34), .C1 (n_69_35), .C2 (n_75_32) );
AOI211_X1 g_56_40 (.ZN (n_56_40), .A (n_60_38), .B (n_66_35), .C1 (n_70_33), .C2 (n_73_33) );
AOI211_X1 g_54_41 (.ZN (n_54_41), .A (n_58_39), .B (n_64_36), .C1 (n_68_34), .C2 (n_71_34) );
AOI211_X1 g_52_42 (.ZN (n_52_42), .A (n_56_40), .B (n_62_37), .C1 (n_66_35), .C2 (n_69_35) );
AOI211_X1 g_50_43 (.ZN (n_50_43), .A (n_54_41), .B (n_60_38), .C1 (n_64_36), .C2 (n_70_33) );
AOI211_X1 g_48_44 (.ZN (n_48_44), .A (n_52_42), .B (n_58_39), .C1 (n_62_37), .C2 (n_68_34) );
AOI211_X1 g_46_45 (.ZN (n_46_45), .A (n_50_43), .B (n_56_40), .C1 (n_60_38), .C2 (n_66_35) );
AOI211_X1 g_44_46 (.ZN (n_44_46), .A (n_48_44), .B (n_54_41), .C1 (n_58_39), .C2 (n_64_36) );
AOI211_X1 g_42_47 (.ZN (n_42_47), .A (n_46_45), .B (n_52_42), .C1 (n_56_40), .C2 (n_62_37) );
AOI211_X1 g_40_48 (.ZN (n_40_48), .A (n_44_46), .B (n_50_43), .C1 (n_54_41), .C2 (n_60_38) );
AOI211_X1 g_38_49 (.ZN (n_38_49), .A (n_42_47), .B (n_48_44), .C1 (n_52_42), .C2 (n_58_39) );
AOI211_X1 g_36_50 (.ZN (n_36_50), .A (n_40_48), .B (n_46_45), .C1 (n_50_43), .C2 (n_56_40) );
AOI211_X1 g_34_51 (.ZN (n_34_51), .A (n_38_49), .B (n_44_46), .C1 (n_48_44), .C2 (n_54_41) );
AOI211_X1 g_32_52 (.ZN (n_32_52), .A (n_36_50), .B (n_42_47), .C1 (n_46_45), .C2 (n_52_42) );
AOI211_X1 g_30_53 (.ZN (n_30_53), .A (n_34_51), .B (n_40_48), .C1 (n_44_46), .C2 (n_50_43) );
AOI211_X1 g_28_54 (.ZN (n_28_54), .A (n_32_52), .B (n_38_49), .C1 (n_42_47), .C2 (n_48_44) );
AOI211_X1 g_26_53 (.ZN (n_26_53), .A (n_30_53), .B (n_36_50), .C1 (n_40_48), .C2 (n_46_45) );
AOI211_X1 g_24_54 (.ZN (n_24_54), .A (n_28_54), .B (n_34_51), .C1 (n_38_49), .C2 (n_44_46) );
AOI211_X1 g_22_55 (.ZN (n_22_55), .A (n_26_53), .B (n_32_52), .C1 (n_36_50), .C2 (n_42_47) );
AOI211_X1 g_20_56 (.ZN (n_20_56), .A (n_24_54), .B (n_30_53), .C1 (n_34_51), .C2 (n_40_48) );
AOI211_X1 g_18_57 (.ZN (n_18_57), .A (n_22_55), .B (n_28_54), .C1 (n_32_52), .C2 (n_38_49) );
AOI211_X1 g_16_58 (.ZN (n_16_58), .A (n_20_56), .B (n_26_53), .C1 (n_30_53), .C2 (n_36_50) );
AOI211_X1 g_15_60 (.ZN (n_15_60), .A (n_18_57), .B (n_24_54), .C1 (n_28_54), .C2 (n_34_51) );
AOI211_X1 g_17_59 (.ZN (n_17_59), .A (n_16_58), .B (n_22_55), .C1 (n_26_53), .C2 (n_32_52) );
AOI211_X1 g_15_58 (.ZN (n_15_58), .A (n_15_60), .B (n_20_56), .C1 (n_24_54), .C2 (n_30_53) );
AOI211_X1 g_17_57 (.ZN (n_17_57), .A (n_17_59), .B (n_18_57), .C1 (n_22_55), .C2 (n_28_54) );
AOI211_X1 g_18_59 (.ZN (n_18_59), .A (n_15_58), .B (n_16_58), .C1 (n_20_56), .C2 (n_26_53) );
AOI211_X1 g_16_60 (.ZN (n_16_60), .A (n_17_57), .B (n_15_60), .C1 (n_18_57), .C2 (n_24_54) );
AOI211_X1 g_14_61 (.ZN (n_14_61), .A (n_18_59), .B (n_17_59), .C1 (n_16_58), .C2 (n_22_55) );
AOI211_X1 g_12_62 (.ZN (n_12_62), .A (n_16_60), .B (n_15_58), .C1 (n_15_60), .C2 (n_20_56) );
AOI211_X1 g_10_63 (.ZN (n_10_63), .A (n_14_61), .B (n_17_57), .C1 (n_17_59), .C2 (n_18_57) );
AOI211_X1 g_11_61 (.ZN (n_11_61), .A (n_12_62), .B (n_18_59), .C1 (n_15_58), .C2 (n_16_58) );
AOI211_X1 g_9_62 (.ZN (n_9_62), .A (n_10_63), .B (n_16_60), .C1 (n_17_57), .C2 (n_15_60) );
AOI211_X1 g_7_63 (.ZN (n_7_63), .A (n_11_61), .B (n_14_61), .C1 (n_18_59), .C2 (n_17_59) );
AOI211_X1 g_6_65 (.ZN (n_6_65), .A (n_9_62), .B (n_12_62), .C1 (n_16_60), .C2 (n_15_58) );
AOI211_X1 g_8_64 (.ZN (n_8_64), .A (n_7_63), .B (n_10_63), .C1 (n_14_61), .C2 (n_17_57) );
AOI211_X1 g_7_66 (.ZN (n_7_66), .A (n_6_65), .B (n_11_61), .C1 (n_12_62), .C2 (n_18_59) );
AOI211_X1 g_6_64 (.ZN (n_6_64), .A (n_8_64), .B (n_9_62), .C1 (n_10_63), .C2 (n_16_60) );
AOI211_X1 g_8_63 (.ZN (n_8_63), .A (n_7_66), .B (n_7_63), .C1 (n_11_61), .C2 (n_14_61) );
AOI211_X1 g_10_62 (.ZN (n_10_62), .A (n_6_64), .B (n_6_65), .C1 (n_9_62), .C2 (n_12_62) );
AOI211_X1 g_12_61 (.ZN (n_12_61), .A (n_8_63), .B (n_8_64), .C1 (n_7_63), .C2 (n_10_63) );
AOI211_X1 g_14_60 (.ZN (n_14_60), .A (n_10_62), .B (n_7_66), .C1 (n_6_65), .C2 (n_11_61) );
AOI211_X1 g_16_59 (.ZN (n_16_59), .A (n_12_61), .B (n_6_64), .C1 (n_8_64), .C2 (n_9_62) );
AOI211_X1 g_18_58 (.ZN (n_18_58), .A (n_14_60), .B (n_8_63), .C1 (n_7_66), .C2 (n_7_63) );
AOI211_X1 g_20_57 (.ZN (n_20_57), .A (n_16_59), .B (n_10_62), .C1 (n_6_64), .C2 (n_6_65) );
AOI211_X1 g_22_56 (.ZN (n_22_56), .A (n_18_58), .B (n_12_61), .C1 (n_8_63), .C2 (n_8_64) );
AOI211_X1 g_24_55 (.ZN (n_24_55), .A (n_20_57), .B (n_14_60), .C1 (n_10_62), .C2 (n_7_66) );
AOI211_X1 g_23_57 (.ZN (n_23_57), .A (n_22_56), .B (n_16_59), .C1 (n_12_61), .C2 (n_6_64) );
AOI211_X1 g_25_56 (.ZN (n_25_56), .A (n_24_55), .B (n_18_58), .C1 (n_14_60), .C2 (n_8_63) );
AOI211_X1 g_27_55 (.ZN (n_27_55), .A (n_23_57), .B (n_20_57), .C1 (n_16_59), .C2 (n_10_62) );
AOI211_X1 g_29_56 (.ZN (n_29_56), .A (n_25_56), .B (n_22_56), .C1 (n_18_58), .C2 (n_12_61) );
AOI211_X1 g_31_55 (.ZN (n_31_55), .A (n_27_55), .B (n_24_55), .C1 (n_20_57), .C2 (n_14_60) );
AOI211_X1 g_32_53 (.ZN (n_32_53), .A (n_29_56), .B (n_23_57), .C1 (n_22_56), .C2 (n_16_59) );
AOI211_X1 g_34_52 (.ZN (n_34_52), .A (n_31_55), .B (n_25_56), .C1 (n_24_55), .C2 (n_18_58) );
AOI211_X1 g_36_51 (.ZN (n_36_51), .A (n_32_53), .B (n_27_55), .C1 (n_23_57), .C2 (n_20_57) );
AOI211_X1 g_34_50 (.ZN (n_34_50), .A (n_34_52), .B (n_29_56), .C1 (n_25_56), .C2 (n_22_56) );
AOI211_X1 g_36_49 (.ZN (n_36_49), .A (n_36_51), .B (n_31_55), .C1 (n_27_55), .C2 (n_24_55) );
AOI211_X1 g_38_48 (.ZN (n_38_48), .A (n_34_50), .B (n_32_53), .C1 (n_29_56), .C2 (n_23_57) );
AOI211_X1 g_40_47 (.ZN (n_40_47), .A (n_36_49), .B (n_34_52), .C1 (n_31_55), .C2 (n_25_56) );
AOI211_X1 g_42_46 (.ZN (n_42_46), .A (n_38_48), .B (n_36_51), .C1 (n_32_53), .C2 (n_27_55) );
AOI211_X1 g_44_45 (.ZN (n_44_45), .A (n_40_47), .B (n_34_50), .C1 (n_34_52), .C2 (n_29_56) );
AOI211_X1 g_43_47 (.ZN (n_43_47), .A (n_42_46), .B (n_36_49), .C1 (n_36_51), .C2 (n_31_55) );
AOI211_X1 g_45_46 (.ZN (n_45_46), .A (n_44_45), .B (n_38_48), .C1 (n_34_50), .C2 (n_32_53) );
AOI211_X1 g_47_45 (.ZN (n_47_45), .A (n_43_47), .B (n_40_47), .C1 (n_36_49), .C2 (n_34_52) );
AOI211_X1 g_49_44 (.ZN (n_49_44), .A (n_45_46), .B (n_42_46), .C1 (n_38_48), .C2 (n_36_51) );
AOI211_X1 g_51_43 (.ZN (n_51_43), .A (n_47_45), .B (n_44_45), .C1 (n_40_47), .C2 (n_34_50) );
AOI211_X1 g_53_42 (.ZN (n_53_42), .A (n_49_44), .B (n_43_47), .C1 (n_42_46), .C2 (n_36_49) );
AOI211_X1 g_55_41 (.ZN (n_55_41), .A (n_51_43), .B (n_45_46), .C1 (n_44_45), .C2 (n_38_48) );
AOI211_X1 g_57_40 (.ZN (n_57_40), .A (n_53_42), .B (n_47_45), .C1 (n_43_47), .C2 (n_40_47) );
AOI211_X1 g_59_39 (.ZN (n_59_39), .A (n_55_41), .B (n_49_44), .C1 (n_45_46), .C2 (n_42_46) );
AOI211_X1 g_58_41 (.ZN (n_58_41), .A (n_57_40), .B (n_51_43), .C1 (n_47_45), .C2 (n_44_45) );
AOI211_X1 g_57_39 (.ZN (n_57_39), .A (n_59_39), .B (n_53_42), .C1 (n_49_44), .C2 (n_43_47) );
AOI211_X1 g_59_38 (.ZN (n_59_38), .A (n_58_41), .B (n_55_41), .C1 (n_51_43), .C2 (n_45_46) );
AOI211_X1 g_60_40 (.ZN (n_60_40), .A (n_57_39), .B (n_57_40), .C1 (n_53_42), .C2 (n_47_45) );
AOI211_X1 g_62_39 (.ZN (n_62_39), .A (n_59_38), .B (n_59_39), .C1 (n_55_41), .C2 (n_49_44) );
AOI211_X1 g_64_38 (.ZN (n_64_38), .A (n_60_40), .B (n_58_41), .C1 (n_57_40), .C2 (n_51_43) );
AOI211_X1 g_66_37 (.ZN (n_66_37), .A (n_62_39), .B (n_57_39), .C1 (n_59_39), .C2 (n_53_42) );
AOI211_X1 g_68_36 (.ZN (n_68_36), .A (n_64_38), .B (n_59_38), .C1 (n_58_41), .C2 (n_55_41) );
AOI211_X1 g_70_35 (.ZN (n_70_35), .A (n_66_37), .B (n_60_40), .C1 (n_57_39), .C2 (n_57_40) );
AOI211_X1 g_71_33 (.ZN (n_71_33), .A (n_68_36), .B (n_62_39), .C1 (n_59_38), .C2 (n_59_39) );
AOI211_X1 g_73_32 (.ZN (n_73_32), .A (n_70_35), .B (n_64_38), .C1 (n_60_40), .C2 (n_58_41) );
AOI211_X1 g_72_34 (.ZN (n_72_34), .A (n_71_33), .B (n_66_37), .C1 (n_62_39), .C2 (n_57_39) );
AOI211_X1 g_74_33 (.ZN (n_74_33), .A (n_73_32), .B (n_68_36), .C1 (n_64_38), .C2 (n_59_38) );
AOI211_X1 g_73_35 (.ZN (n_73_35), .A (n_72_34), .B (n_70_35), .C1 (n_66_37), .C2 (n_60_40) );
AOI211_X1 g_72_33 (.ZN (n_72_33), .A (n_74_33), .B (n_71_33), .C1 (n_68_36), .C2 (n_62_39) );
AOI211_X1 g_74_32 (.ZN (n_74_32), .A (n_73_35), .B (n_73_32), .C1 (n_70_35), .C2 (n_64_38) );
AOI211_X1 g_76_31 (.ZN (n_76_31), .A (n_72_33), .B (n_72_34), .C1 (n_71_33), .C2 (n_66_37) );
AOI211_X1 g_77_33 (.ZN (n_77_33), .A (n_74_32), .B (n_74_33), .C1 (n_73_32), .C2 (n_68_36) );
AOI211_X1 g_75_34 (.ZN (n_75_34), .A (n_76_31), .B (n_73_35), .C1 (n_72_34), .C2 (n_70_35) );
AOI211_X1 g_74_36 (.ZN (n_74_36), .A (n_77_33), .B (n_72_33), .C1 (n_74_33), .C2 (n_71_33) );
AOI211_X1 g_73_34 (.ZN (n_73_34), .A (n_75_34), .B (n_74_32), .C1 (n_73_35), .C2 (n_73_32) );
AOI211_X1 g_75_33 (.ZN (n_75_33), .A (n_74_36), .B (n_76_31), .C1 (n_72_33), .C2 (n_72_34) );
AOI211_X1 g_77_32 (.ZN (n_77_32), .A (n_73_34), .B (n_77_33), .C1 (n_74_32), .C2 (n_74_33) );
AOI211_X1 g_79_31 (.ZN (n_79_31), .A (n_75_33), .B (n_75_34), .C1 (n_76_31), .C2 (n_73_35) );
AOI211_X1 g_81_30 (.ZN (n_81_30), .A (n_77_32), .B (n_74_36), .C1 (n_77_33), .C2 (n_72_33) );
AOI211_X1 g_83_29 (.ZN (n_83_29), .A (n_79_31), .B (n_73_34), .C1 (n_75_34), .C2 (n_74_32) );
AOI211_X1 g_85_28 (.ZN (n_85_28), .A (n_81_30), .B (n_75_33), .C1 (n_74_36), .C2 (n_76_31) );
AOI211_X1 g_87_27 (.ZN (n_87_27), .A (n_83_29), .B (n_77_32), .C1 (n_73_34), .C2 (n_77_33) );
AOI211_X1 g_86_29 (.ZN (n_86_29), .A (n_85_28), .B (n_79_31), .C1 (n_75_33), .C2 (n_75_34) );
AOI211_X1 g_88_28 (.ZN (n_88_28), .A (n_87_27), .B (n_81_30), .C1 (n_77_32), .C2 (n_74_36) );
AOI211_X1 g_90_27 (.ZN (n_90_27), .A (n_86_29), .B (n_83_29), .C1 (n_79_31), .C2 (n_73_34) );
AOI211_X1 g_92_26 (.ZN (n_92_26), .A (n_88_28), .B (n_85_28), .C1 (n_81_30), .C2 (n_75_33) );
AOI211_X1 g_94_25 (.ZN (n_94_25), .A (n_90_27), .B (n_87_27), .C1 (n_83_29), .C2 (n_77_32) );
AOI211_X1 g_96_26 (.ZN (n_96_26), .A (n_92_26), .B (n_86_29), .C1 (n_85_28), .C2 (n_79_31) );
AOI211_X1 g_95_24 (.ZN (n_95_24), .A (n_94_25), .B (n_88_28), .C1 (n_87_27), .C2 (n_81_30) );
AOI211_X1 g_97_23 (.ZN (n_97_23), .A (n_96_26), .B (n_90_27), .C1 (n_86_29), .C2 (n_83_29) );
AOI211_X1 g_99_22 (.ZN (n_99_22), .A (n_95_24), .B (n_92_26), .C1 (n_88_28), .C2 (n_85_28) );
AOI211_X1 g_101_21 (.ZN (n_101_21), .A (n_97_23), .B (n_94_25), .C1 (n_90_27), .C2 (n_87_27) );
AOI211_X1 g_103_20 (.ZN (n_103_20), .A (n_99_22), .B (n_96_26), .C1 (n_92_26), .C2 (n_86_29) );
AOI211_X1 g_105_19 (.ZN (n_105_19), .A (n_101_21), .B (n_95_24), .C1 (n_94_25), .C2 (n_88_28) );
AOI211_X1 g_107_18 (.ZN (n_107_18), .A (n_103_20), .B (n_97_23), .C1 (n_96_26), .C2 (n_90_27) );
AOI211_X1 g_109_17 (.ZN (n_109_17), .A (n_105_19), .B (n_99_22), .C1 (n_95_24), .C2 (n_92_26) );
AOI211_X1 g_111_16 (.ZN (n_111_16), .A (n_107_18), .B (n_101_21), .C1 (n_97_23), .C2 (n_94_25) );
AOI211_X1 g_113_17 (.ZN (n_113_17), .A (n_109_17), .B (n_103_20), .C1 (n_99_22), .C2 (n_96_26) );
AOI211_X1 g_111_18 (.ZN (n_111_18), .A (n_111_16), .B (n_105_19), .C1 (n_101_21), .C2 (n_95_24) );
AOI211_X1 g_109_19 (.ZN (n_109_19), .A (n_113_17), .B (n_107_18), .C1 (n_103_20), .C2 (n_97_23) );
AOI211_X1 g_107_20 (.ZN (n_107_20), .A (n_111_18), .B (n_109_17), .C1 (n_105_19), .C2 (n_99_22) );
AOI211_X1 g_108_18 (.ZN (n_108_18), .A (n_109_19), .B (n_111_16), .C1 (n_107_18), .C2 (n_101_21) );
AOI211_X1 g_106_19 (.ZN (n_106_19), .A (n_107_20), .B (n_113_17), .C1 (n_109_17), .C2 (n_103_20) );
AOI211_X1 g_104_20 (.ZN (n_104_20), .A (n_108_18), .B (n_111_18), .C1 (n_111_16), .C2 (n_105_19) );
AOI211_X1 g_102_21 (.ZN (n_102_21), .A (n_106_19), .B (n_109_19), .C1 (n_113_17), .C2 (n_107_18) );
AOI211_X1 g_101_23 (.ZN (n_101_23), .A (n_104_20), .B (n_107_20), .C1 (n_111_18), .C2 (n_109_17) );
AOI211_X1 g_103_22 (.ZN (n_103_22), .A (n_102_21), .B (n_108_18), .C1 (n_109_19), .C2 (n_111_16) );
AOI211_X1 g_105_21 (.ZN (n_105_21), .A (n_101_23), .B (n_106_19), .C1 (n_107_20), .C2 (n_113_17) );
AOI211_X1 g_104_23 (.ZN (n_104_23), .A (n_103_22), .B (n_104_20), .C1 (n_108_18), .C2 (n_111_18) );
AOI211_X1 g_102_22 (.ZN (n_102_22), .A (n_105_21), .B (n_102_21), .C1 (n_106_19), .C2 (n_109_19) );
AOI211_X1 g_104_21 (.ZN (n_104_21), .A (n_104_23), .B (n_101_23), .C1 (n_104_20), .C2 (n_107_20) );
AOI211_X1 g_106_20 (.ZN (n_106_20), .A (n_102_22), .B (n_103_22), .C1 (n_102_21), .C2 (n_108_18) );
AOI211_X1 g_108_19 (.ZN (n_108_19), .A (n_104_21), .B (n_105_21), .C1 (n_101_23), .C2 (n_106_19) );
AOI211_X1 g_110_18 (.ZN (n_110_18), .A (n_106_20), .B (n_104_23), .C1 (n_103_22), .C2 (n_104_20) );
AOI211_X1 g_112_17 (.ZN (n_112_17), .A (n_108_19), .B (n_102_22), .C1 (n_105_21), .C2 (n_102_21) );
AOI211_X1 g_111_19 (.ZN (n_111_19), .A (n_110_18), .B (n_104_21), .C1 (n_104_23), .C2 (n_101_23) );
AOI211_X1 g_109_20 (.ZN (n_109_20), .A (n_112_17), .B (n_106_20), .C1 (n_102_22), .C2 (n_103_22) );
AOI211_X1 g_107_21 (.ZN (n_107_21), .A (n_111_19), .B (n_108_19), .C1 (n_104_21), .C2 (n_105_21) );
AOI211_X1 g_105_22 (.ZN (n_105_22), .A (n_109_20), .B (n_110_18), .C1 (n_106_20), .C2 (n_104_23) );
AOI211_X1 g_103_23 (.ZN (n_103_23), .A (n_107_21), .B (n_112_17), .C1 (n_108_19), .C2 (n_102_22) );
AOI211_X1 g_101_24 (.ZN (n_101_24), .A (n_105_22), .B (n_111_19), .C1 (n_110_18), .C2 (n_104_21) );
AOI211_X1 g_99_25 (.ZN (n_99_25), .A (n_103_23), .B (n_109_20), .C1 (n_112_17), .C2 (n_106_20) );
AOI211_X1 g_100_23 (.ZN (n_100_23), .A (n_101_24), .B (n_107_21), .C1 (n_111_19), .C2 (n_108_19) );
AOI211_X1 g_98_24 (.ZN (n_98_24), .A (n_99_25), .B (n_105_22), .C1 (n_109_20), .C2 (n_110_18) );
AOI211_X1 g_97_26 (.ZN (n_97_26), .A (n_100_23), .B (n_103_23), .C1 (n_107_21), .C2 (n_112_17) );
AOI211_X1 g_95_27 (.ZN (n_95_27), .A (n_98_24), .B (n_101_24), .C1 (n_105_22), .C2 (n_111_19) );
AOI211_X1 g_96_25 (.ZN (n_96_25), .A (n_97_26), .B (n_99_25), .C1 (n_103_23), .C2 (n_109_20) );
AOI211_X1 g_94_24 (.ZN (n_94_24), .A (n_95_27), .B (n_100_23), .C1 (n_101_24), .C2 (n_107_21) );
AOI211_X1 g_93_26 (.ZN (n_93_26), .A (n_96_25), .B (n_98_24), .C1 (n_99_25), .C2 (n_105_22) );
AOI211_X1 g_91_27 (.ZN (n_91_27), .A (n_94_24), .B (n_97_26), .C1 (n_100_23), .C2 (n_103_23) );
AOI211_X1 g_92_25 (.ZN (n_92_25), .A (n_93_26), .B (n_95_27), .C1 (n_98_24), .C2 (n_101_24) );
AOI211_X1 g_90_26 (.ZN (n_90_26), .A (n_91_27), .B (n_96_25), .C1 (n_97_26), .C2 (n_99_25) );
AOI211_X1 g_89_28 (.ZN (n_89_28), .A (n_92_25), .B (n_94_24), .C1 (n_95_27), .C2 (n_100_23) );
AOI211_X1 g_87_29 (.ZN (n_87_29), .A (n_90_26), .B (n_93_26), .C1 (n_96_25), .C2 (n_98_24) );
AOI211_X1 g_85_30 (.ZN (n_85_30), .A (n_89_28), .B (n_91_27), .C1 (n_94_24), .C2 (n_97_26) );
AOI211_X1 g_83_31 (.ZN (n_83_31), .A (n_87_29), .B (n_92_25), .C1 (n_93_26), .C2 (n_95_27) );
AOI211_X1 g_81_32 (.ZN (n_81_32), .A (n_85_30), .B (n_90_26), .C1 (n_91_27), .C2 (n_96_25) );
AOI211_X1 g_82_30 (.ZN (n_82_30), .A (n_83_31), .B (n_89_28), .C1 (n_92_25), .C2 (n_94_24) );
AOI211_X1 g_80_31 (.ZN (n_80_31), .A (n_81_32), .B (n_87_29), .C1 (n_90_26), .C2 (n_93_26) );
AOI211_X1 g_78_32 (.ZN (n_78_32), .A (n_82_30), .B (n_85_30), .C1 (n_89_28), .C2 (n_91_27) );
AOI211_X1 g_76_33 (.ZN (n_76_33), .A (n_80_31), .B (n_83_31), .C1 (n_87_29), .C2 (n_92_25) );
AOI211_X1 g_74_34 (.ZN (n_74_34), .A (n_78_32), .B (n_81_32), .C1 (n_85_30), .C2 (n_90_26) );
AOI211_X1 g_72_35 (.ZN (n_72_35), .A (n_76_33), .B (n_82_30), .C1 (n_83_31), .C2 (n_89_28) );
AOI211_X1 g_70_34 (.ZN (n_70_34), .A (n_74_34), .B (n_80_31), .C1 (n_81_32), .C2 (n_87_29) );
AOI211_X1 g_68_35 (.ZN (n_68_35), .A (n_72_35), .B (n_78_32), .C1 (n_82_30), .C2 (n_85_30) );
AOI211_X1 g_66_36 (.ZN (n_66_36), .A (n_70_34), .B (n_76_33), .C1 (n_80_31), .C2 (n_83_31) );
AOI211_X1 g_64_37 (.ZN (n_64_37), .A (n_68_35), .B (n_74_34), .C1 (n_78_32), .C2 (n_81_32) );
AOI211_X1 g_62_38 (.ZN (n_62_38), .A (n_66_36), .B (n_72_35), .C1 (n_76_33), .C2 (n_82_30) );
AOI211_X1 g_60_39 (.ZN (n_60_39), .A (n_64_37), .B (n_70_34), .C1 (n_74_34), .C2 (n_80_31) );
AOI211_X1 g_58_40 (.ZN (n_58_40), .A (n_62_38), .B (n_68_35), .C1 (n_72_35), .C2 (n_78_32) );
AOI211_X1 g_56_41 (.ZN (n_56_41), .A (n_60_39), .B (n_66_36), .C1 (n_70_34), .C2 (n_76_33) );
AOI211_X1 g_54_42 (.ZN (n_54_42), .A (n_58_40), .B (n_64_37), .C1 (n_68_35), .C2 (n_74_34) );
AOI211_X1 g_55_40 (.ZN (n_55_40), .A (n_56_41), .B (n_62_38), .C1 (n_66_36), .C2 (n_72_35) );
AOI211_X1 g_53_41 (.ZN (n_53_41), .A (n_54_42), .B (n_60_39), .C1 (n_64_37), .C2 (n_70_34) );
AOI211_X1 g_51_42 (.ZN (n_51_42), .A (n_55_40), .B (n_58_40), .C1 (n_62_38), .C2 (n_68_35) );
AOI211_X1 g_49_43 (.ZN (n_49_43), .A (n_53_41), .B (n_56_41), .C1 (n_60_39), .C2 (n_66_36) );
AOI211_X1 g_47_44 (.ZN (n_47_44), .A (n_51_42), .B (n_54_42), .C1 (n_58_40), .C2 (n_64_37) );
AOI211_X1 g_45_45 (.ZN (n_45_45), .A (n_49_43), .B (n_55_40), .C1 (n_56_41), .C2 (n_62_38) );
AOI211_X1 g_43_46 (.ZN (n_43_46), .A (n_47_44), .B (n_53_41), .C1 (n_54_42), .C2 (n_60_39) );
AOI211_X1 g_41_47 (.ZN (n_41_47), .A (n_45_45), .B (n_51_42), .C1 (n_55_40), .C2 (n_58_40) );
AOI211_X1 g_40_49 (.ZN (n_40_49), .A (n_43_46), .B (n_49_43), .C1 (n_53_41), .C2 (n_56_41) );
AOI211_X1 g_38_50 (.ZN (n_38_50), .A (n_41_47), .B (n_47_44), .C1 (n_51_42), .C2 (n_54_42) );
AOI211_X1 g_37_52 (.ZN (n_37_52), .A (n_40_49), .B (n_45_45), .C1 (n_49_43), .C2 (n_55_40) );
AOI211_X1 g_35_51 (.ZN (n_35_51), .A (n_38_50), .B (n_43_46), .C1 (n_47_44), .C2 (n_53_41) );
AOI211_X1 g_37_50 (.ZN (n_37_50), .A (n_37_52), .B (n_41_47), .C1 (n_45_45), .C2 (n_51_42) );
AOI211_X1 g_39_49 (.ZN (n_39_49), .A (n_35_51), .B (n_40_49), .C1 (n_43_46), .C2 (n_49_43) );
AOI211_X1 g_41_48 (.ZN (n_41_48), .A (n_37_50), .B (n_38_50), .C1 (n_41_47), .C2 (n_47_44) );
AOI211_X1 g_40_50 (.ZN (n_40_50), .A (n_39_49), .B (n_37_52), .C1 (n_40_49), .C2 (n_45_45) );
AOI211_X1 g_42_49 (.ZN (n_42_49), .A (n_41_48), .B (n_35_51), .C1 (n_38_50), .C2 (n_43_46) );
AOI211_X1 g_44_48 (.ZN (n_44_48), .A (n_40_50), .B (n_37_50), .C1 (n_37_52), .C2 (n_41_47) );
AOI211_X1 g_46_47 (.ZN (n_46_47), .A (n_42_49), .B (n_39_49), .C1 (n_35_51), .C2 (n_40_49) );
AOI211_X1 g_48_46 (.ZN (n_48_46), .A (n_44_48), .B (n_41_48), .C1 (n_37_50), .C2 (n_38_50) );
AOI211_X1 g_50_45 (.ZN (n_50_45), .A (n_46_47), .B (n_40_50), .C1 (n_39_49), .C2 (n_37_52) );
AOI211_X1 g_52_44 (.ZN (n_52_44), .A (n_48_46), .B (n_42_49), .C1 (n_41_48), .C2 (n_35_51) );
AOI211_X1 g_54_43 (.ZN (n_54_43), .A (n_50_45), .B (n_44_48), .C1 (n_40_50), .C2 (n_37_50) );
AOI211_X1 g_56_42 (.ZN (n_56_42), .A (n_52_44), .B (n_46_47), .C1 (n_42_49), .C2 (n_39_49) );
AOI211_X1 g_55_44 (.ZN (n_55_44), .A (n_54_43), .B (n_48_46), .C1 (n_44_48), .C2 (n_41_48) );
AOI211_X1 g_53_43 (.ZN (n_53_43), .A (n_56_42), .B (n_50_45), .C1 (n_46_47), .C2 (n_40_50) );
AOI211_X1 g_55_42 (.ZN (n_55_42), .A (n_55_44), .B (n_52_44), .C1 (n_48_46), .C2 (n_42_49) );
AOI211_X1 g_57_41 (.ZN (n_57_41), .A (n_53_43), .B (n_54_43), .C1 (n_50_45), .C2 (n_44_48) );
AOI211_X1 g_59_40 (.ZN (n_59_40), .A (n_55_42), .B (n_56_42), .C1 (n_52_44), .C2 (n_46_47) );
AOI211_X1 g_61_39 (.ZN (n_61_39), .A (n_57_41), .B (n_55_44), .C1 (n_54_43), .C2 (n_48_46) );
AOI211_X1 g_63_38 (.ZN (n_63_38), .A (n_59_40), .B (n_53_43), .C1 (n_56_42), .C2 (n_50_45) );
AOI211_X1 g_65_37 (.ZN (n_65_37), .A (n_61_39), .B (n_55_42), .C1 (n_55_44), .C2 (n_52_44) );
AOI211_X1 g_67_36 (.ZN (n_67_36), .A (n_63_38), .B (n_57_41), .C1 (n_53_43), .C2 (n_54_43) );
AOI211_X1 g_66_38 (.ZN (n_66_38), .A (n_65_37), .B (n_59_40), .C1 (n_55_42), .C2 (n_56_42) );
AOI211_X1 g_68_37 (.ZN (n_68_37), .A (n_67_36), .B (n_61_39), .C1 (n_57_41), .C2 (n_55_44) );
AOI211_X1 g_70_36 (.ZN (n_70_36), .A (n_66_38), .B (n_63_38), .C1 (n_59_40), .C2 (n_53_43) );
AOI211_X1 g_72_37 (.ZN (n_72_37), .A (n_68_37), .B (n_65_37), .C1 (n_61_39), .C2 (n_55_42) );
AOI211_X1 g_71_35 (.ZN (n_71_35), .A (n_70_36), .B (n_67_36), .C1 (n_63_38), .C2 (n_57_41) );
AOI211_X1 g_69_36 (.ZN (n_69_36), .A (n_72_37), .B (n_66_38), .C1 (n_65_37), .C2 (n_59_40) );
AOI211_X1 g_67_37 (.ZN (n_67_37), .A (n_71_35), .B (n_68_37), .C1 (n_67_36), .C2 (n_61_39) );
AOI211_X1 g_65_38 (.ZN (n_65_38), .A (n_69_36), .B (n_70_36), .C1 (n_66_38), .C2 (n_63_38) );
AOI211_X1 g_63_39 (.ZN (n_63_39), .A (n_67_37), .B (n_72_37), .C1 (n_68_37), .C2 (n_65_37) );
AOI211_X1 g_61_40 (.ZN (n_61_40), .A (n_65_38), .B (n_71_35), .C1 (n_70_36), .C2 (n_67_36) );
AOI211_X1 g_59_41 (.ZN (n_59_41), .A (n_63_39), .B (n_69_36), .C1 (n_72_37), .C2 (n_66_38) );
AOI211_X1 g_57_42 (.ZN (n_57_42), .A (n_61_40), .B (n_67_37), .C1 (n_71_35), .C2 (n_68_37) );
AOI211_X1 g_55_43 (.ZN (n_55_43), .A (n_59_41), .B (n_65_38), .C1 (n_69_36), .C2 (n_70_36) );
AOI211_X1 g_53_44 (.ZN (n_53_44), .A (n_57_42), .B (n_63_39), .C1 (n_67_37), .C2 (n_72_37) );
AOI211_X1 g_51_45 (.ZN (n_51_45), .A (n_55_43), .B (n_61_40), .C1 (n_65_38), .C2 (n_71_35) );
AOI211_X1 g_52_43 (.ZN (n_52_43), .A (n_53_44), .B (n_59_41), .C1 (n_63_39), .C2 (n_69_36) );
AOI211_X1 g_50_44 (.ZN (n_50_44), .A (n_51_45), .B (n_57_42), .C1 (n_61_40), .C2 (n_67_37) );
AOI211_X1 g_48_45 (.ZN (n_48_45), .A (n_52_43), .B (n_55_43), .C1 (n_59_41), .C2 (n_65_38) );
AOI211_X1 g_46_46 (.ZN (n_46_46), .A (n_50_44), .B (n_53_44), .C1 (n_57_42), .C2 (n_63_39) );
AOI211_X1 g_44_47 (.ZN (n_44_47), .A (n_48_45), .B (n_51_45), .C1 (n_55_43), .C2 (n_61_40) );
AOI211_X1 g_42_48 (.ZN (n_42_48), .A (n_46_46), .B (n_52_43), .C1 (n_53_44), .C2 (n_59_41) );
AOI211_X1 g_41_50 (.ZN (n_41_50), .A (n_44_47), .B (n_50_44), .C1 (n_51_45), .C2 (n_57_42) );
AOI211_X1 g_39_51 (.ZN (n_39_51), .A (n_42_48), .B (n_48_45), .C1 (n_52_43), .C2 (n_55_43) );
AOI211_X1 g_41_52 (.ZN (n_41_52), .A (n_41_50), .B (n_46_46), .C1 (n_50_44), .C2 (n_53_44) );
AOI211_X1 g_43_51 (.ZN (n_43_51), .A (n_39_51), .B (n_44_47), .C1 (n_48_45), .C2 (n_51_45) );
AOI211_X1 g_44_49 (.ZN (n_44_49), .A (n_41_52), .B (n_42_48), .C1 (n_46_46), .C2 (n_52_43) );
AOI211_X1 g_45_47 (.ZN (n_45_47), .A (n_43_51), .B (n_41_50), .C1 (n_44_47), .C2 (n_50_44) );
AOI211_X1 g_47_46 (.ZN (n_47_46), .A (n_44_49), .B (n_39_51), .C1 (n_42_48), .C2 (n_48_45) );
AOI211_X1 g_49_45 (.ZN (n_49_45), .A (n_45_47), .B (n_41_52), .C1 (n_41_50), .C2 (n_46_46) );
AOI211_X1 g_51_44 (.ZN (n_51_44), .A (n_47_46), .B (n_43_51), .C1 (n_39_51), .C2 (n_44_47) );
AOI211_X1 g_53_45 (.ZN (n_53_45), .A (n_49_45), .B (n_44_49), .C1 (n_41_52), .C2 (n_42_48) );
AOI211_X1 g_51_46 (.ZN (n_51_46), .A (n_51_44), .B (n_45_47), .C1 (n_43_51), .C2 (n_41_50) );
AOI211_X1 g_49_47 (.ZN (n_49_47), .A (n_53_45), .B (n_47_46), .C1 (n_44_49), .C2 (n_39_51) );
AOI211_X1 g_47_48 (.ZN (n_47_48), .A (n_51_46), .B (n_49_45), .C1 (n_45_47), .C2 (n_41_52) );
AOI211_X1 g_45_49 (.ZN (n_45_49), .A (n_49_47), .B (n_51_44), .C1 (n_47_46), .C2 (n_43_51) );
AOI211_X1 g_43_48 (.ZN (n_43_48), .A (n_47_48), .B (n_53_45), .C1 (n_49_45), .C2 (n_44_49) );
AOI211_X1 g_42_50 (.ZN (n_42_50), .A (n_45_49), .B (n_51_46), .C1 (n_51_44), .C2 (n_45_47) );
AOI211_X1 g_40_51 (.ZN (n_40_51), .A (n_43_48), .B (n_49_47), .C1 (n_53_45), .C2 (n_47_46) );
AOI211_X1 g_41_49 (.ZN (n_41_49), .A (n_42_50), .B (n_47_48), .C1 (n_51_46), .C2 (n_49_45) );
AOI211_X1 g_39_50 (.ZN (n_39_50), .A (n_40_51), .B (n_45_49), .C1 (n_49_47), .C2 (n_51_44) );
AOI211_X1 g_37_51 (.ZN (n_37_51), .A (n_41_49), .B (n_43_48), .C1 (n_47_48), .C2 (n_53_45) );
AOI211_X1 g_35_52 (.ZN (n_35_52), .A (n_39_50), .B (n_42_50), .C1 (n_45_49), .C2 (n_51_46) );
AOI211_X1 g_33_53 (.ZN (n_33_53), .A (n_37_51), .B (n_40_51), .C1 (n_43_48), .C2 (n_49_47) );
AOI211_X1 g_31_52 (.ZN (n_31_52), .A (n_35_52), .B (n_41_49), .C1 (n_42_50), .C2 (n_47_48) );
AOI211_X1 g_30_54 (.ZN (n_30_54), .A (n_33_53), .B (n_39_50), .C1 (n_40_51), .C2 (n_45_49) );
AOI211_X1 g_28_55 (.ZN (n_28_55), .A (n_31_52), .B (n_37_51), .C1 (n_41_49), .C2 (n_43_48) );
AOI211_X1 g_29_53 (.ZN (n_29_53), .A (n_30_54), .B (n_35_52), .C1 (n_39_50), .C2 (n_42_50) );
AOI211_X1 g_27_54 (.ZN (n_27_54), .A (n_28_55), .B (n_33_53), .C1 (n_37_51), .C2 (n_40_51) );
AOI211_X1 g_25_55 (.ZN (n_25_55), .A (n_29_53), .B (n_31_52), .C1 (n_35_52), .C2 (n_41_49) );
AOI211_X1 g_23_56 (.ZN (n_23_56), .A (n_27_54), .B (n_30_54), .C1 (n_33_53), .C2 (n_39_50) );
AOI211_X1 g_21_57 (.ZN (n_21_57), .A (n_25_55), .B (n_28_55), .C1 (n_31_52), .C2 (n_37_51) );
AOI211_X1 g_19_58 (.ZN (n_19_58), .A (n_23_56), .B (n_29_53), .C1 (n_30_54), .C2 (n_35_52) );
AOI211_X1 g_18_60 (.ZN (n_18_60), .A (n_21_57), .B (n_27_54), .C1 (n_28_55), .C2 (n_33_53) );
AOI211_X1 g_20_59 (.ZN (n_20_59), .A (n_19_58), .B (n_25_55), .C1 (n_29_53), .C2 (n_31_52) );
AOI211_X1 g_22_58 (.ZN (n_22_58), .A (n_18_60), .B (n_23_56), .C1 (n_27_54), .C2 (n_30_54) );
AOI211_X1 g_24_57 (.ZN (n_24_57), .A (n_20_59), .B (n_21_57), .C1 (n_25_55), .C2 (n_28_55) );
AOI211_X1 g_26_56 (.ZN (n_26_56), .A (n_22_58), .B (n_19_58), .C1 (n_23_56), .C2 (n_29_53) );
AOI211_X1 g_25_58 (.ZN (n_25_58), .A (n_24_57), .B (n_18_60), .C1 (n_21_57), .C2 (n_27_54) );
AOI211_X1 g_27_57 (.ZN (n_27_57), .A (n_26_56), .B (n_20_59), .C1 (n_19_58), .C2 (n_25_55) );
AOI211_X1 g_26_55 (.ZN (n_26_55), .A (n_25_58), .B (n_22_58), .C1 (n_18_60), .C2 (n_23_56) );
AOI211_X1 g_24_56 (.ZN (n_24_56), .A (n_27_57), .B (n_24_57), .C1 (n_20_59), .C2 (n_21_57) );
AOI211_X1 g_22_57 (.ZN (n_22_57), .A (n_26_55), .B (n_26_56), .C1 (n_22_58), .C2 (n_19_58) );
AOI211_X1 g_21_59 (.ZN (n_21_59), .A (n_24_56), .B (n_25_58), .C1 (n_24_57), .C2 (n_18_60) );
AOI211_X1 g_23_58 (.ZN (n_23_58), .A (n_22_57), .B (n_27_57), .C1 (n_26_56), .C2 (n_20_59) );
AOI211_X1 g_25_57 (.ZN (n_25_57), .A (n_21_59), .B (n_26_55), .C1 (n_25_58), .C2 (n_22_58) );
AOI211_X1 g_27_56 (.ZN (n_27_56), .A (n_23_58), .B (n_24_56), .C1 (n_27_57), .C2 (n_24_57) );
AOI211_X1 g_29_55 (.ZN (n_29_55), .A (n_25_57), .B (n_22_57), .C1 (n_26_55), .C2 (n_26_56) );
AOI211_X1 g_31_54 (.ZN (n_31_54), .A (n_27_56), .B (n_21_59), .C1 (n_24_56), .C2 (n_25_58) );
AOI211_X1 g_30_56 (.ZN (n_30_56), .A (n_29_55), .B (n_23_58), .C1 (n_22_57), .C2 (n_27_57) );
AOI211_X1 g_28_57 (.ZN (n_28_57), .A (n_31_54), .B (n_25_57), .C1 (n_21_59), .C2 (n_26_55) );
AOI211_X1 g_26_58 (.ZN (n_26_58), .A (n_30_56), .B (n_27_56), .C1 (n_23_58), .C2 (n_24_56) );
AOI211_X1 g_24_59 (.ZN (n_24_59), .A (n_28_57), .B (n_29_55), .C1 (n_25_57), .C2 (n_22_57) );
AOI211_X1 g_22_60 (.ZN (n_22_60), .A (n_26_58), .B (n_31_54), .C1 (n_27_56), .C2 (n_21_59) );
AOI211_X1 g_21_58 (.ZN (n_21_58), .A (n_24_59), .B (n_30_56), .C1 (n_29_55), .C2 (n_23_58) );
AOI211_X1 g_19_59 (.ZN (n_19_59), .A (n_22_60), .B (n_28_57), .C1 (n_31_54), .C2 (n_25_57) );
AOI211_X1 g_17_60 (.ZN (n_17_60), .A (n_21_58), .B (n_26_58), .C1 (n_30_56), .C2 (n_27_56) );
AOI211_X1 g_15_61 (.ZN (n_15_61), .A (n_19_59), .B (n_24_59), .C1 (n_28_57), .C2 (n_29_55) );
AOI211_X1 g_13_62 (.ZN (n_13_62), .A (n_17_60), .B (n_22_60), .C1 (n_26_58), .C2 (n_31_54) );
AOI211_X1 g_11_63 (.ZN (n_11_63), .A (n_15_61), .B (n_21_58), .C1 (n_24_59), .C2 (n_30_56) );
AOI211_X1 g_9_64 (.ZN (n_9_64), .A (n_13_62), .B (n_19_59), .C1 (n_22_60), .C2 (n_28_57) );
AOI211_X1 g_7_65 (.ZN (n_7_65), .A (n_11_63), .B (n_17_60), .C1 (n_21_58), .C2 (n_26_58) );
AOI211_X1 g_5_66 (.ZN (n_5_66), .A (n_9_64), .B (n_15_61), .C1 (n_19_59), .C2 (n_24_59) );
AOI211_X1 g_3_67 (.ZN (n_3_67), .A (n_7_65), .B (n_13_62), .C1 (n_17_60), .C2 (n_22_60) );
AOI211_X1 g_1_68 (.ZN (n_1_68), .A (n_5_66), .B (n_11_63), .C1 (n_15_61), .C2 (n_21_58) );
AOI211_X1 g_2_66 (.ZN (n_2_66), .A (n_3_67), .B (n_9_64), .C1 (n_13_62), .C2 (n_19_59) );
AOI211_X1 g_3_64 (.ZN (n_3_64), .A (n_1_68), .B (n_7_65), .C1 (n_11_63), .C2 (n_17_60) );
AOI211_X1 g_5_63 (.ZN (n_5_63), .A (n_2_66), .B (n_5_66), .C1 (n_9_64), .C2 (n_15_61) );
AOI211_X1 g_4_65 (.ZN (n_4_65), .A (n_3_64), .B (n_3_67), .C1 (n_7_65), .C2 (n_13_62) );
AOI211_X1 g_5_67 (.ZN (n_5_67), .A (n_5_63), .B (n_1_68), .C1 (n_5_66), .C2 (n_11_63) );
AOI211_X1 g_3_68 (.ZN (n_3_68), .A (n_4_65), .B (n_2_66), .C1 (n_3_67), .C2 (n_9_64) );
AOI211_X1 g_4_66 (.ZN (n_4_66), .A (n_5_67), .B (n_3_64), .C1 (n_1_68), .C2 (n_7_65) );
AOI211_X1 g_6_67 (.ZN (n_6_67), .A (n_3_68), .B (n_5_63), .C1 (n_2_66), .C2 (n_5_66) );
AOI211_X1 g_8_66 (.ZN (n_8_66), .A (n_4_66), .B (n_4_65), .C1 (n_3_64), .C2 (n_3_67) );
AOI211_X1 g_7_64 (.ZN (n_7_64), .A (n_6_67), .B (n_5_67), .C1 (n_5_63), .C2 (n_1_68) );
AOI211_X1 g_9_65 (.ZN (n_9_65), .A (n_8_66), .B (n_3_68), .C1 (n_4_65), .C2 (n_2_66) );
AOI211_X1 g_11_64 (.ZN (n_11_64), .A (n_7_64), .B (n_4_66), .C1 (n_5_67), .C2 (n_3_64) );
AOI211_X1 g_13_63 (.ZN (n_13_63), .A (n_9_65), .B (n_6_67), .C1 (n_3_68), .C2 (n_5_63) );
AOI211_X1 g_15_62 (.ZN (n_15_62), .A (n_11_64), .B (n_8_66), .C1 (n_4_66), .C2 (n_4_65) );
AOI211_X1 g_17_61 (.ZN (n_17_61), .A (n_13_63), .B (n_7_64), .C1 (n_6_67), .C2 (n_5_67) );
AOI211_X1 g_19_60 (.ZN (n_19_60), .A (n_15_62), .B (n_9_65), .C1 (n_8_66), .C2 (n_3_68) );
AOI211_X1 g_18_62 (.ZN (n_18_62), .A (n_17_61), .B (n_11_64), .C1 (n_7_64), .C2 (n_4_66) );
AOI211_X1 g_20_61 (.ZN (n_20_61), .A (n_19_60), .B (n_13_63), .C1 (n_9_65), .C2 (n_6_67) );
AOI211_X1 g_19_63 (.ZN (n_19_63), .A (n_18_62), .B (n_15_62), .C1 (n_11_64), .C2 (n_8_66) );
AOI211_X1 g_18_61 (.ZN (n_18_61), .A (n_20_61), .B (n_17_61), .C1 (n_13_63), .C2 (n_7_64) );
AOI211_X1 g_20_60 (.ZN (n_20_60), .A (n_19_63), .B (n_19_60), .C1 (n_15_62), .C2 (n_9_65) );
AOI211_X1 g_22_59 (.ZN (n_22_59), .A (n_18_61), .B (n_18_62), .C1 (n_17_61), .C2 (n_11_64) );
AOI211_X1 g_24_58 (.ZN (n_24_58), .A (n_20_60), .B (n_20_61), .C1 (n_19_60), .C2 (n_13_63) );
AOI211_X1 g_26_57 (.ZN (n_26_57), .A (n_22_59), .B (n_19_63), .C1 (n_18_62), .C2 (n_15_62) );
AOI211_X1 g_28_56 (.ZN (n_28_56), .A (n_24_58), .B (n_18_61), .C1 (n_20_61), .C2 (n_17_61) );
AOI211_X1 g_30_55 (.ZN (n_30_55), .A (n_26_57), .B (n_20_60), .C1 (n_19_63), .C2 (n_19_60) );
AOI211_X1 g_31_53 (.ZN (n_31_53), .A (n_28_56), .B (n_22_59), .C1 (n_18_61), .C2 (n_18_62) );
AOI211_X1 g_33_52 (.ZN (n_33_52), .A (n_30_55), .B (n_24_58), .C1 (n_20_60), .C2 (n_20_61) );
AOI211_X1 g_32_54 (.ZN (n_32_54), .A (n_31_53), .B (n_26_57), .C1 (n_22_59), .C2 (n_19_63) );
AOI211_X1 g_34_53 (.ZN (n_34_53), .A (n_33_52), .B (n_28_56), .C1 (n_24_58), .C2 (n_18_61) );
AOI211_X1 g_36_52 (.ZN (n_36_52), .A (n_32_54), .B (n_30_55), .C1 (n_26_57), .C2 (n_20_60) );
AOI211_X1 g_38_51 (.ZN (n_38_51), .A (n_34_53), .B (n_31_53), .C1 (n_28_56), .C2 (n_22_59) );
AOI211_X1 g_39_53 (.ZN (n_39_53), .A (n_36_52), .B (n_33_52), .C1 (n_30_55), .C2 (n_24_58) );
AOI211_X1 g_37_54 (.ZN (n_37_54), .A (n_38_51), .B (n_32_54), .C1 (n_31_53), .C2 (n_26_57) );
AOI211_X1 g_38_52 (.ZN (n_38_52), .A (n_39_53), .B (n_34_53), .C1 (n_33_52), .C2 (n_28_56) );
AOI211_X1 g_36_53 (.ZN (n_36_53), .A (n_37_54), .B (n_36_52), .C1 (n_32_54), .C2 (n_30_55) );
AOI211_X1 g_34_54 (.ZN (n_34_54), .A (n_38_52), .B (n_38_51), .C1 (n_34_53), .C2 (n_31_53) );
AOI211_X1 g_32_55 (.ZN (n_32_55), .A (n_36_53), .B (n_39_53), .C1 (n_36_52), .C2 (n_33_52) );
AOI211_X1 g_31_57 (.ZN (n_31_57), .A (n_34_54), .B (n_37_54), .C1 (n_38_51), .C2 (n_32_54) );
AOI211_X1 g_33_56 (.ZN (n_33_56), .A (n_32_55), .B (n_38_52), .C1 (n_39_53), .C2 (n_34_53) );
AOI211_X1 g_35_55 (.ZN (n_35_55), .A (n_31_57), .B (n_36_53), .C1 (n_37_54), .C2 (n_36_52) );
AOI211_X1 g_33_54 (.ZN (n_33_54), .A (n_33_56), .B (n_34_54), .C1 (n_38_52), .C2 (n_38_51) );
AOI211_X1 g_35_53 (.ZN (n_35_53), .A (n_35_55), .B (n_32_55), .C1 (n_36_53), .C2 (n_39_53) );
AOI211_X1 g_34_55 (.ZN (n_34_55), .A (n_33_54), .B (n_31_57), .C1 (n_34_54), .C2 (n_37_54) );
AOI211_X1 g_36_54 (.ZN (n_36_54), .A (n_35_53), .B (n_33_56), .C1 (n_32_55), .C2 (n_38_52) );
AOI211_X1 g_38_53 (.ZN (n_38_53), .A (n_34_55), .B (n_35_55), .C1 (n_31_57), .C2 (n_36_53) );
AOI211_X1 g_40_52 (.ZN (n_40_52), .A (n_36_54), .B (n_33_54), .C1 (n_33_56), .C2 (n_34_54) );
AOI211_X1 g_42_51 (.ZN (n_42_51), .A (n_38_53), .B (n_35_53), .C1 (n_35_55), .C2 (n_32_55) );
AOI211_X1 g_43_49 (.ZN (n_43_49), .A (n_40_52), .B (n_34_55), .C1 (n_33_54), .C2 (n_31_57) );
AOI211_X1 g_45_48 (.ZN (n_45_48), .A (n_42_51), .B (n_36_54), .C1 (n_35_53), .C2 (n_33_56) );
AOI211_X1 g_47_47 (.ZN (n_47_47), .A (n_43_49), .B (n_38_53), .C1 (n_34_55), .C2 (n_35_55) );
AOI211_X1 g_49_46 (.ZN (n_49_46), .A (n_45_48), .B (n_40_52), .C1 (n_36_54), .C2 (n_33_54) );
AOI211_X1 g_48_48 (.ZN (n_48_48), .A (n_47_47), .B (n_42_51), .C1 (n_38_53), .C2 (n_35_53) );
AOI211_X1 g_50_47 (.ZN (n_50_47), .A (n_49_46), .B (n_43_49), .C1 (n_40_52), .C2 (n_34_55) );
AOI211_X1 g_52_46 (.ZN (n_52_46), .A (n_48_48), .B (n_45_48), .C1 (n_42_51), .C2 (n_36_54) );
AOI211_X1 g_54_45 (.ZN (n_54_45), .A (n_50_47), .B (n_47_47), .C1 (n_43_49), .C2 (n_38_53) );
AOI211_X1 g_56_44 (.ZN (n_56_44), .A (n_52_46), .B (n_49_46), .C1 (n_45_48), .C2 (n_40_52) );
AOI211_X1 g_58_43 (.ZN (n_58_43), .A (n_54_45), .B (n_48_48), .C1 (n_47_47), .C2 (n_42_51) );
AOI211_X1 g_60_42 (.ZN (n_60_42), .A (n_56_44), .B (n_50_47), .C1 (n_49_46), .C2 (n_43_49) );
AOI211_X1 g_62_41 (.ZN (n_62_41), .A (n_58_43), .B (n_52_46), .C1 (n_48_48), .C2 (n_45_48) );
AOI211_X1 g_64_40 (.ZN (n_64_40), .A (n_60_42), .B (n_54_45), .C1 (n_50_47), .C2 (n_47_47) );
AOI211_X1 g_66_39 (.ZN (n_66_39), .A (n_62_41), .B (n_56_44), .C1 (n_52_46), .C2 (n_49_46) );
AOI211_X1 g_68_38 (.ZN (n_68_38), .A (n_64_40), .B (n_58_43), .C1 (n_54_45), .C2 (n_48_48) );
AOI211_X1 g_70_37 (.ZN (n_70_37), .A (n_66_39), .B (n_60_42), .C1 (n_56_44), .C2 (n_50_47) );
AOI211_X1 g_72_36 (.ZN (n_72_36), .A (n_68_38), .B (n_62_41), .C1 (n_58_43), .C2 (n_52_46) );
AOI211_X1 g_74_35 (.ZN (n_74_35), .A (n_70_37), .B (n_64_40), .C1 (n_60_42), .C2 (n_54_45) );
AOI211_X1 g_76_34 (.ZN (n_76_34), .A (n_72_36), .B (n_66_39), .C1 (n_62_41), .C2 (n_56_44) );
AOI211_X1 g_78_33 (.ZN (n_78_33), .A (n_74_35), .B (n_68_38), .C1 (n_64_40), .C2 (n_58_43) );
AOI211_X1 g_80_32 (.ZN (n_80_32), .A (n_76_34), .B (n_70_37), .C1 (n_66_39), .C2 (n_60_42) );
AOI211_X1 g_82_31 (.ZN (n_82_31), .A (n_78_33), .B (n_72_36), .C1 (n_68_38), .C2 (n_62_41) );
AOI211_X1 g_84_30 (.ZN (n_84_30), .A (n_80_32), .B (n_74_35), .C1 (n_70_37), .C2 (n_64_40) );
AOI211_X1 g_83_32 (.ZN (n_83_32), .A (n_82_31), .B (n_76_34), .C1 (n_72_36), .C2 (n_66_39) );
AOI211_X1 g_81_31 (.ZN (n_81_31), .A (n_84_30), .B (n_78_33), .C1 (n_74_35), .C2 (n_68_38) );
AOI211_X1 g_83_30 (.ZN (n_83_30), .A (n_83_32), .B (n_80_32), .C1 (n_76_34), .C2 (n_70_37) );
AOI211_X1 g_85_29 (.ZN (n_85_29), .A (n_81_31), .B (n_82_31), .C1 (n_78_33), .C2 (n_72_36) );
AOI211_X1 g_87_28 (.ZN (n_87_28), .A (n_83_30), .B (n_84_30), .C1 (n_80_32), .C2 (n_74_35) );
AOI211_X1 g_89_27 (.ZN (n_89_27), .A (n_85_29), .B (n_83_32), .C1 (n_82_31), .C2 (n_76_34) );
AOI211_X1 g_91_26 (.ZN (n_91_26), .A (n_87_28), .B (n_81_31), .C1 (n_84_30), .C2 (n_78_33) );
AOI211_X1 g_93_25 (.ZN (n_93_25), .A (n_89_27), .B (n_83_30), .C1 (n_83_32), .C2 (n_80_32) );
AOI211_X1 g_94_27 (.ZN (n_94_27), .A (n_91_26), .B (n_85_29), .C1 (n_81_31), .C2 (n_82_31) );
AOI211_X1 g_92_28 (.ZN (n_92_28), .A (n_93_25), .B (n_87_28), .C1 (n_83_30), .C2 (n_84_30) );
AOI211_X1 g_90_29 (.ZN (n_90_29), .A (n_94_27), .B (n_89_27), .C1 (n_85_29), .C2 (n_83_32) );
AOI211_X1 g_88_30 (.ZN (n_88_30), .A (n_92_28), .B (n_91_26), .C1 (n_87_28), .C2 (n_81_31) );
AOI211_X1 g_86_31 (.ZN (n_86_31), .A (n_90_29), .B (n_93_25), .C1 (n_89_27), .C2 (n_83_30) );
AOI211_X1 g_84_32 (.ZN (n_84_32), .A (n_88_30), .B (n_94_27), .C1 (n_91_26), .C2 (n_85_29) );
AOI211_X1 g_82_33 (.ZN (n_82_33), .A (n_86_31), .B (n_92_28), .C1 (n_93_25), .C2 (n_87_28) );
AOI211_X1 g_80_34 (.ZN (n_80_34), .A (n_84_32), .B (n_90_29), .C1 (n_94_27), .C2 (n_89_27) );
AOI211_X1 g_78_35 (.ZN (n_78_35), .A (n_82_33), .B (n_88_30), .C1 (n_92_28), .C2 (n_91_26) );
AOI211_X1 g_79_33 (.ZN (n_79_33), .A (n_80_34), .B (n_86_31), .C1 (n_90_29), .C2 (n_93_25) );
AOI211_X1 g_77_34 (.ZN (n_77_34), .A (n_78_35), .B (n_84_32), .C1 (n_88_30), .C2 (n_94_27) );
AOI211_X1 g_75_35 (.ZN (n_75_35), .A (n_79_33), .B (n_82_33), .C1 (n_86_31), .C2 (n_92_28) );
AOI211_X1 g_73_36 (.ZN (n_73_36), .A (n_77_34), .B (n_80_34), .C1 (n_84_32), .C2 (n_90_29) );
AOI211_X1 g_71_37 (.ZN (n_71_37), .A (n_75_35), .B (n_78_35), .C1 (n_82_33), .C2 (n_88_30) );
AOI211_X1 g_69_38 (.ZN (n_69_38), .A (n_73_36), .B (n_79_33), .C1 (n_80_34), .C2 (n_86_31) );
AOI211_X1 g_67_39 (.ZN (n_67_39), .A (n_71_37), .B (n_77_34), .C1 (n_78_35), .C2 (n_84_32) );
AOI211_X1 g_65_40 (.ZN (n_65_40), .A (n_69_38), .B (n_75_35), .C1 (n_79_33), .C2 (n_82_33) );
AOI211_X1 g_63_41 (.ZN (n_63_41), .A (n_67_39), .B (n_73_36), .C1 (n_77_34), .C2 (n_80_34) );
AOI211_X1 g_64_39 (.ZN (n_64_39), .A (n_65_40), .B (n_71_37), .C1 (n_75_35), .C2 (n_78_35) );
AOI211_X1 g_62_40 (.ZN (n_62_40), .A (n_63_41), .B (n_69_38), .C1 (n_73_36), .C2 (n_79_33) );
AOI211_X1 g_60_41 (.ZN (n_60_41), .A (n_64_39), .B (n_67_39), .C1 (n_71_37), .C2 (n_77_34) );
AOI211_X1 g_58_42 (.ZN (n_58_42), .A (n_62_40), .B (n_65_40), .C1 (n_69_38), .C2 (n_75_35) );
AOI211_X1 g_56_43 (.ZN (n_56_43), .A (n_60_41), .B (n_63_41), .C1 (n_67_39), .C2 (n_73_36) );
AOI211_X1 g_54_44 (.ZN (n_54_44), .A (n_58_42), .B (n_64_39), .C1 (n_65_40), .C2 (n_71_37) );
AOI211_X1 g_52_45 (.ZN (n_52_45), .A (n_56_43), .B (n_62_40), .C1 (n_63_41), .C2 (n_69_38) );
AOI211_X1 g_50_46 (.ZN (n_50_46), .A (n_54_44), .B (n_60_41), .C1 (n_64_39), .C2 (n_67_39) );
AOI211_X1 g_48_47 (.ZN (n_48_47), .A (n_52_45), .B (n_58_42), .C1 (n_62_40), .C2 (n_65_40) );
AOI211_X1 g_46_48 (.ZN (n_46_48), .A (n_50_46), .B (n_56_43), .C1 (n_60_41), .C2 (n_63_41) );
AOI211_X1 g_45_50 (.ZN (n_45_50), .A (n_48_47), .B (n_54_44), .C1 (n_58_42), .C2 (n_64_39) );
AOI211_X1 g_47_49 (.ZN (n_47_49), .A (n_46_48), .B (n_52_45), .C1 (n_56_43), .C2 (n_62_40) );
AOI211_X1 g_49_48 (.ZN (n_49_48), .A (n_45_50), .B (n_50_46), .C1 (n_54_44), .C2 (n_60_41) );
AOI211_X1 g_51_47 (.ZN (n_51_47), .A (n_47_49), .B (n_48_47), .C1 (n_52_45), .C2 (n_58_42) );
AOI211_X1 g_53_46 (.ZN (n_53_46), .A (n_49_48), .B (n_46_48), .C1 (n_50_46), .C2 (n_56_43) );
AOI211_X1 g_55_45 (.ZN (n_55_45), .A (n_51_47), .B (n_45_50), .C1 (n_48_47), .C2 (n_54_44) );
AOI211_X1 g_57_44 (.ZN (n_57_44), .A (n_53_46), .B (n_47_49), .C1 (n_46_48), .C2 (n_52_45) );
AOI211_X1 g_59_43 (.ZN (n_59_43), .A (n_55_45), .B (n_49_48), .C1 (n_45_50), .C2 (n_50_46) );
AOI211_X1 g_61_42 (.ZN (n_61_42), .A (n_57_44), .B (n_51_47), .C1 (n_47_49), .C2 (n_48_47) );
AOI211_X1 g_60_44 (.ZN (n_60_44), .A (n_59_43), .B (n_53_46), .C1 (n_49_48), .C2 (n_46_48) );
AOI211_X1 g_59_42 (.ZN (n_59_42), .A (n_61_42), .B (n_55_45), .C1 (n_51_47), .C2 (n_45_50) );
AOI211_X1 g_57_43 (.ZN (n_57_43), .A (n_60_44), .B (n_57_44), .C1 (n_53_46), .C2 (n_47_49) );
AOI211_X1 g_58_45 (.ZN (n_58_45), .A (n_59_42), .B (n_59_43), .C1 (n_55_45), .C2 (n_49_48) );
AOI211_X1 g_56_46 (.ZN (n_56_46), .A (n_57_43), .B (n_61_42), .C1 (n_57_44), .C2 (n_51_47) );
AOI211_X1 g_54_47 (.ZN (n_54_47), .A (n_58_45), .B (n_60_44), .C1 (n_59_43), .C2 (n_53_46) );
AOI211_X1 g_52_48 (.ZN (n_52_48), .A (n_56_46), .B (n_59_42), .C1 (n_61_42), .C2 (n_55_45) );
AOI211_X1 g_50_49 (.ZN (n_50_49), .A (n_54_47), .B (n_57_43), .C1 (n_60_44), .C2 (n_57_44) );
AOI211_X1 g_48_50 (.ZN (n_48_50), .A (n_52_48), .B (n_58_45), .C1 (n_59_42), .C2 (n_59_43) );
AOI211_X1 g_46_49 (.ZN (n_46_49), .A (n_50_49), .B (n_56_46), .C1 (n_57_43), .C2 (n_61_42) );
AOI211_X1 g_44_50 (.ZN (n_44_50), .A (n_48_50), .B (n_54_47), .C1 (n_58_45), .C2 (n_60_44) );
AOI211_X1 g_46_51 (.ZN (n_46_51), .A (n_46_49), .B (n_52_48), .C1 (n_56_46), .C2 (n_59_42) );
AOI211_X1 g_44_52 (.ZN (n_44_52), .A (n_44_50), .B (n_50_49), .C1 (n_54_47), .C2 (n_57_43) );
AOI211_X1 g_43_50 (.ZN (n_43_50), .A (n_46_51), .B (n_48_50), .C1 (n_52_48), .C2 (n_58_45) );
AOI211_X1 g_41_51 (.ZN (n_41_51), .A (n_44_52), .B (n_46_49), .C1 (n_50_49), .C2 (n_56_46) );
AOI211_X1 g_39_52 (.ZN (n_39_52), .A (n_43_50), .B (n_44_50), .C1 (n_48_50), .C2 (n_54_47) );
AOI211_X1 g_37_53 (.ZN (n_37_53), .A (n_41_51), .B (n_46_51), .C1 (n_46_49), .C2 (n_52_48) );
AOI211_X1 g_35_54 (.ZN (n_35_54), .A (n_39_52), .B (n_44_52), .C1 (n_44_50), .C2 (n_50_49) );
AOI211_X1 g_33_55 (.ZN (n_33_55), .A (n_37_53), .B (n_43_50), .C1 (n_46_51), .C2 (n_48_50) );
AOI211_X1 g_31_56 (.ZN (n_31_56), .A (n_35_54), .B (n_41_51), .C1 (n_44_52), .C2 (n_46_49) );
AOI211_X1 g_29_57 (.ZN (n_29_57), .A (n_33_55), .B (n_39_52), .C1 (n_43_50), .C2 (n_44_50) );
AOI211_X1 g_27_58 (.ZN (n_27_58), .A (n_31_56), .B (n_37_53), .C1 (n_41_51), .C2 (n_46_51) );
AOI211_X1 g_25_59 (.ZN (n_25_59), .A (n_29_57), .B (n_35_54), .C1 (n_39_52), .C2 (n_44_52) );
AOI211_X1 g_23_60 (.ZN (n_23_60), .A (n_27_58), .B (n_33_55), .C1 (n_37_53), .C2 (n_43_50) );
AOI211_X1 g_21_61 (.ZN (n_21_61), .A (n_25_59), .B (n_31_56), .C1 (n_35_54), .C2 (n_41_51) );
AOI211_X1 g_19_62 (.ZN (n_19_62), .A (n_23_60), .B (n_29_57), .C1 (n_33_55), .C2 (n_39_52) );
AOI211_X1 g_17_63 (.ZN (n_17_63), .A (n_21_61), .B (n_27_58), .C1 (n_31_56), .C2 (n_37_53) );
AOI211_X1 g_16_61 (.ZN (n_16_61), .A (n_19_62), .B (n_25_59), .C1 (n_29_57), .C2 (n_35_54) );
AOI211_X1 g_14_62 (.ZN (n_14_62), .A (n_17_63), .B (n_23_60), .C1 (n_27_58), .C2 (n_33_55) );
AOI211_X1 g_12_63 (.ZN (n_12_63), .A (n_16_61), .B (n_21_61), .C1 (n_25_59), .C2 (n_31_56) );
AOI211_X1 g_10_64 (.ZN (n_10_64), .A (n_14_62), .B (n_19_62), .C1 (n_23_60), .C2 (n_29_57) );
AOI211_X1 g_8_65 (.ZN (n_8_65), .A (n_12_63), .B (n_17_63), .C1 (n_21_61), .C2 (n_27_58) );
AOI211_X1 g_6_66 (.ZN (n_6_66), .A (n_10_64), .B (n_16_61), .C1 (n_19_62), .C2 (n_25_59) );
AOI211_X1 g_4_67 (.ZN (n_4_67), .A (n_8_65), .B (n_14_62), .C1 (n_17_63), .C2 (n_23_60) );
AOI211_X1 g_3_69 (.ZN (n_3_69), .A (n_6_66), .B (n_12_63), .C1 (n_16_61), .C2 (n_21_61) );
AOI211_X1 g_5_68 (.ZN (n_5_68), .A (n_4_67), .B (n_10_64), .C1 (n_14_62), .C2 (n_19_62) );
AOI211_X1 g_7_67 (.ZN (n_7_67), .A (n_3_69), .B (n_8_65), .C1 (n_12_63), .C2 (n_17_63) );
AOI211_X1 g_9_66 (.ZN (n_9_66), .A (n_5_68), .B (n_6_66), .C1 (n_10_64), .C2 (n_16_61) );
AOI211_X1 g_11_65 (.ZN (n_11_65), .A (n_7_67), .B (n_4_67), .C1 (n_8_65), .C2 (n_14_62) );
AOI211_X1 g_13_64 (.ZN (n_13_64), .A (n_9_66), .B (n_3_69), .C1 (n_6_66), .C2 (n_12_63) );
AOI211_X1 g_15_63 (.ZN (n_15_63), .A (n_11_65), .B (n_5_68), .C1 (n_4_67), .C2 (n_10_64) );
AOI211_X1 g_17_62 (.ZN (n_17_62), .A (n_13_64), .B (n_7_67), .C1 (n_3_69), .C2 (n_8_65) );
AOI211_X1 g_19_61 (.ZN (n_19_61), .A (n_15_63), .B (n_9_66), .C1 (n_5_68), .C2 (n_6_66) );
AOI211_X1 g_21_60 (.ZN (n_21_60), .A (n_17_62), .B (n_11_65), .C1 (n_7_67), .C2 (n_4_67) );
AOI211_X1 g_23_59 (.ZN (n_23_59), .A (n_19_61), .B (n_13_64), .C1 (n_9_66), .C2 (n_3_69) );
AOI211_X1 g_22_61 (.ZN (n_22_61), .A (n_21_60), .B (n_15_63), .C1 (n_11_65), .C2 (n_5_68) );
AOI211_X1 g_24_60 (.ZN (n_24_60), .A (n_23_59), .B (n_17_62), .C1 (n_13_64), .C2 (n_7_67) );
AOI211_X1 g_26_59 (.ZN (n_26_59), .A (n_22_61), .B (n_19_61), .C1 (n_15_63), .C2 (n_9_66) );
AOI211_X1 g_28_58 (.ZN (n_28_58), .A (n_24_60), .B (n_21_60), .C1 (n_17_62), .C2 (n_11_65) );
AOI211_X1 g_30_57 (.ZN (n_30_57), .A (n_26_59), .B (n_23_59), .C1 (n_19_61), .C2 (n_13_64) );
AOI211_X1 g_32_56 (.ZN (n_32_56), .A (n_28_58), .B (n_22_61), .C1 (n_21_60), .C2 (n_15_63) );
AOI211_X1 g_31_58 (.ZN (n_31_58), .A (n_30_57), .B (n_24_60), .C1 (n_23_59), .C2 (n_17_62) );
AOI211_X1 g_33_57 (.ZN (n_33_57), .A (n_32_56), .B (n_26_59), .C1 (n_22_61), .C2 (n_19_61) );
AOI211_X1 g_35_56 (.ZN (n_35_56), .A (n_31_58), .B (n_28_58), .C1 (n_24_60), .C2 (n_21_60) );
AOI211_X1 g_37_55 (.ZN (n_37_55), .A (n_33_57), .B (n_30_57), .C1 (n_26_59), .C2 (n_23_59) );
AOI211_X1 g_39_54 (.ZN (n_39_54), .A (n_35_56), .B (n_32_56), .C1 (n_28_58), .C2 (n_22_61) );
AOI211_X1 g_41_53 (.ZN (n_41_53), .A (n_37_55), .B (n_31_58), .C1 (n_30_57), .C2 (n_24_60) );
AOI211_X1 g_43_52 (.ZN (n_43_52), .A (n_39_54), .B (n_33_57), .C1 (n_32_56), .C2 (n_26_59) );
AOI211_X1 g_45_51 (.ZN (n_45_51), .A (n_41_53), .B (n_35_56), .C1 (n_31_58), .C2 (n_28_58) );
AOI211_X1 g_47_50 (.ZN (n_47_50), .A (n_43_52), .B (n_37_55), .C1 (n_33_57), .C2 (n_30_57) );
AOI211_X1 g_49_49 (.ZN (n_49_49), .A (n_45_51), .B (n_39_54), .C1 (n_35_56), .C2 (n_32_56) );
AOI211_X1 g_51_48 (.ZN (n_51_48), .A (n_47_50), .B (n_41_53), .C1 (n_37_55), .C2 (n_31_58) );
AOI211_X1 g_53_47 (.ZN (n_53_47), .A (n_49_49), .B (n_43_52), .C1 (n_39_54), .C2 (n_33_57) );
AOI211_X1 g_55_46 (.ZN (n_55_46), .A (n_51_48), .B (n_45_51), .C1 (n_41_53), .C2 (n_35_56) );
AOI211_X1 g_57_45 (.ZN (n_57_45), .A (n_53_47), .B (n_47_50), .C1 (n_43_52), .C2 (n_37_55) );
AOI211_X1 g_59_44 (.ZN (n_59_44), .A (n_55_46), .B (n_49_49), .C1 (n_45_51), .C2 (n_39_54) );
AOI211_X1 g_61_43 (.ZN (n_61_43), .A (n_57_45), .B (n_51_48), .C1 (n_47_50), .C2 (n_41_53) );
AOI211_X1 g_63_42 (.ZN (n_63_42), .A (n_59_44), .B (n_53_47), .C1 (n_49_49), .C2 (n_43_52) );
AOI211_X1 g_61_41 (.ZN (n_61_41), .A (n_61_43), .B (n_55_46), .C1 (n_51_48), .C2 (n_45_51) );
AOI211_X1 g_63_40 (.ZN (n_63_40), .A (n_63_42), .B (n_57_45), .C1 (n_53_47), .C2 (n_47_50) );
AOI211_X1 g_65_39 (.ZN (n_65_39), .A (n_61_41), .B (n_59_44), .C1 (n_55_46), .C2 (n_49_49) );
AOI211_X1 g_67_38 (.ZN (n_67_38), .A (n_63_40), .B (n_61_43), .C1 (n_57_45), .C2 (n_51_48) );
AOI211_X1 g_69_37 (.ZN (n_69_37), .A (n_65_39), .B (n_63_42), .C1 (n_59_44), .C2 (n_53_47) );
AOI211_X1 g_71_36 (.ZN (n_71_36), .A (n_67_38), .B (n_61_41), .C1 (n_61_43), .C2 (n_55_46) );
AOI211_X1 g_70_38 (.ZN (n_70_38), .A (n_69_37), .B (n_63_40), .C1 (n_63_42), .C2 (n_57_45) );
AOI211_X1 g_68_39 (.ZN (n_68_39), .A (n_71_36), .B (n_65_39), .C1 (n_61_41), .C2 (n_59_44) );
AOI211_X1 g_66_40 (.ZN (n_66_40), .A (n_70_38), .B (n_67_38), .C1 (n_63_40), .C2 (n_61_43) );
AOI211_X1 g_64_41 (.ZN (n_64_41), .A (n_68_39), .B (n_69_37), .C1 (n_65_39), .C2 (n_63_42) );
AOI211_X1 g_62_42 (.ZN (n_62_42), .A (n_66_40), .B (n_71_36), .C1 (n_67_38), .C2 (n_61_41) );
AOI211_X1 g_60_43 (.ZN (n_60_43), .A (n_64_41), .B (n_70_38), .C1 (n_69_37), .C2 (n_63_40) );
AOI211_X1 g_58_44 (.ZN (n_58_44), .A (n_62_42), .B (n_68_39), .C1 (n_71_36), .C2 (n_65_39) );
AOI211_X1 g_56_45 (.ZN (n_56_45), .A (n_60_43), .B (n_66_40), .C1 (n_70_38), .C2 (n_67_38) );
AOI211_X1 g_54_46 (.ZN (n_54_46), .A (n_58_44), .B (n_64_41), .C1 (n_68_39), .C2 (n_69_37) );
AOI211_X1 g_52_47 (.ZN (n_52_47), .A (n_56_45), .B (n_62_42), .C1 (n_66_40), .C2 (n_71_36) );
AOI211_X1 g_50_48 (.ZN (n_50_48), .A (n_54_46), .B (n_60_43), .C1 (n_64_41), .C2 (n_70_38) );
AOI211_X1 g_48_49 (.ZN (n_48_49), .A (n_52_47), .B (n_58_44), .C1 (n_62_42), .C2 (n_68_39) );
AOI211_X1 g_46_50 (.ZN (n_46_50), .A (n_50_48), .B (n_56_45), .C1 (n_60_43), .C2 (n_66_40) );
AOI211_X1 g_44_51 (.ZN (n_44_51), .A (n_48_49), .B (n_54_46), .C1 (n_58_44), .C2 (n_64_41) );
AOI211_X1 g_42_52 (.ZN (n_42_52), .A (n_46_50), .B (n_52_47), .C1 (n_56_45), .C2 (n_62_42) );
AOI211_X1 g_40_53 (.ZN (n_40_53), .A (n_44_51), .B (n_50_48), .C1 (n_54_46), .C2 (n_60_43) );
AOI211_X1 g_38_54 (.ZN (n_38_54), .A (n_42_52), .B (n_48_49), .C1 (n_52_47), .C2 (n_58_44) );
AOI211_X1 g_36_55 (.ZN (n_36_55), .A (n_40_53), .B (n_46_50), .C1 (n_50_48), .C2 (n_56_45) );
AOI211_X1 g_34_56 (.ZN (n_34_56), .A (n_38_54), .B (n_44_51), .C1 (n_48_49), .C2 (n_54_46) );
AOI211_X1 g_32_57 (.ZN (n_32_57), .A (n_36_55), .B (n_42_52), .C1 (n_46_50), .C2 (n_52_47) );
AOI211_X1 g_30_58 (.ZN (n_30_58), .A (n_34_56), .B (n_40_53), .C1 (n_44_51), .C2 (n_50_48) );
AOI211_X1 g_28_59 (.ZN (n_28_59), .A (n_32_57), .B (n_38_54), .C1 (n_42_52), .C2 (n_48_49) );
AOI211_X1 g_26_60 (.ZN (n_26_60), .A (n_30_58), .B (n_36_55), .C1 (n_40_53), .C2 (n_46_50) );
AOI211_X1 g_24_61 (.ZN (n_24_61), .A (n_28_59), .B (n_34_56), .C1 (n_38_54), .C2 (n_44_51) );
AOI211_X1 g_22_62 (.ZN (n_22_62), .A (n_26_60), .B (n_32_57), .C1 (n_36_55), .C2 (n_42_52) );
AOI211_X1 g_20_63 (.ZN (n_20_63), .A (n_24_61), .B (n_30_58), .C1 (n_34_56), .C2 (n_40_53) );
AOI211_X1 g_18_64 (.ZN (n_18_64), .A (n_22_62), .B (n_28_59), .C1 (n_32_57), .C2 (n_38_54) );
AOI211_X1 g_16_63 (.ZN (n_16_63), .A (n_20_63), .B (n_26_60), .C1 (n_30_58), .C2 (n_36_55) );
AOI211_X1 g_14_64 (.ZN (n_14_64), .A (n_18_64), .B (n_24_61), .C1 (n_28_59), .C2 (n_34_56) );
AOI211_X1 g_12_65 (.ZN (n_12_65), .A (n_16_63), .B (n_22_62), .C1 (n_26_60), .C2 (n_32_57) );
AOI211_X1 g_10_66 (.ZN (n_10_66), .A (n_14_64), .B (n_20_63), .C1 (n_24_61), .C2 (n_30_58) );
AOI211_X1 g_8_67 (.ZN (n_8_67), .A (n_12_65), .B (n_18_64), .C1 (n_22_62), .C2 (n_28_59) );
AOI211_X1 g_6_68 (.ZN (n_6_68), .A (n_10_66), .B (n_16_63), .C1 (n_20_63), .C2 (n_26_60) );
AOI211_X1 g_4_69 (.ZN (n_4_69), .A (n_8_67), .B (n_14_64), .C1 (n_18_64), .C2 (n_24_61) );
AOI211_X1 g_2_70 (.ZN (n_2_70), .A (n_6_68), .B (n_12_65), .C1 (n_16_63), .C2 (n_22_62) );
AOI211_X1 g_1_72 (.ZN (n_1_72), .A (n_4_69), .B (n_10_66), .C1 (n_14_64), .C2 (n_20_63) );
AOI211_X1 g_3_71 (.ZN (n_3_71), .A (n_2_70), .B (n_8_67), .C1 (n_12_65), .C2 (n_18_64) );
AOI211_X1 g_5_70 (.ZN (n_5_70), .A (n_1_72), .B (n_6_68), .C1 (n_10_66), .C2 (n_16_63) );
AOI211_X1 g_7_69 (.ZN (n_7_69), .A (n_3_71), .B (n_4_69), .C1 (n_8_67), .C2 (n_14_64) );
AOI211_X1 g_9_68 (.ZN (n_9_68), .A (n_5_70), .B (n_2_70), .C1 (n_6_68), .C2 (n_12_65) );
AOI211_X1 g_11_67 (.ZN (n_11_67), .A (n_7_69), .B (n_1_72), .C1 (n_4_69), .C2 (n_10_66) );
AOI211_X1 g_10_65 (.ZN (n_10_65), .A (n_9_68), .B (n_3_71), .C1 (n_2_70), .C2 (n_8_67) );
AOI211_X1 g_12_64 (.ZN (n_12_64), .A (n_11_67), .B (n_5_70), .C1 (n_1_72), .C2 (n_6_68) );
AOI211_X1 g_14_63 (.ZN (n_14_63), .A (n_10_65), .B (n_7_69), .C1 (n_3_71), .C2 (n_4_69) );
AOI211_X1 g_16_62 (.ZN (n_16_62), .A (n_12_64), .B (n_9_68), .C1 (n_5_70), .C2 (n_2_70) );
AOI211_X1 g_15_64 (.ZN (n_15_64), .A (n_14_63), .B (n_11_67), .C1 (n_7_69), .C2 (n_1_72) );
AOI211_X1 g_13_65 (.ZN (n_13_65), .A (n_16_62), .B (n_10_65), .C1 (n_9_68), .C2 (n_3_71) );
AOI211_X1 g_11_66 (.ZN (n_11_66), .A (n_15_64), .B (n_12_64), .C1 (n_11_67), .C2 (n_5_70) );
AOI211_X1 g_9_67 (.ZN (n_9_67), .A (n_13_65), .B (n_14_63), .C1 (n_10_65), .C2 (n_7_69) );
AOI211_X1 g_7_68 (.ZN (n_7_68), .A (n_11_66), .B (n_16_62), .C1 (n_12_64), .C2 (n_9_68) );
AOI211_X1 g_5_69 (.ZN (n_5_69), .A (n_9_67), .B (n_15_64), .C1 (n_14_63), .C2 (n_11_67) );
AOI211_X1 g_4_71 (.ZN (n_4_71), .A (n_7_68), .B (n_13_65), .C1 (n_16_62), .C2 (n_10_65) );
AOI211_X1 g_3_73 (.ZN (n_3_73), .A (n_5_69), .B (n_11_66), .C1 (n_15_64), .C2 (n_12_64) );
AOI211_X1 g_5_74 (.ZN (n_5_74), .A (n_4_71), .B (n_9_67), .C1 (n_13_65), .C2 (n_14_63) );
AOI211_X1 g_3_75 (.ZN (n_3_75), .A (n_3_73), .B (n_7_68), .C1 (n_11_66), .C2 (n_16_62) );
AOI211_X1 g_1_76 (.ZN (n_1_76), .A (n_5_74), .B (n_5_69), .C1 (n_9_67), .C2 (n_15_64) );
AOI211_X1 g_2_74 (.ZN (n_2_74), .A (n_3_75), .B (n_4_71), .C1 (n_7_68), .C2 (n_13_65) );
AOI211_X1 g_4_73 (.ZN (n_4_73), .A (n_1_76), .B (n_3_73), .C1 (n_5_69), .C2 (n_11_66) );
AOI211_X1 g_6_72 (.ZN (n_6_72), .A (n_2_74), .B (n_5_74), .C1 (n_4_71), .C2 (n_9_67) );
AOI211_X1 g_7_70 (.ZN (n_7_70), .A (n_4_73), .B (n_3_75), .C1 (n_3_73), .C2 (n_7_68) );
AOI211_X1 g_8_68 (.ZN (n_8_68), .A (n_6_72), .B (n_1_76), .C1 (n_5_74), .C2 (n_5_69) );
AOI211_X1 g_10_67 (.ZN (n_10_67), .A (n_7_70), .B (n_2_74), .C1 (n_3_75), .C2 (n_4_71) );
AOI211_X1 g_12_66 (.ZN (n_12_66), .A (n_8_68), .B (n_4_73), .C1 (n_1_76), .C2 (n_3_73) );
AOI211_X1 g_14_65 (.ZN (n_14_65), .A (n_10_67), .B (n_6_72), .C1 (n_2_74), .C2 (n_5_74) );
AOI211_X1 g_16_64 (.ZN (n_16_64), .A (n_12_66), .B (n_7_70), .C1 (n_4_73), .C2 (n_3_75) );
AOI211_X1 g_18_63 (.ZN (n_18_63), .A (n_14_65), .B (n_8_68), .C1 (n_6_72), .C2 (n_1_76) );
AOI211_X1 g_20_62 (.ZN (n_20_62), .A (n_16_64), .B (n_10_67), .C1 (n_7_70), .C2 (n_2_74) );
AOI211_X1 g_19_64 (.ZN (n_19_64), .A (n_18_63), .B (n_12_66), .C1 (n_8_68), .C2 (n_4_73) );
AOI211_X1 g_21_63 (.ZN (n_21_63), .A (n_20_62), .B (n_14_65), .C1 (n_10_67), .C2 (n_6_72) );
AOI211_X1 g_23_62 (.ZN (n_23_62), .A (n_19_64), .B (n_16_64), .C1 (n_12_66), .C2 (n_7_70) );
AOI211_X1 g_25_61 (.ZN (n_25_61), .A (n_21_63), .B (n_18_63), .C1 (n_14_65), .C2 (n_8_68) );
AOI211_X1 g_27_60 (.ZN (n_27_60), .A (n_23_62), .B (n_20_62), .C1 (n_16_64), .C2 (n_10_67) );
AOI211_X1 g_29_59 (.ZN (n_29_59), .A (n_25_61), .B (n_19_64), .C1 (n_18_63), .C2 (n_12_66) );
AOI211_X1 g_28_61 (.ZN (n_28_61), .A (n_27_60), .B (n_21_63), .C1 (n_20_62), .C2 (n_14_65) );
AOI211_X1 g_27_59 (.ZN (n_27_59), .A (n_29_59), .B (n_23_62), .C1 (n_19_64), .C2 (n_16_64) );
AOI211_X1 g_29_58 (.ZN (n_29_58), .A (n_28_61), .B (n_25_61), .C1 (n_21_63), .C2 (n_18_63) );
AOI211_X1 g_30_60 (.ZN (n_30_60), .A (n_27_59), .B (n_27_60), .C1 (n_23_62), .C2 (n_20_62) );
AOI211_X1 g_32_59 (.ZN (n_32_59), .A (n_29_58), .B (n_29_59), .C1 (n_25_61), .C2 (n_19_64) );
AOI211_X1 g_34_58 (.ZN (n_34_58), .A (n_30_60), .B (n_28_61), .C1 (n_27_60), .C2 (n_21_63) );
AOI211_X1 g_36_57 (.ZN (n_36_57), .A (n_32_59), .B (n_27_59), .C1 (n_29_59), .C2 (n_23_62) );
AOI211_X1 g_38_56 (.ZN (n_38_56), .A (n_34_58), .B (n_29_58), .C1 (n_28_61), .C2 (n_25_61) );
AOI211_X1 g_40_55 (.ZN (n_40_55), .A (n_36_57), .B (n_30_60), .C1 (n_27_59), .C2 (n_27_60) );
AOI211_X1 g_42_54 (.ZN (n_42_54), .A (n_38_56), .B (n_32_59), .C1 (n_29_58), .C2 (n_29_59) );
AOI211_X1 g_44_53 (.ZN (n_44_53), .A (n_40_55), .B (n_34_58), .C1 (n_30_60), .C2 (n_28_61) );
AOI211_X1 g_46_52 (.ZN (n_46_52), .A (n_42_54), .B (n_36_57), .C1 (n_32_59), .C2 (n_27_59) );
AOI211_X1 g_48_51 (.ZN (n_48_51), .A (n_44_53), .B (n_38_56), .C1 (n_34_58), .C2 (n_29_58) );
AOI211_X1 g_50_50 (.ZN (n_50_50), .A (n_46_52), .B (n_40_55), .C1 (n_36_57), .C2 (n_30_60) );
AOI211_X1 g_52_49 (.ZN (n_52_49), .A (n_48_51), .B (n_42_54), .C1 (n_38_56), .C2 (n_32_59) );
AOI211_X1 g_54_48 (.ZN (n_54_48), .A (n_50_50), .B (n_44_53), .C1 (n_40_55), .C2 (n_34_58) );
AOI211_X1 g_56_47 (.ZN (n_56_47), .A (n_52_49), .B (n_46_52), .C1 (n_42_54), .C2 (n_36_57) );
AOI211_X1 g_58_46 (.ZN (n_58_46), .A (n_54_48), .B (n_48_51), .C1 (n_44_53), .C2 (n_38_56) );
AOI211_X1 g_60_45 (.ZN (n_60_45), .A (n_56_47), .B (n_50_50), .C1 (n_46_52), .C2 (n_40_55) );
AOI211_X1 g_62_44 (.ZN (n_62_44), .A (n_58_46), .B (n_52_49), .C1 (n_48_51), .C2 (n_42_54) );
AOI211_X1 g_64_43 (.ZN (n_64_43), .A (n_60_45), .B (n_54_48), .C1 (n_50_50), .C2 (n_44_53) );
AOI211_X1 g_65_41 (.ZN (n_65_41), .A (n_62_44), .B (n_56_47), .C1 (n_52_49), .C2 (n_46_52) );
AOI211_X1 g_67_40 (.ZN (n_67_40), .A (n_64_43), .B (n_58_46), .C1 (n_54_48), .C2 (n_48_51) );
AOI211_X1 g_69_39 (.ZN (n_69_39), .A (n_65_41), .B (n_60_45), .C1 (n_56_47), .C2 (n_50_50) );
AOI211_X1 g_71_38 (.ZN (n_71_38), .A (n_67_40), .B (n_62_44), .C1 (n_58_46), .C2 (n_52_49) );
AOI211_X1 g_73_37 (.ZN (n_73_37), .A (n_69_39), .B (n_64_43), .C1 (n_60_45), .C2 (n_54_48) );
AOI211_X1 g_75_36 (.ZN (n_75_36), .A (n_71_38), .B (n_65_41), .C1 (n_62_44), .C2 (n_56_47) );
AOI211_X1 g_77_35 (.ZN (n_77_35), .A (n_73_37), .B (n_67_40), .C1 (n_64_43), .C2 (n_58_46) );
AOI211_X1 g_79_34 (.ZN (n_79_34), .A (n_75_36), .B (n_69_39), .C1 (n_65_41), .C2 (n_60_45) );
AOI211_X1 g_81_33 (.ZN (n_81_33), .A (n_77_35), .B (n_71_38), .C1 (n_67_40), .C2 (n_62_44) );
AOI211_X1 g_80_35 (.ZN (n_80_35), .A (n_79_34), .B (n_73_37), .C1 (n_69_39), .C2 (n_64_43) );
AOI211_X1 g_78_34 (.ZN (n_78_34), .A (n_81_33), .B (n_75_36), .C1 (n_71_38), .C2 (n_65_41) );
AOI211_X1 g_76_35 (.ZN (n_76_35), .A (n_80_35), .B (n_77_35), .C1 (n_73_37), .C2 (n_67_40) );
AOI211_X1 g_78_36 (.ZN (n_78_36), .A (n_78_34), .B (n_79_34), .C1 (n_75_36), .C2 (n_69_39) );
AOI211_X1 g_76_37 (.ZN (n_76_37), .A (n_76_35), .B (n_81_33), .C1 (n_77_35), .C2 (n_71_38) );
AOI211_X1 g_74_38 (.ZN (n_74_38), .A (n_78_36), .B (n_80_35), .C1 (n_79_34), .C2 (n_73_37) );
AOI211_X1 g_72_39 (.ZN (n_72_39), .A (n_76_37), .B (n_78_34), .C1 (n_81_33), .C2 (n_75_36) );
AOI211_X1 g_70_40 (.ZN (n_70_40), .A (n_74_38), .B (n_76_35), .C1 (n_80_35), .C2 (n_77_35) );
AOI211_X1 g_68_41 (.ZN (n_68_41), .A (n_72_39), .B (n_78_36), .C1 (n_78_34), .C2 (n_79_34) );
AOI211_X1 g_66_42 (.ZN (n_66_42), .A (n_70_40), .B (n_76_37), .C1 (n_76_35), .C2 (n_81_33) );
AOI211_X1 g_65_44 (.ZN (n_65_44), .A (n_68_41), .B (n_74_38), .C1 (n_78_36), .C2 (n_80_35) );
AOI211_X1 g_64_42 (.ZN (n_64_42), .A (n_66_42), .B (n_72_39), .C1 (n_76_37), .C2 (n_78_34) );
AOI211_X1 g_62_43 (.ZN (n_62_43), .A (n_65_44), .B (n_70_40), .C1 (n_74_38), .C2 (n_76_35) );
AOI211_X1 g_61_45 (.ZN (n_61_45), .A (n_64_42), .B (n_68_41), .C1 (n_72_39), .C2 (n_78_36) );
AOI211_X1 g_63_44 (.ZN (n_63_44), .A (n_62_43), .B (n_66_42), .C1 (n_70_40), .C2 (n_76_37) );
AOI211_X1 g_65_43 (.ZN (n_65_43), .A (n_61_45), .B (n_65_44), .C1 (n_68_41), .C2 (n_74_38) );
AOI211_X1 g_66_41 (.ZN (n_66_41), .A (n_63_44), .B (n_64_42), .C1 (n_66_42), .C2 (n_72_39) );
AOI211_X1 g_68_40 (.ZN (n_68_40), .A (n_65_43), .B (n_62_43), .C1 (n_65_44), .C2 (n_70_40) );
AOI211_X1 g_70_39 (.ZN (n_70_39), .A (n_66_41), .B (n_61_45), .C1 (n_64_42), .C2 (n_68_41) );
AOI211_X1 g_72_38 (.ZN (n_72_38), .A (n_68_40), .B (n_63_44), .C1 (n_62_43), .C2 (n_66_42) );
AOI211_X1 g_74_37 (.ZN (n_74_37), .A (n_70_39), .B (n_65_43), .C1 (n_61_45), .C2 (n_65_44) );
AOI211_X1 g_76_36 (.ZN (n_76_36), .A (n_72_38), .B (n_66_41), .C1 (n_63_44), .C2 (n_64_42) );
AOI211_X1 g_75_38 (.ZN (n_75_38), .A (n_74_37), .B (n_68_40), .C1 (n_65_43), .C2 (n_62_43) );
AOI211_X1 g_77_37 (.ZN (n_77_37), .A (n_76_36), .B (n_70_39), .C1 (n_66_41), .C2 (n_61_45) );
AOI211_X1 g_79_36 (.ZN (n_79_36), .A (n_75_38), .B (n_72_38), .C1 (n_68_40), .C2 (n_63_44) );
AOI211_X1 g_81_35 (.ZN (n_81_35), .A (n_77_37), .B (n_74_37), .C1 (n_70_39), .C2 (n_65_43) );
AOI211_X1 g_80_33 (.ZN (n_80_33), .A (n_79_36), .B (n_76_36), .C1 (n_72_38), .C2 (n_66_41) );
AOI211_X1 g_82_32 (.ZN (n_82_32), .A (n_81_35), .B (n_75_38), .C1 (n_74_37), .C2 (n_68_40) );
AOI211_X1 g_84_31 (.ZN (n_84_31), .A (n_80_33), .B (n_77_37), .C1 (n_76_36), .C2 (n_70_39) );
AOI211_X1 g_86_30 (.ZN (n_86_30), .A (n_82_32), .B (n_79_36), .C1 (n_75_38), .C2 (n_72_38) );
AOI211_X1 g_88_29 (.ZN (n_88_29), .A (n_84_31), .B (n_81_35), .C1 (n_77_37), .C2 (n_74_37) );
AOI211_X1 g_90_28 (.ZN (n_90_28), .A (n_86_30), .B (n_80_33), .C1 (n_79_36), .C2 (n_76_36) );
AOI211_X1 g_92_27 (.ZN (n_92_27), .A (n_88_29), .B (n_82_32), .C1 (n_81_35), .C2 (n_75_38) );
AOI211_X1 g_94_26 (.ZN (n_94_26), .A (n_90_28), .B (n_84_31), .C1 (n_80_33), .C2 (n_77_37) );
AOI211_X1 g_93_28 (.ZN (n_93_28), .A (n_92_27), .B (n_86_30), .C1 (n_82_32), .C2 (n_79_36) );
AOI211_X1 g_91_29 (.ZN (n_91_29), .A (n_94_26), .B (n_88_29), .C1 (n_84_31), .C2 (n_81_35) );
AOI211_X1 g_89_30 (.ZN (n_89_30), .A (n_93_28), .B (n_90_28), .C1 (n_86_30), .C2 (n_80_33) );
AOI211_X1 g_87_31 (.ZN (n_87_31), .A (n_91_29), .B (n_92_27), .C1 (n_88_29), .C2 (n_82_32) );
AOI211_X1 g_85_32 (.ZN (n_85_32), .A (n_89_30), .B (n_94_26), .C1 (n_90_28), .C2 (n_84_31) );
AOI211_X1 g_83_33 (.ZN (n_83_33), .A (n_87_31), .B (n_93_28), .C1 (n_92_27), .C2 (n_86_30) );
AOI211_X1 g_81_34 (.ZN (n_81_34), .A (n_85_32), .B (n_91_29), .C1 (n_94_26), .C2 (n_88_29) );
AOI211_X1 g_79_35 (.ZN (n_79_35), .A (n_83_33), .B (n_89_30), .C1 (n_93_28), .C2 (n_90_28) );
AOI211_X1 g_77_36 (.ZN (n_77_36), .A (n_81_34), .B (n_87_31), .C1 (n_91_29), .C2 (n_92_27) );
AOI211_X1 g_75_37 (.ZN (n_75_37), .A (n_79_35), .B (n_85_32), .C1 (n_89_30), .C2 (n_94_26) );
AOI211_X1 g_73_38 (.ZN (n_73_38), .A (n_77_36), .B (n_83_33), .C1 (n_87_31), .C2 (n_93_28) );
AOI211_X1 g_71_39 (.ZN (n_71_39), .A (n_75_37), .B (n_81_34), .C1 (n_85_32), .C2 (n_91_29) );
AOI211_X1 g_69_40 (.ZN (n_69_40), .A (n_73_38), .B (n_79_35), .C1 (n_83_33), .C2 (n_89_30) );
AOI211_X1 g_67_41 (.ZN (n_67_41), .A (n_71_39), .B (n_77_36), .C1 (n_81_34), .C2 (n_87_31) );
AOI211_X1 g_65_42 (.ZN (n_65_42), .A (n_69_40), .B (n_75_37), .C1 (n_79_35), .C2 (n_85_32) );
AOI211_X1 g_63_43 (.ZN (n_63_43), .A (n_67_41), .B (n_73_38), .C1 (n_77_36), .C2 (n_83_33) );
AOI211_X1 g_61_44 (.ZN (n_61_44), .A (n_65_42), .B (n_71_39), .C1 (n_75_37), .C2 (n_81_34) );
AOI211_X1 g_59_45 (.ZN (n_59_45), .A (n_63_43), .B (n_69_40), .C1 (n_73_38), .C2 (n_79_35) );
AOI211_X1 g_57_46 (.ZN (n_57_46), .A (n_61_44), .B (n_67_41), .C1 (n_71_39), .C2 (n_77_36) );
AOI211_X1 g_55_47 (.ZN (n_55_47), .A (n_59_45), .B (n_65_42), .C1 (n_69_40), .C2 (n_75_37) );
AOI211_X1 g_53_48 (.ZN (n_53_48), .A (n_57_46), .B (n_63_43), .C1 (n_67_41), .C2 (n_73_38) );
AOI211_X1 g_51_49 (.ZN (n_51_49), .A (n_55_47), .B (n_61_44), .C1 (n_65_42), .C2 (n_71_39) );
AOI211_X1 g_49_50 (.ZN (n_49_50), .A (n_53_48), .B (n_59_45), .C1 (n_63_43), .C2 (n_69_40) );
AOI211_X1 g_47_51 (.ZN (n_47_51), .A (n_51_49), .B (n_57_46), .C1 (n_61_44), .C2 (n_67_41) );
AOI211_X1 g_45_52 (.ZN (n_45_52), .A (n_49_50), .B (n_55_47), .C1 (n_59_45), .C2 (n_65_42) );
AOI211_X1 g_43_53 (.ZN (n_43_53), .A (n_47_51), .B (n_53_48), .C1 (n_57_46), .C2 (n_63_43) );
AOI211_X1 g_41_54 (.ZN (n_41_54), .A (n_45_52), .B (n_51_49), .C1 (n_55_47), .C2 (n_61_44) );
AOI211_X1 g_39_55 (.ZN (n_39_55), .A (n_43_53), .B (n_49_50), .C1 (n_53_48), .C2 (n_59_45) );
AOI211_X1 g_37_56 (.ZN (n_37_56), .A (n_41_54), .B (n_47_51), .C1 (n_51_49), .C2 (n_57_46) );
AOI211_X1 g_35_57 (.ZN (n_35_57), .A (n_39_55), .B (n_45_52), .C1 (n_49_50), .C2 (n_55_47) );
AOI211_X1 g_33_58 (.ZN (n_33_58), .A (n_37_56), .B (n_43_53), .C1 (n_47_51), .C2 (n_53_48) );
AOI211_X1 g_31_59 (.ZN (n_31_59), .A (n_35_57), .B (n_41_54), .C1 (n_45_52), .C2 (n_51_49) );
AOI211_X1 g_29_60 (.ZN (n_29_60), .A (n_33_58), .B (n_39_55), .C1 (n_43_53), .C2 (n_49_50) );
AOI211_X1 g_27_61 (.ZN (n_27_61), .A (n_31_59), .B (n_37_56), .C1 (n_41_54), .C2 (n_47_51) );
AOI211_X1 g_25_60 (.ZN (n_25_60), .A (n_29_60), .B (n_35_57), .C1 (n_39_55), .C2 (n_45_52) );
AOI211_X1 g_23_61 (.ZN (n_23_61), .A (n_27_61), .B (n_33_58), .C1 (n_37_56), .C2 (n_43_53) );
AOI211_X1 g_21_62 (.ZN (n_21_62), .A (n_25_60), .B (n_31_59), .C1 (n_35_57), .C2 (n_41_54) );
AOI211_X1 g_20_64 (.ZN (n_20_64), .A (n_23_61), .B (n_29_60), .C1 (n_33_58), .C2 (n_39_55) );
AOI211_X1 g_22_63 (.ZN (n_22_63), .A (n_21_62), .B (n_27_61), .C1 (n_31_59), .C2 (n_37_56) );
AOI211_X1 g_24_62 (.ZN (n_24_62), .A (n_20_64), .B (n_25_60), .C1 (n_29_60), .C2 (n_35_57) );
AOI211_X1 g_26_61 (.ZN (n_26_61), .A (n_22_63), .B (n_23_61), .C1 (n_27_61), .C2 (n_33_58) );
AOI211_X1 g_28_60 (.ZN (n_28_60), .A (n_24_62), .B (n_21_62), .C1 (n_25_60), .C2 (n_31_59) );
AOI211_X1 g_30_59 (.ZN (n_30_59), .A (n_26_61), .B (n_20_64), .C1 (n_23_61), .C2 (n_29_60) );
AOI211_X1 g_32_58 (.ZN (n_32_58), .A (n_28_60), .B (n_22_63), .C1 (n_21_62), .C2 (n_27_61) );
AOI211_X1 g_34_57 (.ZN (n_34_57), .A (n_30_59), .B (n_24_62), .C1 (n_20_64), .C2 (n_25_60) );
AOI211_X1 g_36_56 (.ZN (n_36_56), .A (n_32_58), .B (n_26_61), .C1 (n_22_63), .C2 (n_23_61) );
AOI211_X1 g_38_55 (.ZN (n_38_55), .A (n_34_57), .B (n_28_60), .C1 (n_24_62), .C2 (n_21_62) );
AOI211_X1 g_40_54 (.ZN (n_40_54), .A (n_36_56), .B (n_30_59), .C1 (n_26_61), .C2 (n_20_64) );
AOI211_X1 g_42_53 (.ZN (n_42_53), .A (n_38_55), .B (n_32_58), .C1 (n_28_60), .C2 (n_22_63) );
AOI211_X1 g_41_55 (.ZN (n_41_55), .A (n_40_54), .B (n_34_57), .C1 (n_30_59), .C2 (n_24_62) );
AOI211_X1 g_43_54 (.ZN (n_43_54), .A (n_42_53), .B (n_36_56), .C1 (n_32_58), .C2 (n_26_61) );
AOI211_X1 g_45_53 (.ZN (n_45_53), .A (n_41_55), .B (n_38_55), .C1 (n_34_57), .C2 (n_28_60) );
AOI211_X1 g_47_52 (.ZN (n_47_52), .A (n_43_54), .B (n_40_54), .C1 (n_36_56), .C2 (n_30_59) );
AOI211_X1 g_49_51 (.ZN (n_49_51), .A (n_45_53), .B (n_42_53), .C1 (n_38_55), .C2 (n_32_58) );
AOI211_X1 g_51_50 (.ZN (n_51_50), .A (n_47_52), .B (n_41_55), .C1 (n_40_54), .C2 (n_34_57) );
AOI211_X1 g_53_49 (.ZN (n_53_49), .A (n_49_51), .B (n_43_54), .C1 (n_42_53), .C2 (n_36_56) );
AOI211_X1 g_55_48 (.ZN (n_55_48), .A (n_51_50), .B (n_45_53), .C1 (n_41_55), .C2 (n_38_55) );
AOI211_X1 g_57_47 (.ZN (n_57_47), .A (n_53_49), .B (n_47_52), .C1 (n_43_54), .C2 (n_40_54) );
AOI211_X1 g_59_46 (.ZN (n_59_46), .A (n_55_48), .B (n_49_51), .C1 (n_45_53), .C2 (n_42_53) );
AOI211_X1 g_58_48 (.ZN (n_58_48), .A (n_57_47), .B (n_51_50), .C1 (n_47_52), .C2 (n_41_55) );
AOI211_X1 g_60_47 (.ZN (n_60_47), .A (n_59_46), .B (n_53_49), .C1 (n_49_51), .C2 (n_43_54) );
AOI211_X1 g_62_46 (.ZN (n_62_46), .A (n_58_48), .B (n_55_48), .C1 (n_51_50), .C2 (n_45_53) );
AOI211_X1 g_64_45 (.ZN (n_64_45), .A (n_60_47), .B (n_57_47), .C1 (n_53_49), .C2 (n_47_52) );
AOI211_X1 g_66_44 (.ZN (n_66_44), .A (n_62_46), .B (n_59_46), .C1 (n_55_48), .C2 (n_49_51) );
AOI211_X1 g_67_42 (.ZN (n_67_42), .A (n_64_45), .B (n_58_48), .C1 (n_57_47), .C2 (n_51_50) );
AOI211_X1 g_69_41 (.ZN (n_69_41), .A (n_66_44), .B (n_60_47), .C1 (n_59_46), .C2 (n_53_49) );
AOI211_X1 g_71_40 (.ZN (n_71_40), .A (n_67_42), .B (n_62_46), .C1 (n_58_48), .C2 (n_55_48) );
AOI211_X1 g_73_39 (.ZN (n_73_39), .A (n_69_41), .B (n_64_45), .C1 (n_60_47), .C2 (n_57_47) );
AOI211_X1 g_72_41 (.ZN (n_72_41), .A (n_71_40), .B (n_66_44), .C1 (n_62_46), .C2 (n_59_46) );
AOI211_X1 g_74_40 (.ZN (n_74_40), .A (n_73_39), .B (n_67_42), .C1 (n_64_45), .C2 (n_58_48) );
AOI211_X1 g_76_39 (.ZN (n_76_39), .A (n_72_41), .B (n_69_41), .C1 (n_66_44), .C2 (n_60_47) );
AOI211_X1 g_78_38 (.ZN (n_78_38), .A (n_74_40), .B (n_71_40), .C1 (n_67_42), .C2 (n_62_46) );
AOI211_X1 g_80_37 (.ZN (n_80_37), .A (n_76_39), .B (n_73_39), .C1 (n_69_41), .C2 (n_64_45) );
AOI211_X1 g_82_36 (.ZN (n_82_36), .A (n_78_38), .B (n_72_41), .C1 (n_71_40), .C2 (n_66_44) );
AOI211_X1 g_83_34 (.ZN (n_83_34), .A (n_80_37), .B (n_74_40), .C1 (n_73_39), .C2 (n_67_42) );
AOI211_X1 g_85_33 (.ZN (n_85_33), .A (n_82_36), .B (n_76_39), .C1 (n_72_41), .C2 (n_69_41) );
AOI211_X1 g_87_32 (.ZN (n_87_32), .A (n_83_34), .B (n_78_38), .C1 (n_74_40), .C2 (n_71_40) );
AOI211_X1 g_85_31 (.ZN (n_85_31), .A (n_85_33), .B (n_80_37), .C1 (n_76_39), .C2 (n_73_39) );
AOI211_X1 g_87_30 (.ZN (n_87_30), .A (n_87_32), .B (n_82_36), .C1 (n_78_38), .C2 (n_72_41) );
AOI211_X1 g_89_29 (.ZN (n_89_29), .A (n_85_31), .B (n_83_34), .C1 (n_80_37), .C2 (n_74_40) );
AOI211_X1 g_91_28 (.ZN (n_91_28), .A (n_87_30), .B (n_85_33), .C1 (n_82_36), .C2 (n_76_39) );
AOI211_X1 g_93_27 (.ZN (n_93_27), .A (n_89_29), .B (n_87_32), .C1 (n_83_34), .C2 (n_78_38) );
AOI211_X1 g_95_26 (.ZN (n_95_26), .A (n_91_28), .B (n_85_31), .C1 (n_85_33), .C2 (n_80_37) );
AOI211_X1 g_97_25 (.ZN (n_97_25), .A (n_93_27), .B (n_87_30), .C1 (n_87_32), .C2 (n_82_36) );
AOI211_X1 g_99_24 (.ZN (n_99_24), .A (n_95_26), .B (n_89_29), .C1 (n_85_31), .C2 (n_83_34) );
AOI211_X1 g_98_26 (.ZN (n_98_26), .A (n_97_25), .B (n_91_28), .C1 (n_87_30), .C2 (n_85_33) );
AOI211_X1 g_100_25 (.ZN (n_100_25), .A (n_99_24), .B (n_93_27), .C1 (n_89_29), .C2 (n_87_32) );
AOI211_X1 g_102_24 (.ZN (n_102_24), .A (n_98_26), .B (n_95_26), .C1 (n_91_28), .C2 (n_85_31) );
AOI211_X1 g_101_26 (.ZN (n_101_26), .A (n_100_25), .B (n_97_25), .C1 (n_93_27), .C2 (n_87_30) );
AOI211_X1 g_100_24 (.ZN (n_100_24), .A (n_102_24), .B (n_99_24), .C1 (n_95_26), .C2 (n_89_29) );
AOI211_X1 g_98_25 (.ZN (n_98_25), .A (n_101_26), .B (n_98_26), .C1 (n_97_25), .C2 (n_91_28) );
AOI211_X1 g_99_27 (.ZN (n_99_27), .A (n_100_24), .B (n_100_25), .C1 (n_99_24), .C2 (n_93_27) );
AOI211_X1 g_97_28 (.ZN (n_97_28), .A (n_98_25), .B (n_102_24), .C1 (n_98_26), .C2 (n_95_26) );
AOI211_X1 g_95_29 (.ZN (n_95_29), .A (n_99_27), .B (n_101_26), .C1 (n_100_25), .C2 (n_97_25) );
AOI211_X1 g_96_27 (.ZN (n_96_27), .A (n_97_28), .B (n_100_24), .C1 (n_102_24), .C2 (n_99_24) );
AOI211_X1 g_94_28 (.ZN (n_94_28), .A (n_95_29), .B (n_98_25), .C1 (n_101_26), .C2 (n_98_26) );
AOI211_X1 g_92_29 (.ZN (n_92_29), .A (n_96_27), .B (n_99_27), .C1 (n_100_24), .C2 (n_100_25) );
AOI211_X1 g_90_30 (.ZN (n_90_30), .A (n_94_28), .B (n_97_28), .C1 (n_98_25), .C2 (n_102_24) );
AOI211_X1 g_88_31 (.ZN (n_88_31), .A (n_92_29), .B (n_95_29), .C1 (n_99_27), .C2 (n_101_26) );
AOI211_X1 g_86_32 (.ZN (n_86_32), .A (n_90_30), .B (n_96_27), .C1 (n_97_28), .C2 (n_100_24) );
AOI211_X1 g_84_33 (.ZN (n_84_33), .A (n_88_31), .B (n_94_28), .C1 (n_95_29), .C2 (n_98_25) );
AOI211_X1 g_82_34 (.ZN (n_82_34), .A (n_86_32), .B (n_92_29), .C1 (n_96_27), .C2 (n_99_27) );
AOI211_X1 g_84_35 (.ZN (n_84_35), .A (n_84_33), .B (n_90_30), .C1 (n_94_28), .C2 (n_97_28) );
AOI211_X1 g_86_34 (.ZN (n_86_34), .A (n_82_34), .B (n_88_31), .C1 (n_92_29), .C2 (n_95_29) );
AOI211_X1 g_88_33 (.ZN (n_88_33), .A (n_84_35), .B (n_86_32), .C1 (n_90_30), .C2 (n_96_27) );
AOI211_X1 g_89_31 (.ZN (n_89_31), .A (n_86_34), .B (n_84_33), .C1 (n_88_31), .C2 (n_94_28) );
AOI211_X1 g_91_30 (.ZN (n_91_30), .A (n_88_33), .B (n_82_34), .C1 (n_86_32), .C2 (n_92_29) );
AOI211_X1 g_93_29 (.ZN (n_93_29), .A (n_89_31), .B (n_84_35), .C1 (n_84_33), .C2 (n_90_30) );
AOI211_X1 g_95_28 (.ZN (n_95_28), .A (n_91_30), .B (n_86_34), .C1 (n_82_34), .C2 (n_88_31) );
AOI211_X1 g_97_27 (.ZN (n_97_27), .A (n_93_29), .B (n_88_33), .C1 (n_84_35), .C2 (n_86_32) );
AOI211_X1 g_99_26 (.ZN (n_99_26), .A (n_95_28), .B (n_89_31), .C1 (n_86_34), .C2 (n_84_33) );
AOI211_X1 g_101_25 (.ZN (n_101_25), .A (n_97_27), .B (n_91_30), .C1 (n_88_33), .C2 (n_82_34) );
AOI211_X1 g_102_23 (.ZN (n_102_23), .A (n_99_26), .B (n_93_29), .C1 (n_89_31), .C2 (n_84_35) );
AOI211_X1 g_104_22 (.ZN (n_104_22), .A (n_101_25), .B (n_95_28), .C1 (n_91_30), .C2 (n_86_34) );
AOI211_X1 g_106_21 (.ZN (n_106_21), .A (n_102_23), .B (n_97_27), .C1 (n_93_29), .C2 (n_88_33) );
AOI211_X1 g_108_20 (.ZN (n_108_20), .A (n_104_22), .B (n_99_26), .C1 (n_95_28), .C2 (n_89_31) );
AOI211_X1 g_110_19 (.ZN (n_110_19), .A (n_106_21), .B (n_101_25), .C1 (n_97_27), .C2 (n_91_30) );
AOI211_X1 g_112_18 (.ZN (n_112_18), .A (n_108_20), .B (n_102_23), .C1 (n_99_26), .C2 (n_93_29) );
AOI211_X1 g_114_17 (.ZN (n_114_17), .A (n_110_19), .B (n_104_22), .C1 (n_101_25), .C2 (n_95_28) );
AOI211_X1 g_116_16 (.ZN (n_116_16), .A (n_112_18), .B (n_106_21), .C1 (n_102_23), .C2 (n_97_27) );
AOI211_X1 g_118_17 (.ZN (n_118_17), .A (n_114_17), .B (n_108_20), .C1 (n_104_22), .C2 (n_99_26) );
AOI211_X1 g_116_18 (.ZN (n_116_18), .A (n_116_16), .B (n_110_19), .C1 (n_106_21), .C2 (n_101_25) );
AOI211_X1 g_114_19 (.ZN (n_114_19), .A (n_118_17), .B (n_112_18), .C1 (n_108_20), .C2 (n_102_23) );
AOI211_X1 g_112_20 (.ZN (n_112_20), .A (n_116_18), .B (n_114_17), .C1 (n_110_19), .C2 (n_104_22) );
AOI211_X1 g_110_21 (.ZN (n_110_21), .A (n_114_19), .B (n_116_16), .C1 (n_112_18), .C2 (n_106_21) );
AOI211_X1 g_108_22 (.ZN (n_108_22), .A (n_112_20), .B (n_118_17), .C1 (n_114_17), .C2 (n_108_20) );
AOI211_X1 g_106_23 (.ZN (n_106_23), .A (n_110_21), .B (n_116_18), .C1 (n_116_16), .C2 (n_110_19) );
AOI211_X1 g_104_24 (.ZN (n_104_24), .A (n_108_22), .B (n_114_19), .C1 (n_118_17), .C2 (n_112_18) );
AOI211_X1 g_102_25 (.ZN (n_102_25), .A (n_106_23), .B (n_112_20), .C1 (n_116_18), .C2 (n_114_17) );
AOI211_X1 g_100_26 (.ZN (n_100_26), .A (n_104_24), .B (n_110_21), .C1 (n_114_19), .C2 (n_116_16) );
AOI211_X1 g_98_27 (.ZN (n_98_27), .A (n_102_25), .B (n_108_22), .C1 (n_112_20), .C2 (n_118_17) );
AOI211_X1 g_96_28 (.ZN (n_96_28), .A (n_100_26), .B (n_106_23), .C1 (n_110_21), .C2 (n_116_18) );
AOI211_X1 g_94_29 (.ZN (n_94_29), .A (n_98_27), .B (n_104_24), .C1 (n_108_22), .C2 (n_114_19) );
AOI211_X1 g_92_30 (.ZN (n_92_30), .A (n_96_28), .B (n_102_25), .C1 (n_106_23), .C2 (n_112_20) );
AOI211_X1 g_90_31 (.ZN (n_90_31), .A (n_94_29), .B (n_100_26), .C1 (n_104_24), .C2 (n_110_21) );
AOI211_X1 g_88_32 (.ZN (n_88_32), .A (n_92_30), .B (n_98_27), .C1 (n_102_25), .C2 (n_108_22) );
AOI211_X1 g_86_33 (.ZN (n_86_33), .A (n_90_31), .B (n_96_28), .C1 (n_100_26), .C2 (n_106_23) );
AOI211_X1 g_84_34 (.ZN (n_84_34), .A (n_88_32), .B (n_94_29), .C1 (n_98_27), .C2 (n_104_24) );
AOI211_X1 g_82_35 (.ZN (n_82_35), .A (n_86_33), .B (n_92_30), .C1 (n_96_28), .C2 (n_102_25) );
AOI211_X1 g_80_36 (.ZN (n_80_36), .A (n_84_34), .B (n_90_31), .C1 (n_94_29), .C2 (n_100_26) );
AOI211_X1 g_78_37 (.ZN (n_78_37), .A (n_82_35), .B (n_88_32), .C1 (n_92_30), .C2 (n_98_27) );
AOI211_X1 g_76_38 (.ZN (n_76_38), .A (n_80_36), .B (n_86_33), .C1 (n_90_31), .C2 (n_96_28) );
AOI211_X1 g_74_39 (.ZN (n_74_39), .A (n_78_37), .B (n_84_34), .C1 (n_88_32), .C2 (n_94_29) );
AOI211_X1 g_72_40 (.ZN (n_72_40), .A (n_76_38), .B (n_82_35), .C1 (n_86_33), .C2 (n_92_30) );
AOI211_X1 g_70_41 (.ZN (n_70_41), .A (n_74_39), .B (n_80_36), .C1 (n_84_34), .C2 (n_90_31) );
AOI211_X1 g_68_42 (.ZN (n_68_42), .A (n_72_40), .B (n_78_37), .C1 (n_82_35), .C2 (n_88_32) );
AOI211_X1 g_66_43 (.ZN (n_66_43), .A (n_70_41), .B (n_76_38), .C1 (n_80_36), .C2 (n_86_33) );
AOI211_X1 g_64_44 (.ZN (n_64_44), .A (n_68_42), .B (n_74_39), .C1 (n_78_37), .C2 (n_84_34) );
AOI211_X1 g_62_45 (.ZN (n_62_45), .A (n_66_43), .B (n_72_40), .C1 (n_76_38), .C2 (n_82_35) );
AOI211_X1 g_60_46 (.ZN (n_60_46), .A (n_64_44), .B (n_70_41), .C1 (n_74_39), .C2 (n_80_36) );
AOI211_X1 g_58_47 (.ZN (n_58_47), .A (n_62_45), .B (n_68_42), .C1 (n_72_40), .C2 (n_78_37) );
AOI211_X1 g_56_48 (.ZN (n_56_48), .A (n_60_46), .B (n_66_43), .C1 (n_70_41), .C2 (n_76_38) );
AOI211_X1 g_54_49 (.ZN (n_54_49), .A (n_58_47), .B (n_64_44), .C1 (n_68_42), .C2 (n_74_39) );
AOI211_X1 g_52_50 (.ZN (n_52_50), .A (n_56_48), .B (n_62_45), .C1 (n_66_43), .C2 (n_72_40) );
AOI211_X1 g_50_51 (.ZN (n_50_51), .A (n_54_49), .B (n_60_46), .C1 (n_64_44), .C2 (n_70_41) );
AOI211_X1 g_48_52 (.ZN (n_48_52), .A (n_52_50), .B (n_58_47), .C1 (n_62_45), .C2 (n_68_42) );
AOI211_X1 g_46_53 (.ZN (n_46_53), .A (n_50_51), .B (n_56_48), .C1 (n_60_46), .C2 (n_66_43) );
AOI211_X1 g_44_54 (.ZN (n_44_54), .A (n_48_52), .B (n_54_49), .C1 (n_58_47), .C2 (n_64_44) );
AOI211_X1 g_42_55 (.ZN (n_42_55), .A (n_46_53), .B (n_52_50), .C1 (n_56_48), .C2 (n_62_45) );
AOI211_X1 g_40_56 (.ZN (n_40_56), .A (n_44_54), .B (n_50_51), .C1 (n_54_49), .C2 (n_60_46) );
AOI211_X1 g_38_57 (.ZN (n_38_57), .A (n_42_55), .B (n_48_52), .C1 (n_52_50), .C2 (n_58_47) );
AOI211_X1 g_36_58 (.ZN (n_36_58), .A (n_40_56), .B (n_46_53), .C1 (n_50_51), .C2 (n_56_48) );
AOI211_X1 g_34_59 (.ZN (n_34_59), .A (n_38_57), .B (n_44_54), .C1 (n_48_52), .C2 (n_54_49) );
AOI211_X1 g_32_60 (.ZN (n_32_60), .A (n_36_58), .B (n_42_55), .C1 (n_46_53), .C2 (n_52_50) );
AOI211_X1 g_30_61 (.ZN (n_30_61), .A (n_34_59), .B (n_40_56), .C1 (n_44_54), .C2 (n_50_51) );
AOI211_X1 g_28_62 (.ZN (n_28_62), .A (n_32_60), .B (n_38_57), .C1 (n_42_55), .C2 (n_48_52) );
AOI211_X1 g_26_63 (.ZN (n_26_63), .A (n_30_61), .B (n_36_58), .C1 (n_40_56), .C2 (n_46_53) );
AOI211_X1 g_24_64 (.ZN (n_24_64), .A (n_28_62), .B (n_34_59), .C1 (n_38_57), .C2 (n_44_54) );
AOI211_X1 g_25_62 (.ZN (n_25_62), .A (n_26_63), .B (n_32_60), .C1 (n_36_58), .C2 (n_42_55) );
AOI211_X1 g_23_63 (.ZN (n_23_63), .A (n_24_64), .B (n_30_61), .C1 (n_34_59), .C2 (n_40_56) );
AOI211_X1 g_21_64 (.ZN (n_21_64), .A (n_25_62), .B (n_28_62), .C1 (n_32_60), .C2 (n_38_57) );
AOI211_X1 g_19_65 (.ZN (n_19_65), .A (n_23_63), .B (n_26_63), .C1 (n_30_61), .C2 (n_36_58) );
AOI211_X1 g_17_64 (.ZN (n_17_64), .A (n_21_64), .B (n_24_64), .C1 (n_28_62), .C2 (n_34_59) );
AOI211_X1 g_15_65 (.ZN (n_15_65), .A (n_19_65), .B (n_25_62), .C1 (n_26_63), .C2 (n_32_60) );
AOI211_X1 g_13_66 (.ZN (n_13_66), .A (n_17_64), .B (n_23_63), .C1 (n_24_64), .C2 (n_30_61) );
AOI211_X1 g_12_68 (.ZN (n_12_68), .A (n_15_65), .B (n_21_64), .C1 (n_25_62), .C2 (n_28_62) );
AOI211_X1 g_14_67 (.ZN (n_14_67), .A (n_13_66), .B (n_19_65), .C1 (n_23_63), .C2 (n_26_63) );
AOI211_X1 g_16_66 (.ZN (n_16_66), .A (n_12_68), .B (n_17_64), .C1 (n_21_64), .C2 (n_24_64) );
AOI211_X1 g_18_65 (.ZN (n_18_65), .A (n_14_67), .B (n_15_65), .C1 (n_19_65), .C2 (n_25_62) );
AOI211_X1 g_20_66 (.ZN (n_20_66), .A (n_16_66), .B (n_13_66), .C1 (n_17_64), .C2 (n_23_63) );
AOI211_X1 g_22_65 (.ZN (n_22_65), .A (n_18_65), .B (n_12_68), .C1 (n_15_65), .C2 (n_21_64) );
AOI211_X1 g_21_67 (.ZN (n_21_67), .A (n_20_66), .B (n_14_67), .C1 (n_13_66), .C2 (n_19_65) );
AOI211_X1 g_20_65 (.ZN (n_20_65), .A (n_22_65), .B (n_16_66), .C1 (n_12_68), .C2 (n_17_64) );
AOI211_X1 g_22_64 (.ZN (n_22_64), .A (n_21_67), .B (n_18_65), .C1 (n_14_67), .C2 (n_15_65) );
AOI211_X1 g_24_63 (.ZN (n_24_63), .A (n_20_65), .B (n_20_66), .C1 (n_16_66), .C2 (n_13_66) );
AOI211_X1 g_26_62 (.ZN (n_26_62), .A (n_22_64), .B (n_22_65), .C1 (n_18_65), .C2 (n_12_68) );
AOI211_X1 g_25_64 (.ZN (n_25_64), .A (n_24_63), .B (n_21_67), .C1 (n_20_66), .C2 (n_14_67) );
AOI211_X1 g_27_63 (.ZN (n_27_63), .A (n_26_62), .B (n_20_65), .C1 (n_22_65), .C2 (n_16_66) );
AOI211_X1 g_29_62 (.ZN (n_29_62), .A (n_25_64), .B (n_22_64), .C1 (n_21_67), .C2 (n_18_65) );
AOI211_X1 g_31_61 (.ZN (n_31_61), .A (n_27_63), .B (n_24_63), .C1 (n_20_65), .C2 (n_20_66) );
AOI211_X1 g_33_60 (.ZN (n_33_60), .A (n_29_62), .B (n_26_62), .C1 (n_22_64), .C2 (n_22_65) );
AOI211_X1 g_35_59 (.ZN (n_35_59), .A (n_31_61), .B (n_25_64), .C1 (n_24_63), .C2 (n_21_67) );
AOI211_X1 g_37_58 (.ZN (n_37_58), .A (n_33_60), .B (n_27_63), .C1 (n_26_62), .C2 (n_20_65) );
AOI211_X1 g_39_57 (.ZN (n_39_57), .A (n_35_59), .B (n_29_62), .C1 (n_25_64), .C2 (n_22_64) );
AOI211_X1 g_41_56 (.ZN (n_41_56), .A (n_37_58), .B (n_31_61), .C1 (n_27_63), .C2 (n_24_63) );
AOI211_X1 g_43_55 (.ZN (n_43_55), .A (n_39_57), .B (n_33_60), .C1 (n_29_62), .C2 (n_26_62) );
AOI211_X1 g_45_54 (.ZN (n_45_54), .A (n_41_56), .B (n_35_59), .C1 (n_31_61), .C2 (n_25_64) );
AOI211_X1 g_47_53 (.ZN (n_47_53), .A (n_43_55), .B (n_37_58), .C1 (n_33_60), .C2 (n_27_63) );
AOI211_X1 g_49_52 (.ZN (n_49_52), .A (n_45_54), .B (n_39_57), .C1 (n_35_59), .C2 (n_29_62) );
AOI211_X1 g_51_51 (.ZN (n_51_51), .A (n_47_53), .B (n_41_56), .C1 (n_37_58), .C2 (n_31_61) );
AOI211_X1 g_53_50 (.ZN (n_53_50), .A (n_49_52), .B (n_43_55), .C1 (n_39_57), .C2 (n_33_60) );
AOI211_X1 g_55_49 (.ZN (n_55_49), .A (n_51_51), .B (n_45_54), .C1 (n_41_56), .C2 (n_35_59) );
AOI211_X1 g_57_48 (.ZN (n_57_48), .A (n_53_50), .B (n_47_53), .C1 (n_43_55), .C2 (n_37_58) );
AOI211_X1 g_59_47 (.ZN (n_59_47), .A (n_55_49), .B (n_49_52), .C1 (n_45_54), .C2 (n_39_57) );
AOI211_X1 g_61_46 (.ZN (n_61_46), .A (n_57_48), .B (n_51_51), .C1 (n_47_53), .C2 (n_41_56) );
AOI211_X1 g_63_45 (.ZN (n_63_45), .A (n_59_47), .B (n_53_50), .C1 (n_49_52), .C2 (n_43_55) );
AOI211_X1 g_62_47 (.ZN (n_62_47), .A (n_61_46), .B (n_55_49), .C1 (n_51_51), .C2 (n_45_54) );
AOI211_X1 g_64_46 (.ZN (n_64_46), .A (n_63_45), .B (n_57_48), .C1 (n_53_50), .C2 (n_47_53) );
AOI211_X1 g_66_45 (.ZN (n_66_45), .A (n_62_47), .B (n_59_47), .C1 (n_55_49), .C2 (n_49_52) );
AOI211_X1 g_67_43 (.ZN (n_67_43), .A (n_64_46), .B (n_61_46), .C1 (n_57_48), .C2 (n_51_51) );
AOI211_X1 g_69_42 (.ZN (n_69_42), .A (n_66_45), .B (n_63_45), .C1 (n_59_47), .C2 (n_53_50) );
AOI211_X1 g_71_41 (.ZN (n_71_41), .A (n_67_43), .B (n_62_47), .C1 (n_61_46), .C2 (n_55_49) );
AOI211_X1 g_73_40 (.ZN (n_73_40), .A (n_69_42), .B (n_64_46), .C1 (n_63_45), .C2 (n_57_48) );
AOI211_X1 g_75_39 (.ZN (n_75_39), .A (n_71_41), .B (n_66_45), .C1 (n_62_47), .C2 (n_59_47) );
AOI211_X1 g_77_38 (.ZN (n_77_38), .A (n_73_40), .B (n_67_43), .C1 (n_64_46), .C2 (n_61_46) );
AOI211_X1 g_79_37 (.ZN (n_79_37), .A (n_75_39), .B (n_69_42), .C1 (n_66_45), .C2 (n_63_45) );
AOI211_X1 g_81_36 (.ZN (n_81_36), .A (n_77_38), .B (n_71_41), .C1 (n_67_43), .C2 (n_62_47) );
AOI211_X1 g_83_35 (.ZN (n_83_35), .A (n_79_37), .B (n_73_40), .C1 (n_69_42), .C2 (n_64_46) );
AOI211_X1 g_85_34 (.ZN (n_85_34), .A (n_81_36), .B (n_75_39), .C1 (n_71_41), .C2 (n_66_45) );
AOI211_X1 g_87_33 (.ZN (n_87_33), .A (n_83_35), .B (n_77_38), .C1 (n_73_40), .C2 (n_67_43) );
AOI211_X1 g_89_32 (.ZN (n_89_32), .A (n_85_34), .B (n_79_37), .C1 (n_75_39), .C2 (n_69_42) );
AOI211_X1 g_91_31 (.ZN (n_91_31), .A (n_87_33), .B (n_81_36), .C1 (n_77_38), .C2 (n_71_41) );
AOI211_X1 g_93_30 (.ZN (n_93_30), .A (n_89_32), .B (n_83_35), .C1 (n_79_37), .C2 (n_73_40) );
AOI211_X1 g_92_32 (.ZN (n_92_32), .A (n_91_31), .B (n_85_34), .C1 (n_81_36), .C2 (n_75_39) );
AOI211_X1 g_94_31 (.ZN (n_94_31), .A (n_93_30), .B (n_87_33), .C1 (n_83_35), .C2 (n_77_38) );
AOI211_X1 g_96_30 (.ZN (n_96_30), .A (n_92_32), .B (n_89_32), .C1 (n_85_34), .C2 (n_79_37) );
AOI211_X1 g_98_29 (.ZN (n_98_29), .A (n_94_31), .B (n_91_31), .C1 (n_87_33), .C2 (n_81_36) );
AOI211_X1 g_100_28 (.ZN (n_100_28), .A (n_96_30), .B (n_93_30), .C1 (n_89_32), .C2 (n_83_35) );
AOI211_X1 g_102_27 (.ZN (n_102_27), .A (n_98_29), .B (n_92_32), .C1 (n_91_31), .C2 (n_85_34) );
AOI211_X1 g_103_25 (.ZN (n_103_25), .A (n_100_28), .B (n_94_31), .C1 (n_93_30), .C2 (n_87_33) );
AOI211_X1 g_105_24 (.ZN (n_105_24), .A (n_102_27), .B (n_96_30), .C1 (n_92_32), .C2 (n_89_32) );
AOI211_X1 g_106_22 (.ZN (n_106_22), .A (n_103_25), .B (n_98_29), .C1 (n_94_31), .C2 (n_91_31) );
AOI211_X1 g_108_21 (.ZN (n_108_21), .A (n_105_24), .B (n_100_28), .C1 (n_96_30), .C2 (n_93_30) );
AOI211_X1 g_110_20 (.ZN (n_110_20), .A (n_106_22), .B (n_102_27), .C1 (n_98_29), .C2 (n_92_32) );
AOI211_X1 g_112_19 (.ZN (n_112_19), .A (n_108_21), .B (n_103_25), .C1 (n_100_28), .C2 (n_94_31) );
AOI211_X1 g_114_18 (.ZN (n_114_18), .A (n_110_20), .B (n_105_24), .C1 (n_102_27), .C2 (n_96_30) );
AOI211_X1 g_116_17 (.ZN (n_116_17), .A (n_112_19), .B (n_106_22), .C1 (n_103_25), .C2 (n_98_29) );
AOI211_X1 g_118_16 (.ZN (n_118_16), .A (n_114_18), .B (n_108_21), .C1 (n_105_24), .C2 (n_100_28) );
AOI211_X1 g_120_15 (.ZN (n_120_15), .A (n_116_17), .B (n_110_20), .C1 (n_106_22), .C2 (n_102_27) );
AOI211_X1 g_119_17 (.ZN (n_119_17), .A (n_118_16), .B (n_112_19), .C1 (n_108_21), .C2 (n_103_25) );
AOI211_X1 g_117_18 (.ZN (n_117_18), .A (n_120_15), .B (n_114_18), .C1 (n_110_20), .C2 (n_105_24) );
AOI211_X1 g_115_19 (.ZN (n_115_19), .A (n_119_17), .B (n_116_17), .C1 (n_112_19), .C2 (n_106_22) );
AOI211_X1 g_113_20 (.ZN (n_113_20), .A (n_117_18), .B (n_118_16), .C1 (n_114_18), .C2 (n_108_21) );
AOI211_X1 g_111_21 (.ZN (n_111_21), .A (n_115_19), .B (n_120_15), .C1 (n_116_17), .C2 (n_110_20) );
AOI211_X1 g_109_22 (.ZN (n_109_22), .A (n_113_20), .B (n_119_17), .C1 (n_118_16), .C2 (n_112_19) );
AOI211_X1 g_107_23 (.ZN (n_107_23), .A (n_111_21), .B (n_117_18), .C1 (n_120_15), .C2 (n_114_18) );
AOI211_X1 g_106_25 (.ZN (n_106_25), .A (n_109_22), .B (n_115_19), .C1 (n_119_17), .C2 (n_116_17) );
AOI211_X1 g_105_23 (.ZN (n_105_23), .A (n_107_23), .B (n_113_20), .C1 (n_117_18), .C2 (n_118_16) );
AOI211_X1 g_103_24 (.ZN (n_103_24), .A (n_106_25), .B (n_111_21), .C1 (n_115_19), .C2 (n_120_15) );
AOI211_X1 g_104_26 (.ZN (n_104_26), .A (n_105_23), .B (n_109_22), .C1 (n_113_20), .C2 (n_119_17) );
AOI211_X1 g_103_28 (.ZN (n_103_28), .A (n_103_24), .B (n_107_23), .C1 (n_111_21), .C2 (n_117_18) );
AOI211_X1 g_102_26 (.ZN (n_102_26), .A (n_104_26), .B (n_106_25), .C1 (n_109_22), .C2 (n_115_19) );
AOI211_X1 g_104_25 (.ZN (n_104_25), .A (n_103_28), .B (n_105_23), .C1 (n_107_23), .C2 (n_113_20) );
AOI211_X1 g_106_24 (.ZN (n_106_24), .A (n_102_26), .B (n_103_24), .C1 (n_106_25), .C2 (n_111_21) );
AOI211_X1 g_107_22 (.ZN (n_107_22), .A (n_104_25), .B (n_104_26), .C1 (n_105_23), .C2 (n_109_22) );
AOI211_X1 g_109_21 (.ZN (n_109_21), .A (n_106_24), .B (n_103_28), .C1 (n_103_24), .C2 (n_107_23) );
AOI211_X1 g_111_20 (.ZN (n_111_20), .A (n_107_22), .B (n_102_26), .C1 (n_104_26), .C2 (n_106_25) );
AOI211_X1 g_113_19 (.ZN (n_113_19), .A (n_109_21), .B (n_104_25), .C1 (n_103_28), .C2 (n_105_23) );
AOI211_X1 g_115_18 (.ZN (n_115_18), .A (n_111_20), .B (n_106_24), .C1 (n_102_26), .C2 (n_103_24) );
AOI211_X1 g_114_20 (.ZN (n_114_20), .A (n_113_19), .B (n_107_22), .C1 (n_104_25), .C2 (n_104_26) );
AOI211_X1 g_116_19 (.ZN (n_116_19), .A (n_115_18), .B (n_109_21), .C1 (n_106_24), .C2 (n_103_28) );
AOI211_X1 g_118_18 (.ZN (n_118_18), .A (n_114_20), .B (n_111_20), .C1 (n_107_22), .C2 (n_102_26) );
AOI211_X1 g_120_17 (.ZN (n_120_17), .A (n_116_19), .B (n_113_19), .C1 (n_109_21), .C2 (n_104_25) );
AOI211_X1 g_122_16 (.ZN (n_122_16), .A (n_118_18), .B (n_115_18), .C1 (n_111_20), .C2 (n_106_24) );
AOI211_X1 g_124_15 (.ZN (n_124_15), .A (n_120_17), .B (n_114_20), .C1 (n_113_19), .C2 (n_107_22) );
AOI211_X1 g_126_14 (.ZN (n_126_14), .A (n_122_16), .B (n_116_19), .C1 (n_115_18), .C2 (n_109_21) );
AOI211_X1 g_128_13 (.ZN (n_128_13), .A (n_124_15), .B (n_118_18), .C1 (n_114_20), .C2 (n_111_20) );
AOI211_X1 g_127_15 (.ZN (n_127_15), .A (n_126_14), .B (n_120_17), .C1 (n_116_19), .C2 (n_113_19) );
AOI211_X1 g_125_16 (.ZN (n_125_16), .A (n_128_13), .B (n_122_16), .C1 (n_118_18), .C2 (n_115_18) );
AOI211_X1 g_123_17 (.ZN (n_123_17), .A (n_127_15), .B (n_124_15), .C1 (n_120_17), .C2 (n_114_20) );
AOI211_X1 g_121_18 (.ZN (n_121_18), .A (n_125_16), .B (n_126_14), .C1 (n_122_16), .C2 (n_116_19) );
AOI211_X1 g_119_19 (.ZN (n_119_19), .A (n_123_17), .B (n_128_13), .C1 (n_124_15), .C2 (n_118_18) );
AOI211_X1 g_117_20 (.ZN (n_117_20), .A (n_121_18), .B (n_127_15), .C1 (n_126_14), .C2 (n_120_17) );
AOI211_X1 g_115_21 (.ZN (n_115_21), .A (n_119_19), .B (n_125_16), .C1 (n_128_13), .C2 (n_122_16) );
AOI211_X1 g_113_22 (.ZN (n_113_22), .A (n_117_20), .B (n_123_17), .C1 (n_127_15), .C2 (n_124_15) );
AOI211_X1 g_111_23 (.ZN (n_111_23), .A (n_115_21), .B (n_121_18), .C1 (n_125_16), .C2 (n_126_14) );
AOI211_X1 g_112_21 (.ZN (n_112_21), .A (n_113_22), .B (n_119_19), .C1 (n_123_17), .C2 (n_128_13) );
AOI211_X1 g_110_22 (.ZN (n_110_22), .A (n_111_23), .B (n_117_20), .C1 (n_121_18), .C2 (n_127_15) );
AOI211_X1 g_108_23 (.ZN (n_108_23), .A (n_112_21), .B (n_115_21), .C1 (n_119_19), .C2 (n_125_16) );
AOI211_X1 g_107_25 (.ZN (n_107_25), .A (n_110_22), .B (n_113_22), .C1 (n_117_20), .C2 (n_123_17) );
AOI211_X1 g_109_24 (.ZN (n_109_24), .A (n_108_23), .B (n_111_23), .C1 (n_115_21), .C2 (n_121_18) );
AOI211_X1 g_108_26 (.ZN (n_108_26), .A (n_107_25), .B (n_112_21), .C1 (n_113_22), .C2 (n_119_19) );
AOI211_X1 g_107_24 (.ZN (n_107_24), .A (n_109_24), .B (n_110_22), .C1 (n_111_23), .C2 (n_117_20) );
AOI211_X1 g_109_23 (.ZN (n_109_23), .A (n_108_26), .B (n_108_23), .C1 (n_112_21), .C2 (n_115_21) );
AOI211_X1 g_111_22 (.ZN (n_111_22), .A (n_107_24), .B (n_107_25), .C1 (n_110_22), .C2 (n_113_22) );
AOI211_X1 g_113_21 (.ZN (n_113_21), .A (n_109_23), .B (n_109_24), .C1 (n_108_23), .C2 (n_111_23) );
AOI211_X1 g_115_20 (.ZN (n_115_20), .A (n_111_22), .B (n_108_26), .C1 (n_107_25), .C2 (n_112_21) );
AOI211_X1 g_117_19 (.ZN (n_117_19), .A (n_113_21), .B (n_107_24), .C1 (n_109_24), .C2 (n_110_22) );
AOI211_X1 g_119_18 (.ZN (n_119_18), .A (n_115_20), .B (n_109_23), .C1 (n_108_26), .C2 (n_108_23) );
AOI211_X1 g_121_17 (.ZN (n_121_17), .A (n_117_19), .B (n_111_22), .C1 (n_107_24), .C2 (n_107_25) );
AOI211_X1 g_120_19 (.ZN (n_120_19), .A (n_119_18), .B (n_113_21), .C1 (n_109_23), .C2 (n_109_24) );
AOI211_X1 g_122_18 (.ZN (n_122_18), .A (n_121_17), .B (n_115_20), .C1 (n_111_22), .C2 (n_108_26) );
AOI211_X1 g_124_17 (.ZN (n_124_17), .A (n_120_19), .B (n_117_19), .C1 (n_113_21), .C2 (n_107_24) );
AOI211_X1 g_126_16 (.ZN (n_126_16), .A (n_122_18), .B (n_119_18), .C1 (n_115_20), .C2 (n_109_23) );
AOI211_X1 g_128_15 (.ZN (n_128_15), .A (n_124_17), .B (n_121_17), .C1 (n_117_19), .C2 (n_111_22) );
AOI211_X1 g_130_14 (.ZN (n_130_14), .A (n_126_16), .B (n_120_19), .C1 (n_119_18), .C2 (n_113_21) );
AOI211_X1 g_129_16 (.ZN (n_129_16), .A (n_128_15), .B (n_122_18), .C1 (n_121_17), .C2 (n_115_20) );
AOI211_X1 g_131_15 (.ZN (n_131_15), .A (n_130_14), .B (n_124_17), .C1 (n_120_19), .C2 (n_117_19) );
AOI211_X1 g_133_16 (.ZN (n_133_16), .A (n_129_16), .B (n_126_16), .C1 (n_122_18), .C2 (n_119_18) );
AOI211_X1 g_131_17 (.ZN (n_131_17), .A (n_131_15), .B (n_128_15), .C1 (n_124_17), .C2 (n_121_17) );
AOI211_X1 g_132_15 (.ZN (n_132_15), .A (n_133_16), .B (n_130_14), .C1 (n_126_16), .C2 (n_120_19) );
AOI211_X1 g_133_13 (.ZN (n_133_13), .A (n_131_17), .B (n_129_16), .C1 (n_128_15), .C2 (n_122_18) );
AOI211_X1 g_131_14 (.ZN (n_131_14), .A (n_132_15), .B (n_131_15), .C1 (n_130_14), .C2 (n_124_17) );
AOI211_X1 g_129_15 (.ZN (n_129_15), .A (n_133_13), .B (n_133_16), .C1 (n_129_16), .C2 (n_126_16) );
AOI211_X1 g_127_16 (.ZN (n_127_16), .A (n_131_14), .B (n_131_17), .C1 (n_131_15), .C2 (n_128_15) );
AOI211_X1 g_125_17 (.ZN (n_125_17), .A (n_129_15), .B (n_132_15), .C1 (n_133_16), .C2 (n_130_14) );
AOI211_X1 g_123_18 (.ZN (n_123_18), .A (n_127_16), .B (n_133_13), .C1 (n_131_17), .C2 (n_129_16) );
AOI211_X1 g_121_19 (.ZN (n_121_19), .A (n_125_17), .B (n_131_14), .C1 (n_132_15), .C2 (n_131_15) );
AOI211_X1 g_119_20 (.ZN (n_119_20), .A (n_123_18), .B (n_129_15), .C1 (n_133_13), .C2 (n_133_16) );
AOI211_X1 g_117_21 (.ZN (n_117_21), .A (n_121_19), .B (n_127_16), .C1 (n_131_14), .C2 (n_131_17) );
AOI211_X1 g_118_19 (.ZN (n_118_19), .A (n_119_20), .B (n_125_17), .C1 (n_129_15), .C2 (n_132_15) );
AOI211_X1 g_116_20 (.ZN (n_116_20), .A (n_117_21), .B (n_123_18), .C1 (n_127_16), .C2 (n_133_13) );
AOI211_X1 g_114_21 (.ZN (n_114_21), .A (n_118_19), .B (n_121_19), .C1 (n_125_17), .C2 (n_131_14) );
AOI211_X1 g_112_22 (.ZN (n_112_22), .A (n_116_20), .B (n_119_20), .C1 (n_123_18), .C2 (n_129_15) );
AOI211_X1 g_110_23 (.ZN (n_110_23), .A (n_114_21), .B (n_117_21), .C1 (n_121_19), .C2 (n_127_16) );
AOI211_X1 g_108_24 (.ZN (n_108_24), .A (n_112_22), .B (n_118_19), .C1 (n_119_20), .C2 (n_125_17) );
AOI211_X1 g_110_25 (.ZN (n_110_25), .A (n_110_23), .B (n_116_20), .C1 (n_117_21), .C2 (n_123_18) );
AOI211_X1 g_112_24 (.ZN (n_112_24), .A (n_108_24), .B (n_114_21), .C1 (n_118_19), .C2 (n_121_19) );
AOI211_X1 g_114_23 (.ZN (n_114_23), .A (n_110_25), .B (n_112_22), .C1 (n_116_20), .C2 (n_119_20) );
AOI211_X1 g_116_22 (.ZN (n_116_22), .A (n_112_24), .B (n_110_23), .C1 (n_114_21), .C2 (n_117_21) );
AOI211_X1 g_118_21 (.ZN (n_118_21), .A (n_114_23), .B (n_108_24), .C1 (n_112_22), .C2 (n_118_19) );
AOI211_X1 g_120_20 (.ZN (n_120_20), .A (n_116_22), .B (n_110_25), .C1 (n_110_23), .C2 (n_116_20) );
AOI211_X1 g_122_19 (.ZN (n_122_19), .A (n_118_21), .B (n_112_24), .C1 (n_108_24), .C2 (n_114_21) );
AOI211_X1 g_124_18 (.ZN (n_124_18), .A (n_120_20), .B (n_114_23), .C1 (n_110_25), .C2 (n_112_22) );
AOI211_X1 g_126_17 (.ZN (n_126_17), .A (n_122_19), .B (n_116_22), .C1 (n_112_24), .C2 (n_110_23) );
AOI211_X1 g_128_16 (.ZN (n_128_16), .A (n_124_18), .B (n_118_21), .C1 (n_114_23), .C2 (n_108_24) );
AOI211_X1 g_127_18 (.ZN (n_127_18), .A (n_126_17), .B (n_120_20), .C1 (n_116_22), .C2 (n_110_25) );
AOI211_X1 g_129_17 (.ZN (n_129_17), .A (n_128_16), .B (n_122_19), .C1 (n_118_21), .C2 (n_112_24) );
AOI211_X1 g_131_16 (.ZN (n_131_16), .A (n_127_18), .B (n_124_18), .C1 (n_120_20), .C2 (n_114_23) );
AOI211_X1 g_133_15 (.ZN (n_133_15), .A (n_129_17), .B (n_126_17), .C1 (n_122_19), .C2 (n_116_22) );
AOI211_X1 g_135_14 (.ZN (n_135_14), .A (n_131_16), .B (n_128_16), .C1 (n_124_18), .C2 (n_118_21) );
AOI211_X1 g_134_16 (.ZN (n_134_16), .A (n_133_15), .B (n_127_18), .C1 (n_126_17), .C2 (n_120_20) );
AOI211_X1 g_132_17 (.ZN (n_132_17), .A (n_135_14), .B (n_129_17), .C1 (n_128_16), .C2 (n_122_19) );
AOI211_X1 g_130_16 (.ZN (n_130_16), .A (n_134_16), .B (n_131_16), .C1 (n_127_18), .C2 (n_124_18) );
AOI211_X1 g_128_17 (.ZN (n_128_17), .A (n_132_17), .B (n_133_15), .C1 (n_129_17), .C2 (n_126_17) );
AOI211_X1 g_126_18 (.ZN (n_126_18), .A (n_130_16), .B (n_135_14), .C1 (n_131_16), .C2 (n_128_16) );
AOI211_X1 g_124_19 (.ZN (n_124_19), .A (n_128_17), .B (n_134_16), .C1 (n_133_15), .C2 (n_127_18) );
AOI211_X1 g_122_20 (.ZN (n_122_20), .A (n_126_18), .B (n_132_17), .C1 (n_135_14), .C2 (n_129_17) );
AOI211_X1 g_120_21 (.ZN (n_120_21), .A (n_124_19), .B (n_130_16), .C1 (n_134_16), .C2 (n_131_16) );
AOI211_X1 g_118_20 (.ZN (n_118_20), .A (n_122_20), .B (n_128_17), .C1 (n_132_17), .C2 (n_133_15) );
AOI211_X1 g_116_21 (.ZN (n_116_21), .A (n_120_21), .B (n_126_18), .C1 (n_130_16), .C2 (n_135_14) );
AOI211_X1 g_114_22 (.ZN (n_114_22), .A (n_118_20), .B (n_124_19), .C1 (n_128_17), .C2 (n_134_16) );
AOI211_X1 g_112_23 (.ZN (n_112_23), .A (n_116_21), .B (n_122_20), .C1 (n_126_18), .C2 (n_132_17) );
AOI211_X1 g_110_24 (.ZN (n_110_24), .A (n_114_22), .B (n_120_21), .C1 (n_124_19), .C2 (n_130_16) );
AOI211_X1 g_108_25 (.ZN (n_108_25), .A (n_112_23), .B (n_118_20), .C1 (n_122_20), .C2 (n_128_17) );
AOI211_X1 g_106_26 (.ZN (n_106_26), .A (n_110_24), .B (n_116_21), .C1 (n_120_21), .C2 (n_126_18) );
AOI211_X1 g_104_27 (.ZN (n_104_27), .A (n_108_25), .B (n_114_22), .C1 (n_118_20), .C2 (n_124_19) );
AOI211_X1 g_105_25 (.ZN (n_105_25), .A (n_106_26), .B (n_112_23), .C1 (n_116_21), .C2 (n_122_20) );
AOI211_X1 g_103_26 (.ZN (n_103_26), .A (n_104_27), .B (n_110_24), .C1 (n_114_22), .C2 (n_120_21) );
AOI211_X1 g_101_27 (.ZN (n_101_27), .A (n_105_25), .B (n_108_25), .C1 (n_112_23), .C2 (n_118_20) );
AOI211_X1 g_99_28 (.ZN (n_99_28), .A (n_103_26), .B (n_106_26), .C1 (n_110_24), .C2 (n_116_21) );
AOI211_X1 g_97_29 (.ZN (n_97_29), .A (n_101_27), .B (n_104_27), .C1 (n_108_25), .C2 (n_114_22) );
AOI211_X1 g_95_30 (.ZN (n_95_30), .A (n_99_28), .B (n_105_25), .C1 (n_106_26), .C2 (n_112_23) );
AOI211_X1 g_93_31 (.ZN (n_93_31), .A (n_97_29), .B (n_103_26), .C1 (n_104_27), .C2 (n_110_24) );
AOI211_X1 g_91_32 (.ZN (n_91_32), .A (n_95_30), .B (n_101_27), .C1 (n_105_25), .C2 (n_108_25) );
AOI211_X1 g_89_33 (.ZN (n_89_33), .A (n_93_31), .B (n_99_28), .C1 (n_103_26), .C2 (n_106_26) );
AOI211_X1 g_87_34 (.ZN (n_87_34), .A (n_91_32), .B (n_97_29), .C1 (n_101_27), .C2 (n_104_27) );
AOI211_X1 g_85_35 (.ZN (n_85_35), .A (n_89_33), .B (n_95_30), .C1 (n_99_28), .C2 (n_105_25) );
AOI211_X1 g_83_36 (.ZN (n_83_36), .A (n_87_34), .B (n_93_31), .C1 (n_97_29), .C2 (n_103_26) );
AOI211_X1 g_81_37 (.ZN (n_81_37), .A (n_85_35), .B (n_91_32), .C1 (n_95_30), .C2 (n_101_27) );
AOI211_X1 g_79_38 (.ZN (n_79_38), .A (n_83_36), .B (n_89_33), .C1 (n_93_31), .C2 (n_99_28) );
AOI211_X1 g_77_39 (.ZN (n_77_39), .A (n_81_37), .B (n_87_34), .C1 (n_91_32), .C2 (n_97_29) );
AOI211_X1 g_75_40 (.ZN (n_75_40), .A (n_79_38), .B (n_85_35), .C1 (n_89_33), .C2 (n_95_30) );
AOI211_X1 g_73_41 (.ZN (n_73_41), .A (n_77_39), .B (n_83_36), .C1 (n_87_34), .C2 (n_93_31) );
AOI211_X1 g_71_42 (.ZN (n_71_42), .A (n_75_40), .B (n_81_37), .C1 (n_85_35), .C2 (n_91_32) );
AOI211_X1 g_69_43 (.ZN (n_69_43), .A (n_73_41), .B (n_79_38), .C1 (n_83_36), .C2 (n_89_33) );
AOI211_X1 g_67_44 (.ZN (n_67_44), .A (n_71_42), .B (n_77_39), .C1 (n_81_37), .C2 (n_87_34) );
AOI211_X1 g_65_45 (.ZN (n_65_45), .A (n_69_43), .B (n_75_40), .C1 (n_79_38), .C2 (n_85_35) );
AOI211_X1 g_63_46 (.ZN (n_63_46), .A (n_67_44), .B (n_73_41), .C1 (n_77_39), .C2 (n_83_36) );
AOI211_X1 g_61_47 (.ZN (n_61_47), .A (n_65_45), .B (n_71_42), .C1 (n_75_40), .C2 (n_81_37) );
AOI211_X1 g_59_48 (.ZN (n_59_48), .A (n_63_46), .B (n_69_43), .C1 (n_73_41), .C2 (n_79_38) );
AOI211_X1 g_57_49 (.ZN (n_57_49), .A (n_61_47), .B (n_67_44), .C1 (n_71_42), .C2 (n_77_39) );
AOI211_X1 g_55_50 (.ZN (n_55_50), .A (n_59_48), .B (n_65_45), .C1 (n_69_43), .C2 (n_75_40) );
AOI211_X1 g_53_51 (.ZN (n_53_51), .A (n_57_49), .B (n_63_46), .C1 (n_67_44), .C2 (n_73_41) );
AOI211_X1 g_51_52 (.ZN (n_51_52), .A (n_55_50), .B (n_61_47), .C1 (n_65_45), .C2 (n_71_42) );
AOI211_X1 g_49_53 (.ZN (n_49_53), .A (n_53_51), .B (n_59_48), .C1 (n_63_46), .C2 (n_69_43) );
AOI211_X1 g_47_54 (.ZN (n_47_54), .A (n_51_52), .B (n_57_49), .C1 (n_61_47), .C2 (n_67_44) );
AOI211_X1 g_45_55 (.ZN (n_45_55), .A (n_49_53), .B (n_55_50), .C1 (n_59_48), .C2 (n_65_45) );
AOI211_X1 g_43_56 (.ZN (n_43_56), .A (n_47_54), .B (n_53_51), .C1 (n_57_49), .C2 (n_63_46) );
AOI211_X1 g_41_57 (.ZN (n_41_57), .A (n_45_55), .B (n_51_52), .C1 (n_55_50), .C2 (n_61_47) );
AOI211_X1 g_39_56 (.ZN (n_39_56), .A (n_43_56), .B (n_49_53), .C1 (n_53_51), .C2 (n_59_48) );
AOI211_X1 g_37_57 (.ZN (n_37_57), .A (n_41_57), .B (n_47_54), .C1 (n_51_52), .C2 (n_57_49) );
AOI211_X1 g_35_58 (.ZN (n_35_58), .A (n_39_56), .B (n_45_55), .C1 (n_49_53), .C2 (n_55_50) );
AOI211_X1 g_33_59 (.ZN (n_33_59), .A (n_37_57), .B (n_43_56), .C1 (n_47_54), .C2 (n_53_51) );
AOI211_X1 g_31_60 (.ZN (n_31_60), .A (n_35_58), .B (n_41_57), .C1 (n_45_55), .C2 (n_51_52) );
AOI211_X1 g_29_61 (.ZN (n_29_61), .A (n_33_59), .B (n_39_56), .C1 (n_43_56), .C2 (n_49_53) );
AOI211_X1 g_27_62 (.ZN (n_27_62), .A (n_31_60), .B (n_37_57), .C1 (n_41_57), .C2 (n_47_54) );
AOI211_X1 g_25_63 (.ZN (n_25_63), .A (n_29_61), .B (n_35_58), .C1 (n_39_56), .C2 (n_45_55) );
AOI211_X1 g_23_64 (.ZN (n_23_64), .A (n_27_62), .B (n_33_59), .C1 (n_37_57), .C2 (n_43_56) );
AOI211_X1 g_21_65 (.ZN (n_21_65), .A (n_25_63), .B (n_31_60), .C1 (n_35_58), .C2 (n_41_57) );
AOI211_X1 g_19_66 (.ZN (n_19_66), .A (n_23_64), .B (n_29_61), .C1 (n_33_59), .C2 (n_39_56) );
AOI211_X1 g_17_65 (.ZN (n_17_65), .A (n_21_65), .B (n_27_62), .C1 (n_31_60), .C2 (n_37_57) );
AOI211_X1 g_15_66 (.ZN (n_15_66), .A (n_19_66), .B (n_25_63), .C1 (n_29_61), .C2 (n_35_58) );
AOI211_X1 g_13_67 (.ZN (n_13_67), .A (n_17_65), .B (n_23_64), .C1 (n_27_62), .C2 (n_33_59) );
AOI211_X1 g_11_68 (.ZN (n_11_68), .A (n_15_66), .B (n_21_65), .C1 (n_25_63), .C2 (n_31_60) );
AOI211_X1 g_9_69 (.ZN (n_9_69), .A (n_13_67), .B (n_19_66), .C1 (n_23_64), .C2 (n_29_61) );
AOI211_X1 g_8_71 (.ZN (n_8_71), .A (n_11_68), .B (n_17_65), .C1 (n_21_65), .C2 (n_27_62) );
AOI211_X1 g_6_70 (.ZN (n_6_70), .A (n_9_69), .B (n_15_66), .C1 (n_19_66), .C2 (n_25_63) );
AOI211_X1 g_8_69 (.ZN (n_8_69), .A (n_8_71), .B (n_13_67), .C1 (n_17_65), .C2 (n_23_64) );
AOI211_X1 g_10_68 (.ZN (n_10_68), .A (n_6_70), .B (n_11_68), .C1 (n_15_66), .C2 (n_21_65) );
AOI211_X1 g_12_67 (.ZN (n_12_67), .A (n_8_69), .B (n_9_69), .C1 (n_13_67), .C2 (n_19_66) );
AOI211_X1 g_14_66 (.ZN (n_14_66), .A (n_10_68), .B (n_8_71), .C1 (n_11_68), .C2 (n_17_65) );
AOI211_X1 g_16_65 (.ZN (n_16_65), .A (n_12_67), .B (n_6_70), .C1 (n_9_69), .C2 (n_15_66) );
AOI211_X1 g_17_67 (.ZN (n_17_67), .A (n_14_66), .B (n_8_69), .C1 (n_8_71), .C2 (n_13_67) );
AOI211_X1 g_15_68 (.ZN (n_15_68), .A (n_16_65), .B (n_10_68), .C1 (n_6_70), .C2 (n_11_68) );
AOI211_X1 g_13_69 (.ZN (n_13_69), .A (n_17_67), .B (n_12_67), .C1 (n_8_69), .C2 (n_9_69) );
AOI211_X1 g_11_70 (.ZN (n_11_70), .A (n_15_68), .B (n_14_66), .C1 (n_10_68), .C2 (n_8_71) );
AOI211_X1 g_9_71 (.ZN (n_9_71), .A (n_13_69), .B (n_16_65), .C1 (n_12_67), .C2 (n_6_70) );
AOI211_X1 g_10_69 (.ZN (n_10_69), .A (n_11_70), .B (n_17_67), .C1 (n_14_66), .C2 (n_8_69) );
AOI211_X1 g_8_70 (.ZN (n_8_70), .A (n_9_71), .B (n_15_68), .C1 (n_16_65), .C2 (n_10_68) );
AOI211_X1 g_6_69 (.ZN (n_6_69), .A (n_10_69), .B (n_13_69), .C1 (n_17_67), .C2 (n_12_67) );
AOI211_X1 g_4_70 (.ZN (n_4_70), .A (n_8_70), .B (n_11_70), .C1 (n_15_68), .C2 (n_14_66) );
AOI211_X1 g_3_72 (.ZN (n_3_72), .A (n_6_69), .B (n_9_71), .C1 (n_13_69), .C2 (n_16_65) );
AOI211_X1 g_5_71 (.ZN (n_5_71), .A (n_4_70), .B (n_10_69), .C1 (n_11_70), .C2 (n_17_67) );
AOI211_X1 g_7_72 (.ZN (n_7_72), .A (n_3_72), .B (n_8_70), .C1 (n_9_71), .C2 (n_15_68) );
AOI211_X1 g_5_73 (.ZN (n_5_73), .A (n_5_71), .B (n_6_69), .C1 (n_10_69), .C2 (n_13_69) );
AOI211_X1 g_6_71 (.ZN (n_6_71), .A (n_7_72), .B (n_4_70), .C1 (n_8_70), .C2 (n_11_70) );
AOI211_X1 g_7_73 (.ZN (n_7_73), .A (n_5_73), .B (n_3_72), .C1 (n_6_69), .C2 (n_9_71) );
AOI211_X1 g_5_72 (.ZN (n_5_72), .A (n_6_71), .B (n_5_71), .C1 (n_4_70), .C2 (n_10_69) );
AOI211_X1 g_7_71 (.ZN (n_7_71), .A (n_7_73), .B (n_7_72), .C1 (n_3_72), .C2 (n_8_70) );
AOI211_X1 g_9_70 (.ZN (n_9_70), .A (n_5_72), .B (n_5_73), .C1 (n_5_71), .C2 (n_6_69) );
AOI211_X1 g_11_69 (.ZN (n_11_69), .A (n_7_71), .B (n_6_71), .C1 (n_7_72), .C2 (n_4_70) );
AOI211_X1 g_13_68 (.ZN (n_13_68), .A (n_9_70), .B (n_7_73), .C1 (n_5_73), .C2 (n_3_72) );
AOI211_X1 g_15_67 (.ZN (n_15_67), .A (n_11_69), .B (n_5_72), .C1 (n_6_71), .C2 (n_5_71) );
AOI211_X1 g_17_66 (.ZN (n_17_66), .A (n_13_68), .B (n_7_71), .C1 (n_7_73), .C2 (n_7_72) );
AOI211_X1 g_16_68 (.ZN (n_16_68), .A (n_15_67), .B (n_9_70), .C1 (n_5_72), .C2 (n_5_73) );
AOI211_X1 g_18_67 (.ZN (n_18_67), .A (n_17_66), .B (n_11_69), .C1 (n_7_71), .C2 (n_6_71) );
AOI211_X1 g_17_69 (.ZN (n_17_69), .A (n_16_68), .B (n_13_68), .C1 (n_9_70), .C2 (n_7_73) );
AOI211_X1 g_19_68 (.ZN (n_19_68), .A (n_18_67), .B (n_15_67), .C1 (n_11_69), .C2 (n_5_72) );
AOI211_X1 g_18_66 (.ZN (n_18_66), .A (n_17_69), .B (n_17_66), .C1 (n_13_68), .C2 (n_7_71) );
AOI211_X1 g_16_67 (.ZN (n_16_67), .A (n_19_68), .B (n_16_68), .C1 (n_15_67), .C2 (n_9_70) );
AOI211_X1 g_14_68 (.ZN (n_14_68), .A (n_18_66), .B (n_18_67), .C1 (n_17_66), .C2 (n_11_69) );
AOI211_X1 g_12_69 (.ZN (n_12_69), .A (n_16_67), .B (n_17_69), .C1 (n_16_68), .C2 (n_13_68) );
AOI211_X1 g_10_70 (.ZN (n_10_70), .A (n_14_68), .B (n_19_68), .C1 (n_18_67), .C2 (n_15_67) );
AOI211_X1 g_9_72 (.ZN (n_9_72), .A (n_12_69), .B (n_18_66), .C1 (n_17_69), .C2 (n_17_66) );
AOI211_X1 g_11_71 (.ZN (n_11_71), .A (n_10_70), .B (n_16_67), .C1 (n_19_68), .C2 (n_16_68) );
AOI211_X1 g_13_70 (.ZN (n_13_70), .A (n_9_72), .B (n_14_68), .C1 (n_18_66), .C2 (n_18_67) );
AOI211_X1 g_15_69 (.ZN (n_15_69), .A (n_11_71), .B (n_12_69), .C1 (n_16_67), .C2 (n_17_69) );
AOI211_X1 g_17_68 (.ZN (n_17_68), .A (n_13_70), .B (n_10_70), .C1 (n_14_68), .C2 (n_19_68) );
AOI211_X1 g_19_67 (.ZN (n_19_67), .A (n_15_69), .B (n_9_72), .C1 (n_12_69), .C2 (n_18_66) );
AOI211_X1 g_21_66 (.ZN (n_21_66), .A (n_17_68), .B (n_11_71), .C1 (n_10_70), .C2 (n_16_67) );
AOI211_X1 g_23_65 (.ZN (n_23_65), .A (n_19_67), .B (n_13_70), .C1 (n_9_72), .C2 (n_14_68) );
AOI211_X1 g_22_67 (.ZN (n_22_67), .A (n_21_66), .B (n_15_69), .C1 (n_11_71), .C2 (n_12_69) );
AOI211_X1 g_24_66 (.ZN (n_24_66), .A (n_23_65), .B (n_17_68), .C1 (n_13_70), .C2 (n_10_70) );
AOI211_X1 g_26_65 (.ZN (n_26_65), .A (n_22_67), .B (n_19_67), .C1 (n_15_69), .C2 (n_9_72) );
AOI211_X1 g_28_64 (.ZN (n_28_64), .A (n_24_66), .B (n_21_66), .C1 (n_17_68), .C2 (n_11_71) );
AOI211_X1 g_30_63 (.ZN (n_30_63), .A (n_26_65), .B (n_23_65), .C1 (n_19_67), .C2 (n_13_70) );
AOI211_X1 g_32_62 (.ZN (n_32_62), .A (n_28_64), .B (n_22_67), .C1 (n_21_66), .C2 (n_15_69) );
AOI211_X1 g_34_61 (.ZN (n_34_61), .A (n_30_63), .B (n_24_66), .C1 (n_23_65), .C2 (n_17_68) );
AOI211_X1 g_36_60 (.ZN (n_36_60), .A (n_32_62), .B (n_26_65), .C1 (n_22_67), .C2 (n_19_67) );
AOI211_X1 g_38_59 (.ZN (n_38_59), .A (n_34_61), .B (n_28_64), .C1 (n_24_66), .C2 (n_21_66) );
AOI211_X1 g_40_58 (.ZN (n_40_58), .A (n_36_60), .B (n_30_63), .C1 (n_26_65), .C2 (n_23_65) );
AOI211_X1 g_42_57 (.ZN (n_42_57), .A (n_38_59), .B (n_32_62), .C1 (n_28_64), .C2 (n_22_67) );
AOI211_X1 g_44_56 (.ZN (n_44_56), .A (n_40_58), .B (n_34_61), .C1 (n_30_63), .C2 (n_24_66) );
AOI211_X1 g_46_55 (.ZN (n_46_55), .A (n_42_57), .B (n_36_60), .C1 (n_32_62), .C2 (n_26_65) );
AOI211_X1 g_48_54 (.ZN (n_48_54), .A (n_44_56), .B (n_38_59), .C1 (n_34_61), .C2 (n_28_64) );
AOI211_X1 g_50_53 (.ZN (n_50_53), .A (n_46_55), .B (n_40_58), .C1 (n_36_60), .C2 (n_30_63) );
AOI211_X1 g_52_52 (.ZN (n_52_52), .A (n_48_54), .B (n_42_57), .C1 (n_38_59), .C2 (n_32_62) );
AOI211_X1 g_54_51 (.ZN (n_54_51), .A (n_50_53), .B (n_44_56), .C1 (n_40_58), .C2 (n_34_61) );
AOI211_X1 g_56_50 (.ZN (n_56_50), .A (n_52_52), .B (n_46_55), .C1 (n_42_57), .C2 (n_36_60) );
AOI211_X1 g_58_49 (.ZN (n_58_49), .A (n_54_51), .B (n_48_54), .C1 (n_44_56), .C2 (n_38_59) );
AOI211_X1 g_60_48 (.ZN (n_60_48), .A (n_56_50), .B (n_50_53), .C1 (n_46_55), .C2 (n_40_58) );
AOI211_X1 g_59_50 (.ZN (n_59_50), .A (n_58_49), .B (n_52_52), .C1 (n_48_54), .C2 (n_42_57) );
AOI211_X1 g_61_49 (.ZN (n_61_49), .A (n_60_48), .B (n_54_51), .C1 (n_50_53), .C2 (n_44_56) );
AOI211_X1 g_63_48 (.ZN (n_63_48), .A (n_59_50), .B (n_56_50), .C1 (n_52_52), .C2 (n_46_55) );
AOI211_X1 g_65_47 (.ZN (n_65_47), .A (n_61_49), .B (n_58_49), .C1 (n_54_51), .C2 (n_48_54) );
AOI211_X1 g_67_46 (.ZN (n_67_46), .A (n_63_48), .B (n_60_48), .C1 (n_56_50), .C2 (n_50_53) );
AOI211_X1 g_68_44 (.ZN (n_68_44), .A (n_65_47), .B (n_59_50), .C1 (n_58_49), .C2 (n_52_52) );
AOI211_X1 g_70_43 (.ZN (n_70_43), .A (n_67_46), .B (n_61_49), .C1 (n_60_48), .C2 (n_54_51) );
AOI211_X1 g_72_42 (.ZN (n_72_42), .A (n_68_44), .B (n_63_48), .C1 (n_59_50), .C2 (n_56_50) );
AOI211_X1 g_74_41 (.ZN (n_74_41), .A (n_70_43), .B (n_65_47), .C1 (n_61_49), .C2 (n_58_49) );
AOI211_X1 g_76_40 (.ZN (n_76_40), .A (n_72_42), .B (n_67_46), .C1 (n_63_48), .C2 (n_60_48) );
AOI211_X1 g_78_39 (.ZN (n_78_39), .A (n_74_41), .B (n_68_44), .C1 (n_65_47), .C2 (n_59_50) );
AOI211_X1 g_80_38 (.ZN (n_80_38), .A (n_76_40), .B (n_70_43), .C1 (n_67_46), .C2 (n_61_49) );
AOI211_X1 g_82_37 (.ZN (n_82_37), .A (n_78_39), .B (n_72_42), .C1 (n_68_44), .C2 (n_63_48) );
AOI211_X1 g_84_36 (.ZN (n_84_36), .A (n_80_38), .B (n_74_41), .C1 (n_70_43), .C2 (n_65_47) );
AOI211_X1 g_86_35 (.ZN (n_86_35), .A (n_82_37), .B (n_76_40), .C1 (n_72_42), .C2 (n_67_46) );
AOI211_X1 g_88_34 (.ZN (n_88_34), .A (n_84_36), .B (n_78_39), .C1 (n_74_41), .C2 (n_68_44) );
AOI211_X1 g_90_33 (.ZN (n_90_33), .A (n_86_35), .B (n_80_38), .C1 (n_76_40), .C2 (n_70_43) );
AOI211_X1 g_89_35 (.ZN (n_89_35), .A (n_88_34), .B (n_82_37), .C1 (n_78_39), .C2 (n_72_42) );
AOI211_X1 g_87_36 (.ZN (n_87_36), .A (n_90_33), .B (n_84_36), .C1 (n_80_38), .C2 (n_74_41) );
AOI211_X1 g_85_37 (.ZN (n_85_37), .A (n_89_35), .B (n_86_35), .C1 (n_82_37), .C2 (n_76_40) );
AOI211_X1 g_83_38 (.ZN (n_83_38), .A (n_87_36), .B (n_88_34), .C1 (n_84_36), .C2 (n_78_39) );
AOI211_X1 g_81_39 (.ZN (n_81_39), .A (n_85_37), .B (n_90_33), .C1 (n_86_35), .C2 (n_80_38) );
AOI211_X1 g_79_40 (.ZN (n_79_40), .A (n_83_38), .B (n_89_35), .C1 (n_88_34), .C2 (n_82_37) );
AOI211_X1 g_77_41 (.ZN (n_77_41), .A (n_81_39), .B (n_87_36), .C1 (n_90_33), .C2 (n_84_36) );
AOI211_X1 g_75_42 (.ZN (n_75_42), .A (n_79_40), .B (n_85_37), .C1 (n_89_35), .C2 (n_86_35) );
AOI211_X1 g_73_43 (.ZN (n_73_43), .A (n_77_41), .B (n_83_38), .C1 (n_87_36), .C2 (n_88_34) );
AOI211_X1 g_71_44 (.ZN (n_71_44), .A (n_75_42), .B (n_81_39), .C1 (n_85_37), .C2 (n_90_33) );
AOI211_X1 g_70_42 (.ZN (n_70_42), .A (n_73_43), .B (n_79_40), .C1 (n_83_38), .C2 (n_89_35) );
AOI211_X1 g_68_43 (.ZN (n_68_43), .A (n_71_44), .B (n_77_41), .C1 (n_81_39), .C2 (n_87_36) );
AOI211_X1 g_69_45 (.ZN (n_69_45), .A (n_70_42), .B (n_75_42), .C1 (n_79_40), .C2 (n_85_37) );
AOI211_X1 g_68_47 (.ZN (n_68_47), .A (n_68_43), .B (n_73_43), .C1 (n_77_41), .C2 (n_83_38) );
AOI211_X1 g_67_45 (.ZN (n_67_45), .A (n_69_45), .B (n_71_44), .C1 (n_75_42), .C2 (n_81_39) );
AOI211_X1 g_69_44 (.ZN (n_69_44), .A (n_68_47), .B (n_70_42), .C1 (n_73_43), .C2 (n_79_40) );
AOI211_X1 g_71_43 (.ZN (n_71_43), .A (n_67_45), .B (n_68_43), .C1 (n_71_44), .C2 (n_77_41) );
AOI211_X1 g_73_42 (.ZN (n_73_42), .A (n_69_44), .B (n_69_45), .C1 (n_70_42), .C2 (n_75_42) );
AOI211_X1 g_75_41 (.ZN (n_75_41), .A (n_71_43), .B (n_68_47), .C1 (n_68_43), .C2 (n_73_43) );
AOI211_X1 g_77_40 (.ZN (n_77_40), .A (n_73_42), .B (n_67_45), .C1 (n_69_45), .C2 (n_71_44) );
AOI211_X1 g_79_39 (.ZN (n_79_39), .A (n_75_41), .B (n_69_44), .C1 (n_68_47), .C2 (n_70_42) );
AOI211_X1 g_81_38 (.ZN (n_81_38), .A (n_77_40), .B (n_71_43), .C1 (n_67_45), .C2 (n_68_43) );
AOI211_X1 g_83_37 (.ZN (n_83_37), .A (n_79_39), .B (n_73_42), .C1 (n_69_44), .C2 (n_69_45) );
AOI211_X1 g_85_36 (.ZN (n_85_36), .A (n_81_38), .B (n_75_41), .C1 (n_71_43), .C2 (n_68_47) );
AOI211_X1 g_87_35 (.ZN (n_87_35), .A (n_83_37), .B (n_77_40), .C1 (n_73_42), .C2 (n_67_45) );
AOI211_X1 g_89_34 (.ZN (n_89_34), .A (n_85_36), .B (n_79_39), .C1 (n_75_41), .C2 (n_69_44) );
AOI211_X1 g_90_32 (.ZN (n_90_32), .A (n_87_35), .B (n_81_38), .C1 (n_77_40), .C2 (n_71_43) );
AOI211_X1 g_92_31 (.ZN (n_92_31), .A (n_89_34), .B (n_83_37), .C1 (n_79_39), .C2 (n_73_42) );
AOI211_X1 g_94_30 (.ZN (n_94_30), .A (n_90_32), .B (n_85_36), .C1 (n_81_38), .C2 (n_75_41) );
AOI211_X1 g_96_29 (.ZN (n_96_29), .A (n_92_31), .B (n_87_35), .C1 (n_83_37), .C2 (n_77_40) );
AOI211_X1 g_98_28 (.ZN (n_98_28), .A (n_94_30), .B (n_89_34), .C1 (n_85_36), .C2 (n_79_39) );
AOI211_X1 g_100_27 (.ZN (n_100_27), .A (n_96_29), .B (n_90_32), .C1 (n_87_35), .C2 (n_81_38) );
AOI211_X1 g_101_29 (.ZN (n_101_29), .A (n_98_28), .B (n_92_31), .C1 (n_89_34), .C2 (n_83_37) );
AOI211_X1 g_99_30 (.ZN (n_99_30), .A (n_100_27), .B (n_94_30), .C1 (n_90_32), .C2 (n_85_36) );
AOI211_X1 g_97_31 (.ZN (n_97_31), .A (n_101_29), .B (n_96_29), .C1 (n_92_31), .C2 (n_87_35) );
AOI211_X1 g_95_32 (.ZN (n_95_32), .A (n_99_30), .B (n_98_28), .C1 (n_94_30), .C2 (n_89_34) );
AOI211_X1 g_93_33 (.ZN (n_93_33), .A (n_97_31), .B (n_100_27), .C1 (n_96_29), .C2 (n_90_32) );
AOI211_X1 g_91_34 (.ZN (n_91_34), .A (n_95_32), .B (n_101_29), .C1 (n_98_28), .C2 (n_92_31) );
AOI211_X1 g_90_36 (.ZN (n_90_36), .A (n_93_33), .B (n_99_30), .C1 (n_100_27), .C2 (n_94_30) );
AOI211_X1 g_88_35 (.ZN (n_88_35), .A (n_91_34), .B (n_97_31), .C1 (n_101_29), .C2 (n_96_29) );
AOI211_X1 g_90_34 (.ZN (n_90_34), .A (n_90_36), .B (n_95_32), .C1 (n_99_30), .C2 (n_98_28) );
AOI211_X1 g_92_33 (.ZN (n_92_33), .A (n_88_35), .B (n_93_33), .C1 (n_97_31), .C2 (n_100_27) );
AOI211_X1 g_94_32 (.ZN (n_94_32), .A (n_90_34), .B (n_91_34), .C1 (n_95_32), .C2 (n_101_29) );
AOI211_X1 g_96_31 (.ZN (n_96_31), .A (n_92_33), .B (n_90_36), .C1 (n_93_33), .C2 (n_99_30) );
AOI211_X1 g_98_30 (.ZN (n_98_30), .A (n_94_32), .B (n_88_35), .C1 (n_91_34), .C2 (n_97_31) );
AOI211_X1 g_100_29 (.ZN (n_100_29), .A (n_96_31), .B (n_90_34), .C1 (n_90_36), .C2 (n_95_32) );
AOI211_X1 g_102_28 (.ZN (n_102_28), .A (n_98_30), .B (n_92_33), .C1 (n_88_35), .C2 (n_93_33) );
AOI211_X1 g_101_30 (.ZN (n_101_30), .A (n_100_29), .B (n_94_32), .C1 (n_90_34), .C2 (n_91_34) );
AOI211_X1 g_99_29 (.ZN (n_99_29), .A (n_102_28), .B (n_96_31), .C1 (n_92_33), .C2 (n_90_36) );
AOI211_X1 g_101_28 (.ZN (n_101_28), .A (n_101_30), .B (n_98_30), .C1 (n_94_32), .C2 (n_88_35) );
AOI211_X1 g_103_27 (.ZN (n_103_27), .A (n_99_29), .B (n_100_29), .C1 (n_96_31), .C2 (n_90_34) );
AOI211_X1 g_105_26 (.ZN (n_105_26), .A (n_101_28), .B (n_102_28), .C1 (n_98_30), .C2 (n_92_33) );
AOI211_X1 g_104_28 (.ZN (n_104_28), .A (n_103_27), .B (n_101_30), .C1 (n_100_29), .C2 (n_94_32) );
AOI211_X1 g_106_27 (.ZN (n_106_27), .A (n_105_26), .B (n_99_29), .C1 (n_102_28), .C2 (n_96_31) );
AOI211_X1 g_105_29 (.ZN (n_105_29), .A (n_104_28), .B (n_101_28), .C1 (n_101_30), .C2 (n_98_30) );
AOI211_X1 g_103_30 (.ZN (n_103_30), .A (n_106_27), .B (n_103_27), .C1 (n_99_29), .C2 (n_100_29) );
AOI211_X1 g_101_31 (.ZN (n_101_31), .A (n_105_29), .B (n_105_26), .C1 (n_101_28), .C2 (n_102_28) );
AOI211_X1 g_102_29 (.ZN (n_102_29), .A (n_103_30), .B (n_104_28), .C1 (n_103_27), .C2 (n_101_30) );
AOI211_X1 g_100_30 (.ZN (n_100_30), .A (n_101_31), .B (n_106_27), .C1 (n_105_26), .C2 (n_99_29) );
AOI211_X1 g_98_31 (.ZN (n_98_31), .A (n_102_29), .B (n_105_29), .C1 (n_104_28), .C2 (n_101_28) );
AOI211_X1 g_96_32 (.ZN (n_96_32), .A (n_100_30), .B (n_103_30), .C1 (n_106_27), .C2 (n_103_27) );
AOI211_X1 g_97_30 (.ZN (n_97_30), .A (n_98_31), .B (n_101_31), .C1 (n_105_29), .C2 (n_105_26) );
AOI211_X1 g_95_31 (.ZN (n_95_31), .A (n_96_32), .B (n_102_29), .C1 (n_103_30), .C2 (n_104_28) );
AOI211_X1 g_93_32 (.ZN (n_93_32), .A (n_97_30), .B (n_100_30), .C1 (n_101_31), .C2 (n_106_27) );
AOI211_X1 g_91_33 (.ZN (n_91_33), .A (n_95_31), .B (n_98_31), .C1 (n_102_29), .C2 (n_105_29) );
AOI211_X1 g_92_35 (.ZN (n_92_35), .A (n_93_32), .B (n_96_32), .C1 (n_100_30), .C2 (n_103_30) );
AOI211_X1 g_94_34 (.ZN (n_94_34), .A (n_91_33), .B (n_97_30), .C1 (n_98_31), .C2 (n_101_31) );
AOI211_X1 g_96_33 (.ZN (n_96_33), .A (n_92_35), .B (n_95_31), .C1 (n_96_32), .C2 (n_102_29) );
AOI211_X1 g_98_32 (.ZN (n_98_32), .A (n_94_34), .B (n_93_32), .C1 (n_97_30), .C2 (n_100_30) );
AOI211_X1 g_100_31 (.ZN (n_100_31), .A (n_96_33), .B (n_91_33), .C1 (n_95_31), .C2 (n_98_31) );
AOI211_X1 g_102_30 (.ZN (n_102_30), .A (n_98_32), .B (n_92_35), .C1 (n_93_32), .C2 (n_96_32) );
AOI211_X1 g_104_29 (.ZN (n_104_29), .A (n_100_31), .B (n_94_34), .C1 (n_91_33), .C2 (n_97_30) );
AOI211_X1 g_105_27 (.ZN (n_105_27), .A (n_102_30), .B (n_96_33), .C1 (n_92_35), .C2 (n_95_31) );
AOI211_X1 g_107_26 (.ZN (n_107_26), .A (n_104_29), .B (n_98_32), .C1 (n_94_34), .C2 (n_93_32) );
AOI211_X1 g_109_25 (.ZN (n_109_25), .A (n_105_27), .B (n_100_31), .C1 (n_96_33), .C2 (n_91_33) );
AOI211_X1 g_111_24 (.ZN (n_111_24), .A (n_107_26), .B (n_102_30), .C1 (n_98_32), .C2 (n_92_35) );
AOI211_X1 g_113_23 (.ZN (n_113_23), .A (n_109_25), .B (n_104_29), .C1 (n_100_31), .C2 (n_94_34) );
AOI211_X1 g_115_22 (.ZN (n_115_22), .A (n_111_24), .B (n_105_27), .C1 (n_102_30), .C2 (n_96_33) );
AOI211_X1 g_114_24 (.ZN (n_114_24), .A (n_113_23), .B (n_107_26), .C1 (n_104_29), .C2 (n_98_32) );
AOI211_X1 g_116_23 (.ZN (n_116_23), .A (n_115_22), .B (n_109_25), .C1 (n_105_27), .C2 (n_100_31) );
AOI211_X1 g_118_22 (.ZN (n_118_22), .A (n_114_24), .B (n_111_24), .C1 (n_107_26), .C2 (n_102_30) );
AOI211_X1 g_117_24 (.ZN (n_117_24), .A (n_116_23), .B (n_113_23), .C1 (n_109_25), .C2 (n_104_29) );
AOI211_X1 g_115_23 (.ZN (n_115_23), .A (n_118_22), .B (n_115_22), .C1 (n_111_24), .C2 (n_105_27) );
AOI211_X1 g_117_22 (.ZN (n_117_22), .A (n_117_24), .B (n_114_24), .C1 (n_113_23), .C2 (n_107_26) );
AOI211_X1 g_119_21 (.ZN (n_119_21), .A (n_115_23), .B (n_116_23), .C1 (n_115_22), .C2 (n_109_25) );
AOI211_X1 g_121_20 (.ZN (n_121_20), .A (n_117_22), .B (n_118_22), .C1 (n_114_24), .C2 (n_111_24) );
AOI211_X1 g_123_19 (.ZN (n_123_19), .A (n_119_21), .B (n_117_24), .C1 (n_116_23), .C2 (n_113_23) );
AOI211_X1 g_125_18 (.ZN (n_125_18), .A (n_121_20), .B (n_115_23), .C1 (n_118_22), .C2 (n_115_22) );
AOI211_X1 g_127_17 (.ZN (n_127_17), .A (n_123_19), .B (n_117_22), .C1 (n_117_24), .C2 (n_114_24) );
AOI211_X1 g_129_18 (.ZN (n_129_18), .A (n_125_18), .B (n_119_21), .C1 (n_115_23), .C2 (n_116_23) );
AOI211_X1 g_127_19 (.ZN (n_127_19), .A (n_127_17), .B (n_121_20), .C1 (n_117_22), .C2 (n_118_22) );
AOI211_X1 g_125_20 (.ZN (n_125_20), .A (n_129_18), .B (n_123_19), .C1 (n_119_21), .C2 (n_117_24) );
AOI211_X1 g_123_21 (.ZN (n_123_21), .A (n_127_19), .B (n_125_18), .C1 (n_121_20), .C2 (n_115_23) );
AOI211_X1 g_121_22 (.ZN (n_121_22), .A (n_125_20), .B (n_127_17), .C1 (n_123_19), .C2 (n_117_22) );
AOI211_X1 g_119_23 (.ZN (n_119_23), .A (n_123_21), .B (n_129_18), .C1 (n_125_18), .C2 (n_119_21) );
AOI211_X1 g_118_25 (.ZN (n_118_25), .A (n_121_22), .B (n_127_19), .C1 (n_127_17), .C2 (n_121_20) );
AOI211_X1 g_117_23 (.ZN (n_117_23), .A (n_119_23), .B (n_125_20), .C1 (n_129_18), .C2 (n_123_19) );
AOI211_X1 g_119_22 (.ZN (n_119_22), .A (n_118_25), .B (n_123_21), .C1 (n_127_19), .C2 (n_125_18) );
AOI211_X1 g_121_21 (.ZN (n_121_21), .A (n_117_23), .B (n_121_22), .C1 (n_125_20), .C2 (n_127_17) );
AOI211_X1 g_123_20 (.ZN (n_123_20), .A (n_119_22), .B (n_119_23), .C1 (n_123_21), .C2 (n_129_18) );
AOI211_X1 g_125_19 (.ZN (n_125_19), .A (n_121_21), .B (n_118_25), .C1 (n_121_22), .C2 (n_127_19) );
AOI211_X1 g_124_21 (.ZN (n_124_21), .A (n_123_20), .B (n_117_23), .C1 (n_119_23), .C2 (n_125_20) );
AOI211_X1 g_126_20 (.ZN (n_126_20), .A (n_125_19), .B (n_119_22), .C1 (n_118_25), .C2 (n_123_21) );
AOI211_X1 g_128_19 (.ZN (n_128_19), .A (n_124_21), .B (n_121_21), .C1 (n_117_23), .C2 (n_121_22) );
AOI211_X1 g_130_18 (.ZN (n_130_18), .A (n_126_20), .B (n_123_20), .C1 (n_119_22), .C2 (n_119_23) );
AOI211_X1 g_129_20 (.ZN (n_129_20), .A (n_128_19), .B (n_125_19), .C1 (n_121_21), .C2 (n_118_25) );
AOI211_X1 g_128_18 (.ZN (n_128_18), .A (n_130_18), .B (n_124_21), .C1 (n_123_20), .C2 (n_117_23) );
AOI211_X1 g_130_17 (.ZN (n_130_17), .A (n_129_20), .B (n_126_20), .C1 (n_125_19), .C2 (n_119_22) );
AOI211_X1 g_132_16 (.ZN (n_132_16), .A (n_128_18), .B (n_128_19), .C1 (n_124_21), .C2 (n_121_21) );
AOI211_X1 g_134_15 (.ZN (n_134_15), .A (n_130_17), .B (n_130_18), .C1 (n_126_20), .C2 (n_123_20) );
AOI211_X1 g_135_17 (.ZN (n_135_17), .A (n_132_16), .B (n_129_20), .C1 (n_128_19), .C2 (n_125_19) );
AOI211_X1 g_133_18 (.ZN (n_133_18), .A (n_134_15), .B (n_128_18), .C1 (n_130_18), .C2 (n_124_21) );
AOI211_X1 g_131_19 (.ZN (n_131_19), .A (n_135_17), .B (n_130_17), .C1 (n_129_20), .C2 (n_126_20) );
AOI211_X1 g_130_21 (.ZN (n_130_21), .A (n_133_18), .B (n_132_16), .C1 (n_128_18), .C2 (n_128_19) );
AOI211_X1 g_129_19 (.ZN (n_129_19), .A (n_131_19), .B (n_134_15), .C1 (n_130_17), .C2 (n_130_18) );
AOI211_X1 g_131_18 (.ZN (n_131_18), .A (n_130_21), .B (n_135_17), .C1 (n_132_16), .C2 (n_129_20) );
AOI211_X1 g_133_17 (.ZN (n_133_17), .A (n_129_19), .B (n_133_18), .C1 (n_134_15), .C2 (n_128_18) );
AOI211_X1 g_135_16 (.ZN (n_135_16), .A (n_131_18), .B (n_131_19), .C1 (n_135_17), .C2 (n_130_17) );
AOI211_X1 g_137_15 (.ZN (n_137_15), .A (n_133_17), .B (n_130_21), .C1 (n_133_18), .C2 (n_132_16) );
AOI211_X1 g_139_16 (.ZN (n_139_16), .A (n_135_16), .B (n_129_19), .C1 (n_131_19), .C2 (n_134_15) );
AOI211_X1 g_137_17 (.ZN (n_137_17), .A (n_137_15), .B (n_131_18), .C1 (n_130_21), .C2 (n_135_17) );
AOI211_X1 g_139_18 (.ZN (n_139_18), .A (n_139_16), .B (n_133_17), .C1 (n_129_19), .C2 (n_133_18) );
AOI211_X1 g_141_19 (.ZN (n_141_19), .A (n_137_17), .B (n_135_16), .C1 (n_131_18), .C2 (n_131_19) );
AOI211_X1 g_142_17 (.ZN (n_142_17), .A (n_139_18), .B (n_137_15), .C1 (n_133_17), .C2 (n_130_21) );
AOI211_X1 g_143_19 (.ZN (n_143_19), .A (n_141_19), .B (n_139_16), .C1 (n_135_16), .C2 (n_129_19) );
AOI211_X1 g_141_20 (.ZN (n_141_20), .A (n_142_17), .B (n_137_17), .C1 (n_137_15), .C2 (n_131_18) );
AOI211_X1 g_140_18 (.ZN (n_140_18), .A (n_143_19), .B (n_139_18), .C1 (n_139_16), .C2 (n_133_17) );
AOI211_X1 g_138_17 (.ZN (n_138_17), .A (n_141_20), .B (n_141_19), .C1 (n_137_17), .C2 (n_135_16) );
AOI211_X1 g_136_16 (.ZN (n_136_16), .A (n_140_18), .B (n_142_17), .C1 (n_139_18), .C2 (n_137_15) );
AOI211_X1 g_134_17 (.ZN (n_134_17), .A (n_138_17), .B (n_143_19), .C1 (n_141_19), .C2 (n_139_16) );
AOI211_X1 g_132_18 (.ZN (n_132_18), .A (n_136_16), .B (n_141_20), .C1 (n_142_17), .C2 (n_137_17) );
AOI211_X1 g_130_19 (.ZN (n_130_19), .A (n_134_17), .B (n_140_18), .C1 (n_143_19), .C2 (n_139_18) );
AOI211_X1 g_128_20 (.ZN (n_128_20), .A (n_132_18), .B (n_138_17), .C1 (n_141_20), .C2 (n_141_19) );
AOI211_X1 g_126_19 (.ZN (n_126_19), .A (n_130_19), .B (n_136_16), .C1 (n_140_18), .C2 (n_142_17) );
AOI211_X1 g_124_20 (.ZN (n_124_20), .A (n_128_20), .B (n_134_17), .C1 (n_138_17), .C2 (n_143_19) );
AOI211_X1 g_122_21 (.ZN (n_122_21), .A (n_126_19), .B (n_132_18), .C1 (n_136_16), .C2 (n_141_20) );
AOI211_X1 g_120_22 (.ZN (n_120_22), .A (n_124_20), .B (n_130_19), .C1 (n_134_17), .C2 (n_140_18) );
AOI211_X1 g_118_23 (.ZN (n_118_23), .A (n_122_21), .B (n_128_20), .C1 (n_132_18), .C2 (n_138_17) );
AOI211_X1 g_116_24 (.ZN (n_116_24), .A (n_120_22), .B (n_126_19), .C1 (n_130_19), .C2 (n_136_16) );
AOI211_X1 g_114_25 (.ZN (n_114_25), .A (n_118_23), .B (n_124_20), .C1 (n_128_20), .C2 (n_134_17) );
AOI211_X1 g_112_26 (.ZN (n_112_26), .A (n_116_24), .B (n_122_21), .C1 (n_126_19), .C2 (n_132_18) );
AOI211_X1 g_113_24 (.ZN (n_113_24), .A (n_114_25), .B (n_120_22), .C1 (n_124_20), .C2 (n_130_19) );
AOI211_X1 g_111_25 (.ZN (n_111_25), .A (n_112_26), .B (n_118_23), .C1 (n_122_21), .C2 (n_128_20) );
AOI211_X1 g_109_26 (.ZN (n_109_26), .A (n_113_24), .B (n_116_24), .C1 (n_120_22), .C2 (n_126_19) );
AOI211_X1 g_107_27 (.ZN (n_107_27), .A (n_111_25), .B (n_114_25), .C1 (n_118_23), .C2 (n_124_20) );
AOI211_X1 g_105_28 (.ZN (n_105_28), .A (n_109_26), .B (n_112_26), .C1 (n_116_24), .C2 (n_122_21) );
AOI211_X1 g_103_29 (.ZN (n_103_29), .A (n_107_27), .B (n_113_24), .C1 (n_114_25), .C2 (n_120_22) );
AOI211_X1 g_102_31 (.ZN (n_102_31), .A (n_105_28), .B (n_111_25), .C1 (n_112_26), .C2 (n_118_23) );
AOI211_X1 g_104_30 (.ZN (n_104_30), .A (n_103_29), .B (n_109_26), .C1 (n_113_24), .C2 (n_116_24) );
AOI211_X1 g_106_29 (.ZN (n_106_29), .A (n_102_31), .B (n_107_27), .C1 (n_111_25), .C2 (n_114_25) );
AOI211_X1 g_108_28 (.ZN (n_108_28), .A (n_104_30), .B (n_105_28), .C1 (n_109_26), .C2 (n_112_26) );
AOI211_X1 g_110_27 (.ZN (n_110_27), .A (n_106_29), .B (n_103_29), .C1 (n_107_27), .C2 (n_113_24) );
AOI211_X1 g_109_29 (.ZN (n_109_29), .A (n_108_28), .B (n_102_31), .C1 (n_105_28), .C2 (n_111_25) );
AOI211_X1 g_107_28 (.ZN (n_107_28), .A (n_110_27), .B (n_104_30), .C1 (n_103_29), .C2 (n_109_26) );
AOI211_X1 g_109_27 (.ZN (n_109_27), .A (n_109_29), .B (n_106_29), .C1 (n_102_31), .C2 (n_107_27) );
AOI211_X1 g_111_26 (.ZN (n_111_26), .A (n_107_28), .B (n_108_28), .C1 (n_104_30), .C2 (n_105_28) );
AOI211_X1 g_113_25 (.ZN (n_113_25), .A (n_109_27), .B (n_110_27), .C1 (n_106_29), .C2 (n_103_29) );
AOI211_X1 g_115_24 (.ZN (n_115_24), .A (n_111_26), .B (n_109_29), .C1 (n_108_28), .C2 (n_102_31) );
AOI211_X1 g_116_26 (.ZN (n_116_26), .A (n_113_25), .B (n_107_28), .C1 (n_110_27), .C2 (n_104_30) );
AOI211_X1 g_114_27 (.ZN (n_114_27), .A (n_115_24), .B (n_109_27), .C1 (n_109_29), .C2 (n_106_29) );
AOI211_X1 g_115_25 (.ZN (n_115_25), .A (n_116_26), .B (n_111_26), .C1 (n_107_28), .C2 (n_108_28) );
AOI211_X1 g_113_26 (.ZN (n_113_26), .A (n_114_27), .B (n_113_25), .C1 (n_109_27), .C2 (n_110_27) );
AOI211_X1 g_112_28 (.ZN (n_112_28), .A (n_115_25), .B (n_115_24), .C1 (n_111_26), .C2 (n_109_29) );
AOI211_X1 g_110_29 (.ZN (n_110_29), .A (n_113_26), .B (n_116_26), .C1 (n_113_25), .C2 (n_107_28) );
AOI211_X1 g_111_27 (.ZN (n_111_27), .A (n_112_28), .B (n_114_27), .C1 (n_115_24), .C2 (n_109_27) );
AOI211_X1 g_112_25 (.ZN (n_112_25), .A (n_110_29), .B (n_115_25), .C1 (n_116_26), .C2 (n_111_26) );
AOI211_X1 g_110_26 (.ZN (n_110_26), .A (n_111_27), .B (n_113_26), .C1 (n_114_27), .C2 (n_113_25) );
AOI211_X1 g_108_27 (.ZN (n_108_27), .A (n_112_25), .B (n_112_28), .C1 (n_115_25), .C2 (n_115_24) );
AOI211_X1 g_106_28 (.ZN (n_106_28), .A (n_110_26), .B (n_110_29), .C1 (n_113_26), .C2 (n_116_26) );
AOI211_X1 g_107_30 (.ZN (n_107_30), .A (n_108_27), .B (n_111_27), .C1 (n_112_28), .C2 (n_114_27) );
AOI211_X1 g_105_31 (.ZN (n_105_31), .A (n_106_28), .B (n_112_25), .C1 (n_110_29), .C2 (n_115_25) );
AOI211_X1 g_103_32 (.ZN (n_103_32), .A (n_107_30), .B (n_110_26), .C1 (n_111_27), .C2 (n_113_26) );
AOI211_X1 g_101_33 (.ZN (n_101_33), .A (n_105_31), .B (n_108_27), .C1 (n_112_25), .C2 (n_112_28) );
AOI211_X1 g_99_32 (.ZN (n_99_32), .A (n_103_32), .B (n_106_28), .C1 (n_110_26), .C2 (n_110_29) );
AOI211_X1 g_97_33 (.ZN (n_97_33), .A (n_101_33), .B (n_107_30), .C1 (n_108_27), .C2 (n_111_27) );
AOI211_X1 g_95_34 (.ZN (n_95_34), .A (n_99_32), .B (n_105_31), .C1 (n_106_28), .C2 (n_112_25) );
AOI211_X1 g_93_35 (.ZN (n_93_35), .A (n_97_33), .B (n_103_32), .C1 (n_107_30), .C2 (n_110_26) );
AOI211_X1 g_94_33 (.ZN (n_94_33), .A (n_95_34), .B (n_101_33), .C1 (n_105_31), .C2 (n_108_27) );
AOI211_X1 g_92_34 (.ZN (n_92_34), .A (n_93_35), .B (n_99_32), .C1 (n_103_32), .C2 (n_106_28) );
AOI211_X1 g_90_35 (.ZN (n_90_35), .A (n_94_33), .B (n_97_33), .C1 (n_101_33), .C2 (n_107_30) );
AOI211_X1 g_88_36 (.ZN (n_88_36), .A (n_92_34), .B (n_95_34), .C1 (n_99_32), .C2 (n_105_31) );
AOI211_X1 g_86_37 (.ZN (n_86_37), .A (n_90_35), .B (n_93_35), .C1 (n_97_33), .C2 (n_103_32) );
AOI211_X1 g_84_38 (.ZN (n_84_38), .A (n_88_36), .B (n_94_33), .C1 (n_95_34), .C2 (n_101_33) );
AOI211_X1 g_82_39 (.ZN (n_82_39), .A (n_86_37), .B (n_92_34), .C1 (n_93_35), .C2 (n_99_32) );
AOI211_X1 g_80_40 (.ZN (n_80_40), .A (n_84_38), .B (n_90_35), .C1 (n_94_33), .C2 (n_97_33) );
AOI211_X1 g_78_41 (.ZN (n_78_41), .A (n_82_39), .B (n_88_36), .C1 (n_92_34), .C2 (n_95_34) );
AOI211_X1 g_76_42 (.ZN (n_76_42), .A (n_80_40), .B (n_86_37), .C1 (n_90_35), .C2 (n_93_35) );
AOI211_X1 g_74_43 (.ZN (n_74_43), .A (n_78_41), .B (n_84_38), .C1 (n_88_36), .C2 (n_94_33) );
AOI211_X1 g_72_44 (.ZN (n_72_44), .A (n_76_42), .B (n_82_39), .C1 (n_86_37), .C2 (n_92_34) );
AOI211_X1 g_70_45 (.ZN (n_70_45), .A (n_74_43), .B (n_80_40), .C1 (n_84_38), .C2 (n_90_35) );
AOI211_X1 g_68_46 (.ZN (n_68_46), .A (n_72_44), .B (n_78_41), .C1 (n_82_39), .C2 (n_88_36) );
AOI211_X1 g_66_47 (.ZN (n_66_47), .A (n_70_45), .B (n_76_42), .C1 (n_80_40), .C2 (n_86_37) );
AOI211_X1 g_64_48 (.ZN (n_64_48), .A (n_68_46), .B (n_74_43), .C1 (n_78_41), .C2 (n_84_38) );
AOI211_X1 g_65_46 (.ZN (n_65_46), .A (n_66_47), .B (n_72_44), .C1 (n_76_42), .C2 (n_82_39) );
AOI211_X1 g_63_47 (.ZN (n_63_47), .A (n_64_48), .B (n_70_45), .C1 (n_74_43), .C2 (n_80_40) );
AOI211_X1 g_61_48 (.ZN (n_61_48), .A (n_65_46), .B (n_68_46), .C1 (n_72_44), .C2 (n_78_41) );
AOI211_X1 g_59_49 (.ZN (n_59_49), .A (n_63_47), .B (n_66_47), .C1 (n_70_45), .C2 (n_76_42) );
AOI211_X1 g_57_50 (.ZN (n_57_50), .A (n_61_48), .B (n_64_48), .C1 (n_68_46), .C2 (n_74_43) );
AOI211_X1 g_55_51 (.ZN (n_55_51), .A (n_59_49), .B (n_65_46), .C1 (n_66_47), .C2 (n_72_44) );
AOI211_X1 g_56_49 (.ZN (n_56_49), .A (n_57_50), .B (n_63_47), .C1 (n_64_48), .C2 (n_70_45) );
AOI211_X1 g_54_50 (.ZN (n_54_50), .A (n_55_51), .B (n_61_48), .C1 (n_65_46), .C2 (n_68_46) );
AOI211_X1 g_52_51 (.ZN (n_52_51), .A (n_56_49), .B (n_59_49), .C1 (n_63_47), .C2 (n_66_47) );
AOI211_X1 g_50_52 (.ZN (n_50_52), .A (n_54_50), .B (n_57_50), .C1 (n_61_48), .C2 (n_64_48) );
AOI211_X1 g_48_53 (.ZN (n_48_53), .A (n_52_51), .B (n_55_51), .C1 (n_59_49), .C2 (n_65_46) );
AOI211_X1 g_46_54 (.ZN (n_46_54), .A (n_50_52), .B (n_56_49), .C1 (n_57_50), .C2 (n_63_47) );
AOI211_X1 g_44_55 (.ZN (n_44_55), .A (n_48_53), .B (n_54_50), .C1 (n_55_51), .C2 (n_61_48) );
AOI211_X1 g_42_56 (.ZN (n_42_56), .A (n_46_54), .B (n_52_51), .C1 (n_56_49), .C2 (n_59_49) );
AOI211_X1 g_40_57 (.ZN (n_40_57), .A (n_44_55), .B (n_50_52), .C1 (n_54_50), .C2 (n_57_50) );
AOI211_X1 g_38_58 (.ZN (n_38_58), .A (n_42_56), .B (n_48_53), .C1 (n_52_51), .C2 (n_55_51) );
AOI211_X1 g_36_59 (.ZN (n_36_59), .A (n_40_57), .B (n_46_54), .C1 (n_50_52), .C2 (n_56_49) );
AOI211_X1 g_34_60 (.ZN (n_34_60), .A (n_38_58), .B (n_44_55), .C1 (n_48_53), .C2 (n_54_50) );
AOI211_X1 g_32_61 (.ZN (n_32_61), .A (n_36_59), .B (n_42_56), .C1 (n_46_54), .C2 (n_52_51) );
AOI211_X1 g_30_62 (.ZN (n_30_62), .A (n_34_60), .B (n_40_57), .C1 (n_44_55), .C2 (n_50_52) );
AOI211_X1 g_28_63 (.ZN (n_28_63), .A (n_32_61), .B (n_38_58), .C1 (n_42_56), .C2 (n_48_53) );
AOI211_X1 g_26_64 (.ZN (n_26_64), .A (n_30_62), .B (n_36_59), .C1 (n_40_57), .C2 (n_46_54) );
AOI211_X1 g_24_65 (.ZN (n_24_65), .A (n_28_63), .B (n_34_60), .C1 (n_38_58), .C2 (n_44_55) );
AOI211_X1 g_22_66 (.ZN (n_22_66), .A (n_26_64), .B (n_32_61), .C1 (n_36_59), .C2 (n_42_56) );
AOI211_X1 g_20_67 (.ZN (n_20_67), .A (n_24_65), .B (n_30_62), .C1 (n_34_60), .C2 (n_40_57) );
AOI211_X1 g_18_68 (.ZN (n_18_68), .A (n_22_66), .B (n_28_63), .C1 (n_32_61), .C2 (n_38_58) );
AOI211_X1 g_16_69 (.ZN (n_16_69), .A (n_20_67), .B (n_26_64), .C1 (n_30_62), .C2 (n_36_59) );
AOI211_X1 g_14_70 (.ZN (n_14_70), .A (n_18_68), .B (n_24_65), .C1 (n_28_63), .C2 (n_34_60) );
AOI211_X1 g_12_71 (.ZN (n_12_71), .A (n_16_69), .B (n_22_66), .C1 (n_26_64), .C2 (n_32_61) );
AOI211_X1 g_10_72 (.ZN (n_10_72), .A (n_14_70), .B (n_20_67), .C1 (n_24_65), .C2 (n_30_62) );
AOI211_X1 g_8_73 (.ZN (n_8_73), .A (n_12_71), .B (n_18_68), .C1 (n_22_66), .C2 (n_28_63) );
AOI211_X1 g_6_74 (.ZN (n_6_74), .A (n_10_72), .B (n_16_69), .C1 (n_20_67), .C2 (n_26_64) );
AOI211_X1 g_4_75 (.ZN (n_4_75), .A (n_8_73), .B (n_14_70), .C1 (n_18_68), .C2 (n_24_65) );
AOI211_X1 g_3_77 (.ZN (n_3_77), .A (n_6_74), .B (n_12_71), .C1 (n_16_69), .C2 (n_22_66) );
AOI211_X1 g_5_76 (.ZN (n_5_76), .A (n_4_75), .B (n_10_72), .C1 (n_14_70), .C2 (n_20_67) );
AOI211_X1 g_4_74 (.ZN (n_4_74), .A (n_3_77), .B (n_8_73), .C1 (n_12_71), .C2 (n_18_68) );
AOI211_X1 g_6_73 (.ZN (n_6_73), .A (n_5_76), .B (n_6_74), .C1 (n_10_72), .C2 (n_16_69) );
AOI211_X1 g_8_72 (.ZN (n_8_72), .A (n_4_74), .B (n_4_75), .C1 (n_8_73), .C2 (n_14_70) );
AOI211_X1 g_10_71 (.ZN (n_10_71), .A (n_6_73), .B (n_3_77), .C1 (n_6_74), .C2 (n_12_71) );
AOI211_X1 g_12_70 (.ZN (n_12_70), .A (n_8_72), .B (n_5_76), .C1 (n_4_75), .C2 (n_10_72) );
AOI211_X1 g_14_69 (.ZN (n_14_69), .A (n_10_71), .B (n_4_74), .C1 (n_3_77), .C2 (n_8_73) );
AOI211_X1 g_13_71 (.ZN (n_13_71), .A (n_12_70), .B (n_6_73), .C1 (n_5_76), .C2 (n_6_74) );
AOI211_X1 g_15_70 (.ZN (n_15_70), .A (n_14_69), .B (n_8_72), .C1 (n_4_74), .C2 (n_4_75) );
AOI211_X1 g_14_72 (.ZN (n_14_72), .A (n_13_71), .B (n_10_71), .C1 (n_6_73), .C2 (n_3_77) );
AOI211_X1 g_16_71 (.ZN (n_16_71), .A (n_15_70), .B (n_12_70), .C1 (n_8_72), .C2 (n_5_76) );
AOI211_X1 g_18_70 (.ZN (n_18_70), .A (n_14_72), .B (n_14_69), .C1 (n_10_71), .C2 (n_4_74) );
AOI211_X1 g_20_69 (.ZN (n_20_69), .A (n_16_71), .B (n_13_71), .C1 (n_12_70), .C2 (n_6_73) );
AOI211_X1 g_22_68 (.ZN (n_22_68), .A (n_18_70), .B (n_15_70), .C1 (n_14_69), .C2 (n_8_72) );
AOI211_X1 g_23_66 (.ZN (n_23_66), .A (n_20_69), .B (n_14_72), .C1 (n_13_71), .C2 (n_10_71) );
AOI211_X1 g_25_65 (.ZN (n_25_65), .A (n_22_68), .B (n_16_71), .C1 (n_15_70), .C2 (n_12_70) );
AOI211_X1 g_27_64 (.ZN (n_27_64), .A (n_23_66), .B (n_18_70), .C1 (n_14_72), .C2 (n_14_69) );
AOI211_X1 g_29_63 (.ZN (n_29_63), .A (n_25_65), .B (n_20_69), .C1 (n_16_71), .C2 (n_13_71) );
AOI211_X1 g_31_62 (.ZN (n_31_62), .A (n_27_64), .B (n_22_68), .C1 (n_18_70), .C2 (n_15_70) );
AOI211_X1 g_33_61 (.ZN (n_33_61), .A (n_29_63), .B (n_23_66), .C1 (n_20_69), .C2 (n_14_72) );
AOI211_X1 g_35_60 (.ZN (n_35_60), .A (n_31_62), .B (n_25_65), .C1 (n_22_68), .C2 (n_16_71) );
AOI211_X1 g_37_59 (.ZN (n_37_59), .A (n_33_61), .B (n_27_64), .C1 (n_23_66), .C2 (n_18_70) );
AOI211_X1 g_39_58 (.ZN (n_39_58), .A (n_35_60), .B (n_29_63), .C1 (n_25_65), .C2 (n_20_69) );
AOI211_X1 g_38_60 (.ZN (n_38_60), .A (n_37_59), .B (n_31_62), .C1 (n_27_64), .C2 (n_22_68) );
AOI211_X1 g_40_59 (.ZN (n_40_59), .A (n_39_58), .B (n_33_61), .C1 (n_29_63), .C2 (n_23_66) );
AOI211_X1 g_42_58 (.ZN (n_42_58), .A (n_38_60), .B (n_35_60), .C1 (n_31_62), .C2 (n_25_65) );
AOI211_X1 g_44_57 (.ZN (n_44_57), .A (n_40_59), .B (n_37_59), .C1 (n_33_61), .C2 (n_27_64) );
AOI211_X1 g_46_56 (.ZN (n_46_56), .A (n_42_58), .B (n_39_58), .C1 (n_35_60), .C2 (n_29_63) );
AOI211_X1 g_48_55 (.ZN (n_48_55), .A (n_44_57), .B (n_38_60), .C1 (n_37_59), .C2 (n_31_62) );
AOI211_X1 g_50_54 (.ZN (n_50_54), .A (n_46_56), .B (n_40_59), .C1 (n_39_58), .C2 (n_33_61) );
AOI211_X1 g_52_53 (.ZN (n_52_53), .A (n_48_55), .B (n_42_58), .C1 (n_38_60), .C2 (n_35_60) );
AOI211_X1 g_54_52 (.ZN (n_54_52), .A (n_50_54), .B (n_44_57), .C1 (n_40_59), .C2 (n_37_59) );
AOI211_X1 g_56_51 (.ZN (n_56_51), .A (n_52_53), .B (n_46_56), .C1 (n_42_58), .C2 (n_39_58) );
AOI211_X1 g_58_50 (.ZN (n_58_50), .A (n_54_52), .B (n_48_55), .C1 (n_44_57), .C2 (n_38_60) );
AOI211_X1 g_60_49 (.ZN (n_60_49), .A (n_56_51), .B (n_50_54), .C1 (n_46_56), .C2 (n_40_59) );
AOI211_X1 g_62_48 (.ZN (n_62_48), .A (n_58_50), .B (n_52_53), .C1 (n_48_55), .C2 (n_42_58) );
AOI211_X1 g_64_47 (.ZN (n_64_47), .A (n_60_49), .B (n_54_52), .C1 (n_50_54), .C2 (n_44_57) );
AOI211_X1 g_66_46 (.ZN (n_66_46), .A (n_62_48), .B (n_56_51), .C1 (n_52_53), .C2 (n_46_56) );
AOI211_X1 g_68_45 (.ZN (n_68_45), .A (n_64_47), .B (n_58_50), .C1 (n_54_52), .C2 (n_48_55) );
AOI211_X1 g_70_44 (.ZN (n_70_44), .A (n_66_46), .B (n_60_49), .C1 (n_56_51), .C2 (n_50_54) );
AOI211_X1 g_72_43 (.ZN (n_72_43), .A (n_68_45), .B (n_62_48), .C1 (n_58_50), .C2 (n_52_53) );
AOI211_X1 g_74_42 (.ZN (n_74_42), .A (n_70_44), .B (n_64_47), .C1 (n_60_49), .C2 (n_54_52) );
AOI211_X1 g_76_41 (.ZN (n_76_41), .A (n_72_43), .B (n_66_46), .C1 (n_62_48), .C2 (n_56_51) );
AOI211_X1 g_78_40 (.ZN (n_78_40), .A (n_74_42), .B (n_68_45), .C1 (n_64_47), .C2 (n_58_50) );
AOI211_X1 g_80_39 (.ZN (n_80_39), .A (n_76_41), .B (n_70_44), .C1 (n_66_46), .C2 (n_60_49) );
AOI211_X1 g_82_38 (.ZN (n_82_38), .A (n_78_40), .B (n_72_43), .C1 (n_68_45), .C2 (n_62_48) );
AOI211_X1 g_84_37 (.ZN (n_84_37), .A (n_80_39), .B (n_74_42), .C1 (n_70_44), .C2 (n_64_47) );
AOI211_X1 g_86_36 (.ZN (n_86_36), .A (n_82_38), .B (n_76_41), .C1 (n_72_43), .C2 (n_66_46) );
AOI211_X1 g_88_37 (.ZN (n_88_37), .A (n_84_37), .B (n_78_40), .C1 (n_74_42), .C2 (n_68_45) );
AOI211_X1 g_86_38 (.ZN (n_86_38), .A (n_86_36), .B (n_80_39), .C1 (n_76_41), .C2 (n_70_44) );
AOI211_X1 g_84_39 (.ZN (n_84_39), .A (n_88_37), .B (n_82_38), .C1 (n_78_40), .C2 (n_72_43) );
AOI211_X1 g_82_40 (.ZN (n_82_40), .A (n_86_38), .B (n_84_37), .C1 (n_80_39), .C2 (n_74_42) );
AOI211_X1 g_80_41 (.ZN (n_80_41), .A (n_84_39), .B (n_86_36), .C1 (n_82_38), .C2 (n_76_41) );
AOI211_X1 g_78_42 (.ZN (n_78_42), .A (n_82_40), .B (n_88_37), .C1 (n_84_37), .C2 (n_78_40) );
AOI211_X1 g_76_43 (.ZN (n_76_43), .A (n_80_41), .B (n_86_38), .C1 (n_86_36), .C2 (n_80_39) );
AOI211_X1 g_74_44 (.ZN (n_74_44), .A (n_78_42), .B (n_84_39), .C1 (n_88_37), .C2 (n_82_38) );
AOI211_X1 g_72_45 (.ZN (n_72_45), .A (n_76_43), .B (n_82_40), .C1 (n_86_38), .C2 (n_84_37) );
AOI211_X1 g_70_46 (.ZN (n_70_46), .A (n_74_44), .B (n_80_41), .C1 (n_84_39), .C2 (n_86_36) );
AOI211_X1 g_69_48 (.ZN (n_69_48), .A (n_72_45), .B (n_78_42), .C1 (n_82_40), .C2 (n_88_37) );
AOI211_X1 g_67_47 (.ZN (n_67_47), .A (n_70_46), .B (n_76_43), .C1 (n_80_41), .C2 (n_86_38) );
AOI211_X1 g_69_46 (.ZN (n_69_46), .A (n_69_48), .B (n_74_44), .C1 (n_78_42), .C2 (n_84_39) );
AOI211_X1 g_71_45 (.ZN (n_71_45), .A (n_67_47), .B (n_72_45), .C1 (n_76_43), .C2 (n_82_40) );
AOI211_X1 g_73_44 (.ZN (n_73_44), .A (n_69_46), .B (n_70_46), .C1 (n_74_44), .C2 (n_80_41) );
AOI211_X1 g_75_43 (.ZN (n_75_43), .A (n_71_45), .B (n_69_48), .C1 (n_72_45), .C2 (n_78_42) );
AOI211_X1 g_77_42 (.ZN (n_77_42), .A (n_73_44), .B (n_67_47), .C1 (n_70_46), .C2 (n_76_43) );
AOI211_X1 g_79_41 (.ZN (n_79_41), .A (n_75_43), .B (n_69_46), .C1 (n_69_48), .C2 (n_74_44) );
AOI211_X1 g_81_40 (.ZN (n_81_40), .A (n_77_42), .B (n_71_45), .C1 (n_67_47), .C2 (n_72_45) );
AOI211_X1 g_83_39 (.ZN (n_83_39), .A (n_79_41), .B (n_73_44), .C1 (n_69_46), .C2 (n_70_46) );
AOI211_X1 g_85_38 (.ZN (n_85_38), .A (n_81_40), .B (n_75_43), .C1 (n_71_45), .C2 (n_69_48) );
AOI211_X1 g_87_37 (.ZN (n_87_37), .A (n_83_39), .B (n_77_42), .C1 (n_73_44), .C2 (n_67_47) );
AOI211_X1 g_89_36 (.ZN (n_89_36), .A (n_85_38), .B (n_79_41), .C1 (n_75_43), .C2 (n_69_46) );
AOI211_X1 g_91_35 (.ZN (n_91_35), .A (n_87_37), .B (n_81_40), .C1 (n_77_42), .C2 (n_71_45) );
AOI211_X1 g_93_34 (.ZN (n_93_34), .A (n_89_36), .B (n_83_39), .C1 (n_79_41), .C2 (n_73_44) );
AOI211_X1 g_95_33 (.ZN (n_95_33), .A (n_91_35), .B (n_85_38), .C1 (n_81_40), .C2 (n_75_43) );
AOI211_X1 g_97_32 (.ZN (n_97_32), .A (n_93_34), .B (n_87_37), .C1 (n_83_39), .C2 (n_77_42) );
AOI211_X1 g_99_31 (.ZN (n_99_31), .A (n_95_33), .B (n_89_36), .C1 (n_85_38), .C2 (n_79_41) );
AOI211_X1 g_98_33 (.ZN (n_98_33), .A (n_97_32), .B (n_91_35), .C1 (n_87_37), .C2 (n_81_40) );
AOI211_X1 g_100_32 (.ZN (n_100_32), .A (n_99_31), .B (n_93_34), .C1 (n_89_36), .C2 (n_83_39) );
AOI211_X1 g_99_34 (.ZN (n_99_34), .A (n_98_33), .B (n_95_33), .C1 (n_91_35), .C2 (n_85_38) );
AOI211_X1 g_97_35 (.ZN (n_97_35), .A (n_100_32), .B (n_97_32), .C1 (n_93_34), .C2 (n_87_37) );
AOI211_X1 g_95_36 (.ZN (n_95_36), .A (n_99_34), .B (n_99_31), .C1 (n_95_33), .C2 (n_89_36) );
AOI211_X1 g_96_34 (.ZN (n_96_34), .A (n_97_35), .B (n_98_33), .C1 (n_97_32), .C2 (n_91_35) );
AOI211_X1 g_94_35 (.ZN (n_94_35), .A (n_95_36), .B (n_100_32), .C1 (n_99_31), .C2 (n_93_34) );
AOI211_X1 g_92_36 (.ZN (n_92_36), .A (n_96_34), .B (n_99_34), .C1 (n_98_33), .C2 (n_95_33) );
AOI211_X1 g_90_37 (.ZN (n_90_37), .A (n_94_35), .B (n_97_35), .C1 (n_100_32), .C2 (n_97_32) );
AOI211_X1 g_88_38 (.ZN (n_88_38), .A (n_92_36), .B (n_95_36), .C1 (n_99_34), .C2 (n_99_31) );
AOI211_X1 g_86_39 (.ZN (n_86_39), .A (n_90_37), .B (n_96_34), .C1 (n_97_35), .C2 (n_98_33) );
AOI211_X1 g_84_40 (.ZN (n_84_40), .A (n_88_38), .B (n_94_35), .C1 (n_95_36), .C2 (n_100_32) );
AOI211_X1 g_82_41 (.ZN (n_82_41), .A (n_86_39), .B (n_92_36), .C1 (n_96_34), .C2 (n_99_34) );
AOI211_X1 g_80_42 (.ZN (n_80_42), .A (n_84_40), .B (n_90_37), .C1 (n_94_35), .C2 (n_97_35) );
AOI211_X1 g_78_43 (.ZN (n_78_43), .A (n_82_41), .B (n_88_38), .C1 (n_92_36), .C2 (n_95_36) );
AOI211_X1 g_76_44 (.ZN (n_76_44), .A (n_80_42), .B (n_86_39), .C1 (n_90_37), .C2 (n_96_34) );
AOI211_X1 g_74_45 (.ZN (n_74_45), .A (n_78_43), .B (n_84_40), .C1 (n_88_38), .C2 (n_94_35) );
AOI211_X1 g_72_46 (.ZN (n_72_46), .A (n_76_44), .B (n_82_41), .C1 (n_86_39), .C2 (n_92_36) );
AOI211_X1 g_70_47 (.ZN (n_70_47), .A (n_74_45), .B (n_80_42), .C1 (n_84_40), .C2 (n_90_37) );
AOI211_X1 g_68_48 (.ZN (n_68_48), .A (n_72_46), .B (n_78_43), .C1 (n_82_41), .C2 (n_88_38) );
AOI211_X1 g_66_49 (.ZN (n_66_49), .A (n_70_47), .B (n_76_44), .C1 (n_80_42), .C2 (n_86_39) );
AOI211_X1 g_64_50 (.ZN (n_64_50), .A (n_68_48), .B (n_74_45), .C1 (n_78_43), .C2 (n_84_40) );
AOI211_X1 g_65_48 (.ZN (n_65_48), .A (n_66_49), .B (n_72_46), .C1 (n_76_44), .C2 (n_82_41) );
AOI211_X1 g_63_49 (.ZN (n_63_49), .A (n_64_50), .B (n_70_47), .C1 (n_74_45), .C2 (n_80_42) );
AOI211_X1 g_61_50 (.ZN (n_61_50), .A (n_65_48), .B (n_68_48), .C1 (n_72_46), .C2 (n_78_43) );
AOI211_X1 g_59_51 (.ZN (n_59_51), .A (n_63_49), .B (n_66_49), .C1 (n_70_47), .C2 (n_76_44) );
AOI211_X1 g_57_52 (.ZN (n_57_52), .A (n_61_50), .B (n_64_50), .C1 (n_68_48), .C2 (n_74_45) );
AOI211_X1 g_55_53 (.ZN (n_55_53), .A (n_59_51), .B (n_65_48), .C1 (n_66_49), .C2 (n_72_46) );
AOI211_X1 g_53_52 (.ZN (n_53_52), .A (n_57_52), .B (n_63_49), .C1 (n_64_50), .C2 (n_70_47) );
AOI211_X1 g_51_53 (.ZN (n_51_53), .A (n_55_53), .B (n_61_50), .C1 (n_65_48), .C2 (n_68_48) );
AOI211_X1 g_49_54 (.ZN (n_49_54), .A (n_53_52), .B (n_59_51), .C1 (n_63_49), .C2 (n_66_49) );
AOI211_X1 g_47_55 (.ZN (n_47_55), .A (n_51_53), .B (n_57_52), .C1 (n_61_50), .C2 (n_64_50) );
AOI211_X1 g_45_56 (.ZN (n_45_56), .A (n_49_54), .B (n_55_53), .C1 (n_59_51), .C2 (n_65_48) );
AOI211_X1 g_43_57 (.ZN (n_43_57), .A (n_47_55), .B (n_53_52), .C1 (n_57_52), .C2 (n_63_49) );
AOI211_X1 g_41_58 (.ZN (n_41_58), .A (n_45_56), .B (n_51_53), .C1 (n_55_53), .C2 (n_61_50) );
AOI211_X1 g_39_59 (.ZN (n_39_59), .A (n_43_57), .B (n_49_54), .C1 (n_53_52), .C2 (n_59_51) );
AOI211_X1 g_37_60 (.ZN (n_37_60), .A (n_41_58), .B (n_47_55), .C1 (n_51_53), .C2 (n_57_52) );
AOI211_X1 g_35_61 (.ZN (n_35_61), .A (n_39_59), .B (n_45_56), .C1 (n_49_54), .C2 (n_55_53) );
AOI211_X1 g_33_62 (.ZN (n_33_62), .A (n_37_60), .B (n_43_57), .C1 (n_47_55), .C2 (n_53_52) );
AOI211_X1 g_31_63 (.ZN (n_31_63), .A (n_35_61), .B (n_41_58), .C1 (n_45_56), .C2 (n_51_53) );
AOI211_X1 g_29_64 (.ZN (n_29_64), .A (n_33_62), .B (n_39_59), .C1 (n_43_57), .C2 (n_49_54) );
AOI211_X1 g_27_65 (.ZN (n_27_65), .A (n_31_63), .B (n_37_60), .C1 (n_41_58), .C2 (n_47_55) );
AOI211_X1 g_25_66 (.ZN (n_25_66), .A (n_29_64), .B (n_35_61), .C1 (n_39_59), .C2 (n_45_56) );
AOI211_X1 g_23_67 (.ZN (n_23_67), .A (n_27_65), .B (n_33_62), .C1 (n_37_60), .C2 (n_43_57) );
AOI211_X1 g_21_68 (.ZN (n_21_68), .A (n_25_66), .B (n_31_63), .C1 (n_35_61), .C2 (n_41_58) );
AOI211_X1 g_19_69 (.ZN (n_19_69), .A (n_23_67), .B (n_29_64), .C1 (n_33_62), .C2 (n_39_59) );
AOI211_X1 g_17_70 (.ZN (n_17_70), .A (n_21_68), .B (n_27_65), .C1 (n_31_63), .C2 (n_37_60) );
AOI211_X1 g_15_71 (.ZN (n_15_71), .A (n_19_69), .B (n_25_66), .C1 (n_29_64), .C2 (n_35_61) );
AOI211_X1 g_13_72 (.ZN (n_13_72), .A (n_17_70), .B (n_23_67), .C1 (n_27_65), .C2 (n_33_62) );
AOI211_X1 g_11_73 (.ZN (n_11_73), .A (n_15_71), .B (n_21_68), .C1 (n_25_66), .C2 (n_31_63) );
AOI211_X1 g_9_74 (.ZN (n_9_74), .A (n_13_72), .B (n_19_69), .C1 (n_23_67), .C2 (n_29_64) );
AOI211_X1 g_7_75 (.ZN (n_7_75), .A (n_11_73), .B (n_17_70), .C1 (n_21_68), .C2 (n_27_65) );
AOI211_X1 g_6_77 (.ZN (n_6_77), .A (n_9_74), .B (n_15_71), .C1 (n_19_69), .C2 (n_25_66) );
AOI211_X1 g_5_75 (.ZN (n_5_75), .A (n_7_75), .B (n_13_72), .C1 (n_17_70), .C2 (n_23_67) );
AOI211_X1 g_3_76 (.ZN (n_3_76), .A (n_6_77), .B (n_11_73), .C1 (n_15_71), .C2 (n_21_68) );
AOI211_X1 g_4_78 (.ZN (n_4_78), .A (n_5_75), .B (n_9_74), .C1 (n_13_72), .C2 (n_19_69) );
AOI211_X1 g_3_80 (.ZN (n_3_80), .A (n_3_76), .B (n_7_75), .C1 (n_11_73), .C2 (n_17_70) );
AOI211_X1 g_2_78 (.ZN (n_2_78), .A (n_4_78), .B (n_6_77), .C1 (n_9_74), .C2 (n_15_71) );
AOI211_X1 g_1_80 (.ZN (n_1_80), .A (n_3_80), .B (n_5_75), .C1 (n_7_75), .C2 (n_13_72) );
AOI211_X1 g_3_79 (.ZN (n_3_79), .A (n_2_78), .B (n_3_76), .C1 (n_6_77), .C2 (n_11_73) );
AOI211_X1 g_4_77 (.ZN (n_4_77), .A (n_1_80), .B (n_4_78), .C1 (n_5_75), .C2 (n_9_74) );
AOI211_X1 g_5_79 (.ZN (n_5_79), .A (n_3_79), .B (n_3_80), .C1 (n_3_76), .C2 (n_7_75) );
AOI211_X1 g_4_81 (.ZN (n_4_81), .A (n_4_77), .B (n_2_78), .C1 (n_4_78), .C2 (n_6_77) );
AOI211_X1 g_2_82 (.ZN (n_2_82), .A (n_5_79), .B (n_1_80), .C1 (n_3_80), .C2 (n_5_75) );
AOI211_X1 g_1_84 (.ZN (n_1_84), .A (n_4_81), .B (n_3_79), .C1 (n_2_78), .C2 (n_3_76) );
AOI211_X1 g_3_83 (.ZN (n_3_83), .A (n_2_82), .B (n_4_77), .C1 (n_1_80), .C2 (n_4_78) );
AOI211_X1 g_5_82 (.ZN (n_5_82), .A (n_1_84), .B (n_5_79), .C1 (n_3_79), .C2 (n_3_80) );
AOI211_X1 g_3_81 (.ZN (n_3_81), .A (n_3_83), .B (n_4_81), .C1 (n_4_77), .C2 (n_2_78) );
AOI211_X1 g_4_79 (.ZN (n_4_79), .A (n_5_82), .B (n_2_82), .C1 (n_5_79), .C2 (n_1_80) );
AOI211_X1 g_5_77 (.ZN (n_5_77), .A (n_3_81), .B (n_1_84), .C1 (n_4_81), .C2 (n_3_79) );
AOI211_X1 g_6_75 (.ZN (n_6_75), .A (n_4_79), .B (n_3_83), .C1 (n_2_82), .C2 (n_4_77) );
AOI211_X1 g_8_74 (.ZN (n_8_74), .A (n_5_77), .B (n_5_82), .C1 (n_1_84), .C2 (n_5_79) );
AOI211_X1 g_10_73 (.ZN (n_10_73), .A (n_6_75), .B (n_3_81), .C1 (n_3_83), .C2 (n_4_81) );
AOI211_X1 g_12_72 (.ZN (n_12_72), .A (n_8_74), .B (n_4_79), .C1 (n_5_82), .C2 (n_2_82) );
AOI211_X1 g_14_71 (.ZN (n_14_71), .A (n_10_73), .B (n_5_77), .C1 (n_3_81), .C2 (n_1_84) );
AOI211_X1 g_16_70 (.ZN (n_16_70), .A (n_12_72), .B (n_6_75), .C1 (n_4_79), .C2 (n_3_83) );
AOI211_X1 g_18_69 (.ZN (n_18_69), .A (n_14_71), .B (n_8_74), .C1 (n_5_77), .C2 (n_5_82) );
AOI211_X1 g_20_68 (.ZN (n_20_68), .A (n_16_70), .B (n_10_73), .C1 (n_6_75), .C2 (n_3_81) );
AOI211_X1 g_19_70 (.ZN (n_19_70), .A (n_18_69), .B (n_12_72), .C1 (n_8_74), .C2 (n_4_79) );
AOI211_X1 g_21_69 (.ZN (n_21_69), .A (n_20_68), .B (n_14_71), .C1 (n_10_73), .C2 (n_5_77) );
AOI211_X1 g_23_68 (.ZN (n_23_68), .A (n_19_70), .B (n_16_70), .C1 (n_12_72), .C2 (n_6_75) );
AOI211_X1 g_25_67 (.ZN (n_25_67), .A (n_21_69), .B (n_18_69), .C1 (n_14_71), .C2 (n_8_74) );
AOI211_X1 g_27_66 (.ZN (n_27_66), .A (n_23_68), .B (n_20_68), .C1 (n_16_70), .C2 (n_10_73) );
AOI211_X1 g_29_65 (.ZN (n_29_65), .A (n_25_67), .B (n_19_70), .C1 (n_18_69), .C2 (n_12_72) );
AOI211_X1 g_31_64 (.ZN (n_31_64), .A (n_27_66), .B (n_21_69), .C1 (n_20_68), .C2 (n_14_71) );
AOI211_X1 g_33_63 (.ZN (n_33_63), .A (n_29_65), .B (n_23_68), .C1 (n_19_70), .C2 (n_16_70) );
AOI211_X1 g_35_62 (.ZN (n_35_62), .A (n_31_64), .B (n_25_67), .C1 (n_21_69), .C2 (n_18_69) );
AOI211_X1 g_37_61 (.ZN (n_37_61), .A (n_33_63), .B (n_27_66), .C1 (n_23_68), .C2 (n_20_68) );
AOI211_X1 g_39_60 (.ZN (n_39_60), .A (n_35_62), .B (n_29_65), .C1 (n_25_67), .C2 (n_19_70) );
AOI211_X1 g_41_59 (.ZN (n_41_59), .A (n_37_61), .B (n_31_64), .C1 (n_27_66), .C2 (n_21_69) );
AOI211_X1 g_43_58 (.ZN (n_43_58), .A (n_39_60), .B (n_33_63), .C1 (n_29_65), .C2 (n_23_68) );
AOI211_X1 g_45_57 (.ZN (n_45_57), .A (n_41_59), .B (n_35_62), .C1 (n_31_64), .C2 (n_25_67) );
AOI211_X1 g_47_56 (.ZN (n_47_56), .A (n_43_58), .B (n_37_61), .C1 (n_33_63), .C2 (n_27_66) );
AOI211_X1 g_49_55 (.ZN (n_49_55), .A (n_45_57), .B (n_39_60), .C1 (n_35_62), .C2 (n_29_65) );
AOI211_X1 g_51_54 (.ZN (n_51_54), .A (n_47_56), .B (n_41_59), .C1 (n_37_61), .C2 (n_31_64) );
AOI211_X1 g_53_53 (.ZN (n_53_53), .A (n_49_55), .B (n_43_58), .C1 (n_39_60), .C2 (n_33_63) );
AOI211_X1 g_55_52 (.ZN (n_55_52), .A (n_51_54), .B (n_45_57), .C1 (n_41_59), .C2 (n_35_62) );
AOI211_X1 g_57_51 (.ZN (n_57_51), .A (n_53_53), .B (n_47_56), .C1 (n_43_58), .C2 (n_37_61) );
AOI211_X1 g_56_53 (.ZN (n_56_53), .A (n_55_52), .B (n_49_55), .C1 (n_45_57), .C2 (n_39_60) );
AOI211_X1 g_58_52 (.ZN (n_58_52), .A (n_57_51), .B (n_51_54), .C1 (n_47_56), .C2 (n_41_59) );
AOI211_X1 g_60_51 (.ZN (n_60_51), .A (n_56_53), .B (n_53_53), .C1 (n_49_55), .C2 (n_43_58) );
AOI211_X1 g_62_50 (.ZN (n_62_50), .A (n_58_52), .B (n_55_52), .C1 (n_51_54), .C2 (n_45_57) );
AOI211_X1 g_64_49 (.ZN (n_64_49), .A (n_60_51), .B (n_57_51), .C1 (n_53_53), .C2 (n_47_56) );
AOI211_X1 g_66_48 (.ZN (n_66_48), .A (n_62_50), .B (n_56_53), .C1 (n_55_52), .C2 (n_49_55) );
AOI211_X1 g_65_50 (.ZN (n_65_50), .A (n_64_49), .B (n_58_52), .C1 (n_57_51), .C2 (n_51_54) );
AOI211_X1 g_67_49 (.ZN (n_67_49), .A (n_66_48), .B (n_60_51), .C1 (n_56_53), .C2 (n_53_53) );
AOI211_X1 g_66_51 (.ZN (n_66_51), .A (n_65_50), .B (n_62_50), .C1 (n_58_52), .C2 (n_55_52) );
AOI211_X1 g_65_49 (.ZN (n_65_49), .A (n_67_49), .B (n_64_49), .C1 (n_60_51), .C2 (n_57_51) );
AOI211_X1 g_67_48 (.ZN (n_67_48), .A (n_66_51), .B (n_66_48), .C1 (n_62_50), .C2 (n_56_53) );
AOI211_X1 g_69_47 (.ZN (n_69_47), .A (n_65_49), .B (n_65_50), .C1 (n_64_49), .C2 (n_58_52) );
AOI211_X1 g_71_46 (.ZN (n_71_46), .A (n_67_48), .B (n_67_49), .C1 (n_66_48), .C2 (n_60_51) );
AOI211_X1 g_73_45 (.ZN (n_73_45), .A (n_69_47), .B (n_66_51), .C1 (n_65_50), .C2 (n_62_50) );
AOI211_X1 g_75_44 (.ZN (n_75_44), .A (n_71_46), .B (n_65_49), .C1 (n_67_49), .C2 (n_64_49) );
AOI211_X1 g_77_43 (.ZN (n_77_43), .A (n_73_45), .B (n_67_48), .C1 (n_66_51), .C2 (n_66_48) );
AOI211_X1 g_79_42 (.ZN (n_79_42), .A (n_75_44), .B (n_69_47), .C1 (n_65_49), .C2 (n_65_50) );
AOI211_X1 g_81_41 (.ZN (n_81_41), .A (n_77_43), .B (n_71_46), .C1 (n_67_48), .C2 (n_67_49) );
AOI211_X1 g_83_40 (.ZN (n_83_40), .A (n_79_42), .B (n_73_45), .C1 (n_69_47), .C2 (n_66_51) );
AOI211_X1 g_85_39 (.ZN (n_85_39), .A (n_81_41), .B (n_75_44), .C1 (n_71_46), .C2 (n_65_49) );
AOI211_X1 g_87_38 (.ZN (n_87_38), .A (n_83_40), .B (n_77_43), .C1 (n_73_45), .C2 (n_67_48) );
AOI211_X1 g_89_37 (.ZN (n_89_37), .A (n_85_39), .B (n_79_42), .C1 (n_75_44), .C2 (n_69_47) );
AOI211_X1 g_91_36 (.ZN (n_91_36), .A (n_87_38), .B (n_81_41), .C1 (n_77_43), .C2 (n_71_46) );
AOI211_X1 g_93_37 (.ZN (n_93_37), .A (n_89_37), .B (n_83_40), .C1 (n_79_42), .C2 (n_73_45) );
AOI211_X1 g_91_38 (.ZN (n_91_38), .A (n_91_36), .B (n_85_39), .C1 (n_81_41), .C2 (n_75_44) );
AOI211_X1 g_89_39 (.ZN (n_89_39), .A (n_93_37), .B (n_87_38), .C1 (n_83_40), .C2 (n_77_43) );
AOI211_X1 g_87_40 (.ZN (n_87_40), .A (n_91_38), .B (n_89_37), .C1 (n_85_39), .C2 (n_79_42) );
AOI211_X1 g_85_41 (.ZN (n_85_41), .A (n_89_39), .B (n_91_36), .C1 (n_87_38), .C2 (n_81_41) );
AOI211_X1 g_83_42 (.ZN (n_83_42), .A (n_87_40), .B (n_93_37), .C1 (n_89_37), .C2 (n_83_40) );
AOI211_X1 g_81_43 (.ZN (n_81_43), .A (n_85_41), .B (n_91_38), .C1 (n_91_36), .C2 (n_85_39) );
AOI211_X1 g_79_44 (.ZN (n_79_44), .A (n_83_42), .B (n_89_39), .C1 (n_93_37), .C2 (n_87_38) );
AOI211_X1 g_77_45 (.ZN (n_77_45), .A (n_81_43), .B (n_87_40), .C1 (n_91_38), .C2 (n_89_37) );
AOI211_X1 g_75_46 (.ZN (n_75_46), .A (n_79_44), .B (n_85_41), .C1 (n_89_39), .C2 (n_91_36) );
AOI211_X1 g_73_47 (.ZN (n_73_47), .A (n_77_45), .B (n_83_42), .C1 (n_87_40), .C2 (n_93_37) );
AOI211_X1 g_71_48 (.ZN (n_71_48), .A (n_75_46), .B (n_81_43), .C1 (n_85_41), .C2 (n_91_38) );
AOI211_X1 g_69_49 (.ZN (n_69_49), .A (n_73_47), .B (n_79_44), .C1 (n_83_42), .C2 (n_89_39) );
AOI211_X1 g_67_50 (.ZN (n_67_50), .A (n_71_48), .B (n_77_45), .C1 (n_81_43), .C2 (n_87_40) );
AOI211_X1 g_65_51 (.ZN (n_65_51), .A (n_69_49), .B (n_75_46), .C1 (n_79_44), .C2 (n_85_41) );
AOI211_X1 g_63_50 (.ZN (n_63_50), .A (n_67_50), .B (n_73_47), .C1 (n_77_45), .C2 (n_83_42) );
AOI211_X1 g_61_51 (.ZN (n_61_51), .A (n_65_51), .B (n_71_48), .C1 (n_75_46), .C2 (n_81_43) );
AOI211_X1 g_62_49 (.ZN (n_62_49), .A (n_63_50), .B (n_69_49), .C1 (n_73_47), .C2 (n_79_44) );
AOI211_X1 g_60_50 (.ZN (n_60_50), .A (n_61_51), .B (n_67_50), .C1 (n_71_48), .C2 (n_77_45) );
AOI211_X1 g_58_51 (.ZN (n_58_51), .A (n_62_49), .B (n_65_51), .C1 (n_69_49), .C2 (n_75_46) );
AOI211_X1 g_56_52 (.ZN (n_56_52), .A (n_60_50), .B (n_63_50), .C1 (n_67_50), .C2 (n_73_47) );
AOI211_X1 g_54_53 (.ZN (n_54_53), .A (n_58_51), .B (n_61_51), .C1 (n_65_51), .C2 (n_71_48) );
AOI211_X1 g_52_54 (.ZN (n_52_54), .A (n_56_52), .B (n_62_49), .C1 (n_63_50), .C2 (n_69_49) );
AOI211_X1 g_50_55 (.ZN (n_50_55), .A (n_54_53), .B (n_60_50), .C1 (n_61_51), .C2 (n_67_50) );
AOI211_X1 g_48_56 (.ZN (n_48_56), .A (n_52_54), .B (n_58_51), .C1 (n_62_49), .C2 (n_65_51) );
AOI211_X1 g_46_57 (.ZN (n_46_57), .A (n_50_55), .B (n_56_52), .C1 (n_60_50), .C2 (n_63_50) );
AOI211_X1 g_44_58 (.ZN (n_44_58), .A (n_48_56), .B (n_54_53), .C1 (n_58_51), .C2 (n_61_51) );
AOI211_X1 g_42_59 (.ZN (n_42_59), .A (n_46_57), .B (n_52_54), .C1 (n_56_52), .C2 (n_62_49) );
AOI211_X1 g_40_60 (.ZN (n_40_60), .A (n_44_58), .B (n_50_55), .C1 (n_54_53), .C2 (n_60_50) );
AOI211_X1 g_38_61 (.ZN (n_38_61), .A (n_42_59), .B (n_48_56), .C1 (n_52_54), .C2 (n_58_51) );
AOI211_X1 g_36_62 (.ZN (n_36_62), .A (n_40_60), .B (n_46_57), .C1 (n_50_55), .C2 (n_56_52) );
AOI211_X1 g_34_63 (.ZN (n_34_63), .A (n_38_61), .B (n_44_58), .C1 (n_48_56), .C2 (n_54_53) );
AOI211_X1 g_32_64 (.ZN (n_32_64), .A (n_36_62), .B (n_42_59), .C1 (n_46_57), .C2 (n_52_54) );
AOI211_X1 g_30_65 (.ZN (n_30_65), .A (n_34_63), .B (n_40_60), .C1 (n_44_58), .C2 (n_50_55) );
AOI211_X1 g_28_66 (.ZN (n_28_66), .A (n_32_64), .B (n_38_61), .C1 (n_42_59), .C2 (n_48_56) );
AOI211_X1 g_26_67 (.ZN (n_26_67), .A (n_30_65), .B (n_36_62), .C1 (n_40_60), .C2 (n_46_57) );
AOI211_X1 g_24_68 (.ZN (n_24_68), .A (n_28_66), .B (n_34_63), .C1 (n_38_61), .C2 (n_44_58) );
AOI211_X1 g_22_69 (.ZN (n_22_69), .A (n_26_67), .B (n_32_64), .C1 (n_36_62), .C2 (n_42_59) );
AOI211_X1 g_20_70 (.ZN (n_20_70), .A (n_24_68), .B (n_30_65), .C1 (n_34_63), .C2 (n_40_60) );
AOI211_X1 g_18_71 (.ZN (n_18_71), .A (n_22_69), .B (n_28_66), .C1 (n_32_64), .C2 (n_38_61) );
AOI211_X1 g_16_72 (.ZN (n_16_72), .A (n_20_70), .B (n_26_67), .C1 (n_30_65), .C2 (n_36_62) );
AOI211_X1 g_14_73 (.ZN (n_14_73), .A (n_18_71), .B (n_24_68), .C1 (n_28_66), .C2 (n_34_63) );
AOI211_X1 g_12_74 (.ZN (n_12_74), .A (n_16_72), .B (n_22_69), .C1 (n_26_67), .C2 (n_32_64) );
AOI211_X1 g_11_72 (.ZN (n_11_72), .A (n_14_73), .B (n_20_70), .C1 (n_24_68), .C2 (n_30_65) );
AOI211_X1 g_9_73 (.ZN (n_9_73), .A (n_12_74), .B (n_18_71), .C1 (n_22_69), .C2 (n_28_66) );
AOI211_X1 g_7_74 (.ZN (n_7_74), .A (n_11_72), .B (n_16_72), .C1 (n_20_70), .C2 (n_26_67) );
AOI211_X1 g_6_76 (.ZN (n_6_76), .A (n_9_73), .B (n_14_73), .C1 (n_18_71), .C2 (n_24_68) );
AOI211_X1 g_5_78 (.ZN (n_5_78), .A (n_7_74), .B (n_12_74), .C1 (n_16_72), .C2 (n_22_69) );
AOI211_X1 g_6_80 (.ZN (n_6_80), .A (n_6_76), .B (n_11_72), .C1 (n_14_73), .C2 (n_20_70) );
AOI211_X1 g_7_78 (.ZN (n_7_78), .A (n_5_78), .B (n_9_73), .C1 (n_12_74), .C2 (n_18_71) );
AOI211_X1 g_8_76 (.ZN (n_8_76), .A (n_6_80), .B (n_7_74), .C1 (n_11_72), .C2 (n_16_72) );
AOI211_X1 g_10_75 (.ZN (n_10_75), .A (n_7_78), .B (n_6_76), .C1 (n_9_73), .C2 (n_14_73) );
AOI211_X1 g_9_77 (.ZN (n_9_77), .A (n_8_76), .B (n_5_78), .C1 (n_7_74), .C2 (n_12_74) );
AOI211_X1 g_8_75 (.ZN (n_8_75), .A (n_10_75), .B (n_6_80), .C1 (n_6_76), .C2 (n_11_72) );
AOI211_X1 g_10_74 (.ZN (n_10_74), .A (n_9_77), .B (n_7_78), .C1 (n_5_78), .C2 (n_9_73) );
AOI211_X1 g_12_73 (.ZN (n_12_73), .A (n_8_75), .B (n_8_76), .C1 (n_6_80), .C2 (n_7_74) );
AOI211_X1 g_11_75 (.ZN (n_11_75), .A (n_10_74), .B (n_10_75), .C1 (n_7_78), .C2 (n_6_76) );
AOI211_X1 g_13_74 (.ZN (n_13_74), .A (n_12_73), .B (n_9_77), .C1 (n_8_76), .C2 (n_5_78) );
AOI211_X1 g_15_73 (.ZN (n_15_73), .A (n_11_75), .B (n_8_75), .C1 (n_10_75), .C2 (n_6_80) );
AOI211_X1 g_17_72 (.ZN (n_17_72), .A (n_13_74), .B (n_10_74), .C1 (n_9_77), .C2 (n_7_78) );
AOI211_X1 g_19_71 (.ZN (n_19_71), .A (n_15_73), .B (n_12_73), .C1 (n_8_75), .C2 (n_8_76) );
AOI211_X1 g_21_70 (.ZN (n_21_70), .A (n_17_72), .B (n_11_75), .C1 (n_10_74), .C2 (n_10_75) );
AOI211_X1 g_23_69 (.ZN (n_23_69), .A (n_19_71), .B (n_13_74), .C1 (n_12_73), .C2 (n_9_77) );
AOI211_X1 g_24_67 (.ZN (n_24_67), .A (n_21_70), .B (n_15_73), .C1 (n_11_75), .C2 (n_8_75) );
AOI211_X1 g_26_66 (.ZN (n_26_66), .A (n_23_69), .B (n_17_72), .C1 (n_13_74), .C2 (n_10_74) );
AOI211_X1 g_28_65 (.ZN (n_28_65), .A (n_24_67), .B (n_19_71), .C1 (n_15_73), .C2 (n_12_73) );
AOI211_X1 g_30_64 (.ZN (n_30_64), .A (n_26_66), .B (n_21_70), .C1 (n_17_72), .C2 (n_11_75) );
AOI211_X1 g_32_63 (.ZN (n_32_63), .A (n_28_65), .B (n_23_69), .C1 (n_19_71), .C2 (n_13_74) );
AOI211_X1 g_34_62 (.ZN (n_34_62), .A (n_30_64), .B (n_24_67), .C1 (n_21_70), .C2 (n_15_73) );
AOI211_X1 g_36_61 (.ZN (n_36_61), .A (n_32_63), .B (n_26_66), .C1 (n_23_69), .C2 (n_17_72) );
AOI211_X1 g_35_63 (.ZN (n_35_63), .A (n_34_62), .B (n_28_65), .C1 (n_24_67), .C2 (n_19_71) );
AOI211_X1 g_37_62 (.ZN (n_37_62), .A (n_36_61), .B (n_30_64), .C1 (n_26_66), .C2 (n_21_70) );
AOI211_X1 g_39_61 (.ZN (n_39_61), .A (n_35_63), .B (n_32_63), .C1 (n_28_65), .C2 (n_23_69) );
AOI211_X1 g_41_60 (.ZN (n_41_60), .A (n_37_62), .B (n_34_62), .C1 (n_30_64), .C2 (n_24_67) );
AOI211_X1 g_43_59 (.ZN (n_43_59), .A (n_39_61), .B (n_36_61), .C1 (n_32_63), .C2 (n_26_66) );
AOI211_X1 g_45_58 (.ZN (n_45_58), .A (n_41_60), .B (n_35_63), .C1 (n_34_62), .C2 (n_28_65) );
AOI211_X1 g_47_57 (.ZN (n_47_57), .A (n_43_59), .B (n_37_62), .C1 (n_36_61), .C2 (n_30_64) );
AOI211_X1 g_49_56 (.ZN (n_49_56), .A (n_45_58), .B (n_39_61), .C1 (n_35_63), .C2 (n_32_63) );
AOI211_X1 g_51_55 (.ZN (n_51_55), .A (n_47_57), .B (n_41_60), .C1 (n_37_62), .C2 (n_34_62) );
AOI211_X1 g_53_54 (.ZN (n_53_54), .A (n_49_56), .B (n_43_59), .C1 (n_39_61), .C2 (n_36_61) );
AOI211_X1 g_52_56 (.ZN (n_52_56), .A (n_51_55), .B (n_45_58), .C1 (n_41_60), .C2 (n_35_63) );
AOI211_X1 g_54_55 (.ZN (n_54_55), .A (n_53_54), .B (n_47_57), .C1 (n_43_59), .C2 (n_37_62) );
AOI211_X1 g_56_54 (.ZN (n_56_54), .A (n_52_56), .B (n_49_56), .C1 (n_45_58), .C2 (n_39_61) );
AOI211_X1 g_58_53 (.ZN (n_58_53), .A (n_54_55), .B (n_51_55), .C1 (n_47_57), .C2 (n_41_60) );
AOI211_X1 g_60_52 (.ZN (n_60_52), .A (n_56_54), .B (n_53_54), .C1 (n_49_56), .C2 (n_43_59) );
AOI211_X1 g_62_51 (.ZN (n_62_51), .A (n_58_53), .B (n_52_56), .C1 (n_51_55), .C2 (n_45_58) );
AOI211_X1 g_64_52 (.ZN (n_64_52), .A (n_60_52), .B (n_54_55), .C1 (n_53_54), .C2 (n_47_57) );
AOI211_X1 g_62_53 (.ZN (n_62_53), .A (n_62_51), .B (n_56_54), .C1 (n_52_56), .C2 (n_49_56) );
AOI211_X1 g_63_51 (.ZN (n_63_51), .A (n_64_52), .B (n_58_53), .C1 (n_54_55), .C2 (n_51_55) );
AOI211_X1 g_61_52 (.ZN (n_61_52), .A (n_62_53), .B (n_60_52), .C1 (n_56_54), .C2 (n_53_54) );
AOI211_X1 g_59_53 (.ZN (n_59_53), .A (n_63_51), .B (n_62_51), .C1 (n_58_53), .C2 (n_52_56) );
AOI211_X1 g_57_54 (.ZN (n_57_54), .A (n_61_52), .B (n_64_52), .C1 (n_60_52), .C2 (n_54_55) );
AOI211_X1 g_55_55 (.ZN (n_55_55), .A (n_59_53), .B (n_62_53), .C1 (n_62_51), .C2 (n_56_54) );
AOI211_X1 g_53_56 (.ZN (n_53_56), .A (n_57_54), .B (n_63_51), .C1 (n_64_52), .C2 (n_58_53) );
AOI211_X1 g_54_54 (.ZN (n_54_54), .A (n_55_55), .B (n_61_52), .C1 (n_62_53), .C2 (n_60_52) );
AOI211_X1 g_52_55 (.ZN (n_52_55), .A (n_53_56), .B (n_59_53), .C1 (n_63_51), .C2 (n_62_51) );
AOI211_X1 g_50_56 (.ZN (n_50_56), .A (n_54_54), .B (n_57_54), .C1 (n_61_52), .C2 (n_64_52) );
AOI211_X1 g_48_57 (.ZN (n_48_57), .A (n_52_55), .B (n_55_55), .C1 (n_59_53), .C2 (n_62_53) );
AOI211_X1 g_46_58 (.ZN (n_46_58), .A (n_50_56), .B (n_53_56), .C1 (n_57_54), .C2 (n_63_51) );
AOI211_X1 g_44_59 (.ZN (n_44_59), .A (n_48_57), .B (n_54_54), .C1 (n_55_55), .C2 (n_61_52) );
AOI211_X1 g_42_60 (.ZN (n_42_60), .A (n_46_58), .B (n_52_55), .C1 (n_53_56), .C2 (n_59_53) );
AOI211_X1 g_40_61 (.ZN (n_40_61), .A (n_44_59), .B (n_50_56), .C1 (n_54_54), .C2 (n_57_54) );
AOI211_X1 g_38_62 (.ZN (n_38_62), .A (n_42_60), .B (n_48_57), .C1 (n_52_55), .C2 (n_55_55) );
AOI211_X1 g_36_63 (.ZN (n_36_63), .A (n_40_61), .B (n_46_58), .C1 (n_50_56), .C2 (n_53_56) );
AOI211_X1 g_34_64 (.ZN (n_34_64), .A (n_38_62), .B (n_44_59), .C1 (n_48_57), .C2 (n_54_54) );
AOI211_X1 g_32_65 (.ZN (n_32_65), .A (n_36_63), .B (n_42_60), .C1 (n_46_58), .C2 (n_52_55) );
AOI211_X1 g_30_66 (.ZN (n_30_66), .A (n_34_64), .B (n_40_61), .C1 (n_44_59), .C2 (n_50_56) );
AOI211_X1 g_28_67 (.ZN (n_28_67), .A (n_32_65), .B (n_38_62), .C1 (n_42_60), .C2 (n_48_57) );
AOI211_X1 g_26_68 (.ZN (n_26_68), .A (n_30_66), .B (n_36_63), .C1 (n_40_61), .C2 (n_46_58) );
AOI211_X1 g_24_69 (.ZN (n_24_69), .A (n_28_67), .B (n_34_64), .C1 (n_38_62), .C2 (n_44_59) );
AOI211_X1 g_22_70 (.ZN (n_22_70), .A (n_26_68), .B (n_32_65), .C1 (n_36_63), .C2 (n_42_60) );
AOI211_X1 g_20_71 (.ZN (n_20_71), .A (n_24_69), .B (n_30_66), .C1 (n_34_64), .C2 (n_40_61) );
AOI211_X1 g_18_72 (.ZN (n_18_72), .A (n_22_70), .B (n_28_67), .C1 (n_32_65), .C2 (n_38_62) );
AOI211_X1 g_16_73 (.ZN (n_16_73), .A (n_20_71), .B (n_26_68), .C1 (n_30_66), .C2 (n_36_63) );
AOI211_X1 g_17_71 (.ZN (n_17_71), .A (n_18_72), .B (n_24_69), .C1 (n_28_67), .C2 (n_34_64) );
AOI211_X1 g_15_72 (.ZN (n_15_72), .A (n_16_73), .B (n_22_70), .C1 (n_26_68), .C2 (n_32_65) );
AOI211_X1 g_13_73 (.ZN (n_13_73), .A (n_17_71), .B (n_20_71), .C1 (n_24_69), .C2 (n_30_66) );
AOI211_X1 g_11_74 (.ZN (n_11_74), .A (n_15_72), .B (n_18_72), .C1 (n_22_70), .C2 (n_28_67) );
AOI211_X1 g_9_75 (.ZN (n_9_75), .A (n_13_73), .B (n_16_73), .C1 (n_20_71), .C2 (n_26_68) );
AOI211_X1 g_7_76 (.ZN (n_7_76), .A (n_11_74), .B (n_17_71), .C1 (n_18_72), .C2 (n_24_69) );
AOI211_X1 g_6_78 (.ZN (n_6_78), .A (n_9_75), .B (n_15_72), .C1 (n_16_73), .C2 (n_22_70) );
AOI211_X1 g_8_77 (.ZN (n_8_77), .A (n_7_76), .B (n_13_73), .C1 (n_17_71), .C2 (n_20_71) );
AOI211_X1 g_10_76 (.ZN (n_10_76), .A (n_6_78), .B (n_11_74), .C1 (n_15_72), .C2 (n_18_72) );
AOI211_X1 g_12_75 (.ZN (n_12_75), .A (n_8_77), .B (n_9_75), .C1 (n_13_73), .C2 (n_16_73) );
AOI211_X1 g_14_74 (.ZN (n_14_74), .A (n_10_76), .B (n_7_76), .C1 (n_11_74), .C2 (n_17_71) );
AOI211_X1 g_13_76 (.ZN (n_13_76), .A (n_12_75), .B (n_6_78), .C1 (n_9_75), .C2 (n_15_72) );
AOI211_X1 g_15_75 (.ZN (n_15_75), .A (n_14_74), .B (n_8_77), .C1 (n_7_76), .C2 (n_13_73) );
AOI211_X1 g_17_74 (.ZN (n_17_74), .A (n_13_76), .B (n_10_76), .C1 (n_6_78), .C2 (n_11_74) );
AOI211_X1 g_19_73 (.ZN (n_19_73), .A (n_15_75), .B (n_12_75), .C1 (n_8_77), .C2 (n_9_75) );
AOI211_X1 g_21_72 (.ZN (n_21_72), .A (n_17_74), .B (n_14_74), .C1 (n_10_76), .C2 (n_7_76) );
AOI211_X1 g_23_71 (.ZN (n_23_71), .A (n_19_73), .B (n_13_76), .C1 (n_12_75), .C2 (n_6_78) );
AOI211_X1 g_25_70 (.ZN (n_25_70), .A (n_21_72), .B (n_15_75), .C1 (n_14_74), .C2 (n_8_77) );
AOI211_X1 g_27_69 (.ZN (n_27_69), .A (n_23_71), .B (n_17_74), .C1 (n_13_76), .C2 (n_10_76) );
AOI211_X1 g_25_68 (.ZN (n_25_68), .A (n_25_70), .B (n_19_73), .C1 (n_15_75), .C2 (n_12_75) );
AOI211_X1 g_27_67 (.ZN (n_27_67), .A (n_27_69), .B (n_21_72), .C1 (n_17_74), .C2 (n_14_74) );
AOI211_X1 g_29_66 (.ZN (n_29_66), .A (n_25_68), .B (n_23_71), .C1 (n_19_73), .C2 (n_13_76) );
AOI211_X1 g_31_65 (.ZN (n_31_65), .A (n_27_67), .B (n_25_70), .C1 (n_21_72), .C2 (n_15_75) );
AOI211_X1 g_33_64 (.ZN (n_33_64), .A (n_29_66), .B (n_27_69), .C1 (n_23_71), .C2 (n_17_74) );
AOI211_X1 g_32_66 (.ZN (n_32_66), .A (n_31_65), .B (n_25_68), .C1 (n_25_70), .C2 (n_19_73) );
AOI211_X1 g_34_65 (.ZN (n_34_65), .A (n_33_64), .B (n_27_67), .C1 (n_27_69), .C2 (n_21_72) );
AOI211_X1 g_36_64 (.ZN (n_36_64), .A (n_32_66), .B (n_29_66), .C1 (n_25_68), .C2 (n_23_71) );
AOI211_X1 g_38_63 (.ZN (n_38_63), .A (n_34_65), .B (n_31_65), .C1 (n_27_67), .C2 (n_25_70) );
AOI211_X1 g_40_62 (.ZN (n_40_62), .A (n_36_64), .B (n_33_64), .C1 (n_29_66), .C2 (n_27_69) );
AOI211_X1 g_42_61 (.ZN (n_42_61), .A (n_38_63), .B (n_32_66), .C1 (n_31_65), .C2 (n_25_68) );
AOI211_X1 g_44_60 (.ZN (n_44_60), .A (n_40_62), .B (n_34_65), .C1 (n_33_64), .C2 (n_27_67) );
AOI211_X1 g_46_59 (.ZN (n_46_59), .A (n_42_61), .B (n_36_64), .C1 (n_32_66), .C2 (n_29_66) );
AOI211_X1 g_48_58 (.ZN (n_48_58), .A (n_44_60), .B (n_38_63), .C1 (n_34_65), .C2 (n_31_65) );
AOI211_X1 g_50_57 (.ZN (n_50_57), .A (n_46_59), .B (n_40_62), .C1 (n_36_64), .C2 (n_33_64) );
AOI211_X1 g_49_59 (.ZN (n_49_59), .A (n_48_58), .B (n_42_61), .C1 (n_38_63), .C2 (n_32_66) );
AOI211_X1 g_47_58 (.ZN (n_47_58), .A (n_50_57), .B (n_44_60), .C1 (n_40_62), .C2 (n_34_65) );
AOI211_X1 g_49_57 (.ZN (n_49_57), .A (n_49_59), .B (n_46_59), .C1 (n_42_61), .C2 (n_36_64) );
AOI211_X1 g_51_56 (.ZN (n_51_56), .A (n_47_58), .B (n_48_58), .C1 (n_44_60), .C2 (n_38_63) );
AOI211_X1 g_53_55 (.ZN (n_53_55), .A (n_49_57), .B (n_50_57), .C1 (n_46_59), .C2 (n_40_62) );
AOI211_X1 g_55_54 (.ZN (n_55_54), .A (n_51_56), .B (n_49_59), .C1 (n_48_58), .C2 (n_42_61) );
AOI211_X1 g_57_53 (.ZN (n_57_53), .A (n_53_55), .B (n_47_58), .C1 (n_50_57), .C2 (n_44_60) );
AOI211_X1 g_59_52 (.ZN (n_59_52), .A (n_55_54), .B (n_49_57), .C1 (n_49_59), .C2 (n_46_59) );
AOI211_X1 g_60_54 (.ZN (n_60_54), .A (n_57_53), .B (n_51_56), .C1 (n_47_58), .C2 (n_48_58) );
AOI211_X1 g_58_55 (.ZN (n_58_55), .A (n_59_52), .B (n_53_55), .C1 (n_49_57), .C2 (n_50_57) );
AOI211_X1 g_56_56 (.ZN (n_56_56), .A (n_60_54), .B (n_55_54), .C1 (n_51_56), .C2 (n_49_59) );
AOI211_X1 g_54_57 (.ZN (n_54_57), .A (n_58_55), .B (n_57_53), .C1 (n_53_55), .C2 (n_47_58) );
AOI211_X1 g_52_58 (.ZN (n_52_58), .A (n_56_56), .B (n_59_52), .C1 (n_55_54), .C2 (n_49_57) );
AOI211_X1 g_50_59 (.ZN (n_50_59), .A (n_54_57), .B (n_60_54), .C1 (n_57_53), .C2 (n_51_56) );
AOI211_X1 g_51_57 (.ZN (n_51_57), .A (n_52_58), .B (n_58_55), .C1 (n_59_52), .C2 (n_53_55) );
AOI211_X1 g_49_58 (.ZN (n_49_58), .A (n_50_59), .B (n_56_56), .C1 (n_60_54), .C2 (n_55_54) );
AOI211_X1 g_47_59 (.ZN (n_47_59), .A (n_51_57), .B (n_54_57), .C1 (n_58_55), .C2 (n_57_53) );
AOI211_X1 g_45_60 (.ZN (n_45_60), .A (n_49_58), .B (n_52_58), .C1 (n_56_56), .C2 (n_59_52) );
AOI211_X1 g_43_61 (.ZN (n_43_61), .A (n_47_59), .B (n_50_59), .C1 (n_54_57), .C2 (n_60_54) );
AOI211_X1 g_41_62 (.ZN (n_41_62), .A (n_45_60), .B (n_51_57), .C1 (n_52_58), .C2 (n_58_55) );
AOI211_X1 g_39_63 (.ZN (n_39_63), .A (n_43_61), .B (n_49_58), .C1 (n_50_59), .C2 (n_56_56) );
AOI211_X1 g_37_64 (.ZN (n_37_64), .A (n_41_62), .B (n_47_59), .C1 (n_51_57), .C2 (n_54_57) );
AOI211_X1 g_35_65 (.ZN (n_35_65), .A (n_39_63), .B (n_45_60), .C1 (n_49_58), .C2 (n_52_58) );
AOI211_X1 g_33_66 (.ZN (n_33_66), .A (n_37_64), .B (n_43_61), .C1 (n_47_59), .C2 (n_50_59) );
AOI211_X1 g_31_67 (.ZN (n_31_67), .A (n_35_65), .B (n_41_62), .C1 (n_45_60), .C2 (n_51_57) );
AOI211_X1 g_29_68 (.ZN (n_29_68), .A (n_33_66), .B (n_39_63), .C1 (n_43_61), .C2 (n_49_58) );
AOI211_X1 g_28_70 (.ZN (n_28_70), .A (n_31_67), .B (n_37_64), .C1 (n_41_62), .C2 (n_47_59) );
AOI211_X1 g_27_68 (.ZN (n_27_68), .A (n_29_68), .B (n_35_65), .C1 (n_39_63), .C2 (n_45_60) );
AOI211_X1 g_29_67 (.ZN (n_29_67), .A (n_28_70), .B (n_33_66), .C1 (n_37_64), .C2 (n_43_61) );
AOI211_X1 g_31_66 (.ZN (n_31_66), .A (n_27_68), .B (n_31_67), .C1 (n_35_65), .C2 (n_41_62) );
AOI211_X1 g_33_65 (.ZN (n_33_65), .A (n_29_67), .B (n_29_68), .C1 (n_33_66), .C2 (n_39_63) );
AOI211_X1 g_35_64 (.ZN (n_35_64), .A (n_31_66), .B (n_28_70), .C1 (n_31_67), .C2 (n_37_64) );
AOI211_X1 g_37_63 (.ZN (n_37_63), .A (n_33_65), .B (n_27_68), .C1 (n_29_68), .C2 (n_35_65) );
AOI211_X1 g_39_62 (.ZN (n_39_62), .A (n_35_64), .B (n_29_67), .C1 (n_28_70), .C2 (n_33_66) );
AOI211_X1 g_41_61 (.ZN (n_41_61), .A (n_37_63), .B (n_31_66), .C1 (n_27_68), .C2 (n_31_67) );
AOI211_X1 g_43_60 (.ZN (n_43_60), .A (n_39_62), .B (n_33_65), .C1 (n_29_67), .C2 (n_29_68) );
AOI211_X1 g_45_59 (.ZN (n_45_59), .A (n_41_61), .B (n_35_64), .C1 (n_31_66), .C2 (n_28_70) );
AOI211_X1 g_47_60 (.ZN (n_47_60), .A (n_43_60), .B (n_37_63), .C1 (n_33_65), .C2 (n_27_68) );
AOI211_X1 g_45_61 (.ZN (n_45_61), .A (n_45_59), .B (n_39_62), .C1 (n_35_64), .C2 (n_29_67) );
AOI211_X1 g_43_62 (.ZN (n_43_62), .A (n_47_60), .B (n_41_61), .C1 (n_37_63), .C2 (n_31_66) );
AOI211_X1 g_41_63 (.ZN (n_41_63), .A (n_45_61), .B (n_43_60), .C1 (n_39_62), .C2 (n_33_65) );
AOI211_X1 g_39_64 (.ZN (n_39_64), .A (n_43_62), .B (n_45_59), .C1 (n_41_61), .C2 (n_35_64) );
AOI211_X1 g_37_65 (.ZN (n_37_65), .A (n_41_63), .B (n_47_60), .C1 (n_43_60), .C2 (n_37_63) );
AOI211_X1 g_35_66 (.ZN (n_35_66), .A (n_39_64), .B (n_45_61), .C1 (n_45_59), .C2 (n_39_62) );
AOI211_X1 g_33_67 (.ZN (n_33_67), .A (n_37_65), .B (n_43_62), .C1 (n_47_60), .C2 (n_41_61) );
AOI211_X1 g_31_68 (.ZN (n_31_68), .A (n_35_66), .B (n_41_63), .C1 (n_45_61), .C2 (n_43_60) );
AOI211_X1 g_29_69 (.ZN (n_29_69), .A (n_33_67), .B (n_39_64), .C1 (n_43_62), .C2 (n_45_59) );
AOI211_X1 g_30_67 (.ZN (n_30_67), .A (n_31_68), .B (n_37_65), .C1 (n_41_63), .C2 (n_47_60) );
AOI211_X1 g_28_68 (.ZN (n_28_68), .A (n_29_69), .B (n_35_66), .C1 (n_39_64), .C2 (n_45_61) );
AOI211_X1 g_26_69 (.ZN (n_26_69), .A (n_30_67), .B (n_33_67), .C1 (n_37_65), .C2 (n_43_62) );
AOI211_X1 g_24_70 (.ZN (n_24_70), .A (n_28_68), .B (n_31_68), .C1 (n_35_66), .C2 (n_41_63) );
AOI211_X1 g_22_71 (.ZN (n_22_71), .A (n_26_69), .B (n_29_69), .C1 (n_33_67), .C2 (n_39_64) );
AOI211_X1 g_20_72 (.ZN (n_20_72), .A (n_24_70), .B (n_30_67), .C1 (n_31_68), .C2 (n_37_65) );
AOI211_X1 g_18_73 (.ZN (n_18_73), .A (n_22_71), .B (n_28_68), .C1 (n_29_69), .C2 (n_35_66) );
AOI211_X1 g_16_74 (.ZN (n_16_74), .A (n_20_72), .B (n_26_69), .C1 (n_30_67), .C2 (n_33_67) );
AOI211_X1 g_14_75 (.ZN (n_14_75), .A (n_18_73), .B (n_24_70), .C1 (n_28_68), .C2 (n_31_68) );
AOI211_X1 g_12_76 (.ZN (n_12_76), .A (n_16_74), .B (n_22_71), .C1 (n_26_69), .C2 (n_29_69) );
AOI211_X1 g_10_77 (.ZN (n_10_77), .A (n_14_75), .B (n_20_72), .C1 (n_24_70), .C2 (n_30_67) );
AOI211_X1 g_8_78 (.ZN (n_8_78), .A (n_12_76), .B (n_18_73), .C1 (n_22_71), .C2 (n_28_68) );
AOI211_X1 g_9_76 (.ZN (n_9_76), .A (n_10_77), .B (n_16_74), .C1 (n_20_72), .C2 (n_26_69) );
AOI211_X1 g_7_77 (.ZN (n_7_77), .A (n_8_78), .B (n_14_75), .C1 (n_18_73), .C2 (n_24_70) );
AOI211_X1 g_6_79 (.ZN (n_6_79), .A (n_9_76), .B (n_12_76), .C1 (n_16_74), .C2 (n_22_71) );
AOI211_X1 g_5_81 (.ZN (n_5_81), .A (n_7_77), .B (n_10_77), .C1 (n_14_75), .C2 (n_20_72) );
AOI211_X1 g_7_80 (.ZN (n_7_80), .A (n_6_79), .B (n_8_78), .C1 (n_12_76), .C2 (n_18_73) );
AOI211_X1 g_9_79 (.ZN (n_9_79), .A (n_5_81), .B (n_9_76), .C1 (n_10_77), .C2 (n_16_74) );
AOI211_X1 g_11_78 (.ZN (n_11_78), .A (n_7_80), .B (n_7_77), .C1 (n_8_78), .C2 (n_14_75) );
AOI211_X1 g_13_77 (.ZN (n_13_77), .A (n_9_79), .B (n_6_79), .C1 (n_9_76), .C2 (n_12_76) );
AOI211_X1 g_11_76 (.ZN (n_11_76), .A (n_11_78), .B (n_5_81), .C1 (n_7_77), .C2 (n_10_77) );
AOI211_X1 g_13_75 (.ZN (n_13_75), .A (n_13_77), .B (n_7_80), .C1 (n_6_79), .C2 (n_8_78) );
AOI211_X1 g_15_74 (.ZN (n_15_74), .A (n_11_76), .B (n_9_79), .C1 (n_5_81), .C2 (n_9_76) );
AOI211_X1 g_17_73 (.ZN (n_17_73), .A (n_13_75), .B (n_11_78), .C1 (n_7_80), .C2 (n_7_77) );
AOI211_X1 g_19_72 (.ZN (n_19_72), .A (n_15_74), .B (n_13_77), .C1 (n_9_79), .C2 (n_6_79) );
AOI211_X1 g_21_71 (.ZN (n_21_71), .A (n_17_73), .B (n_11_76), .C1 (n_11_78), .C2 (n_5_81) );
AOI211_X1 g_23_70 (.ZN (n_23_70), .A (n_19_72), .B (n_13_75), .C1 (n_13_77), .C2 (n_7_80) );
AOI211_X1 g_25_69 (.ZN (n_25_69), .A (n_21_71), .B (n_15_74), .C1 (n_11_76), .C2 (n_9_79) );
AOI211_X1 g_26_71 (.ZN (n_26_71), .A (n_23_70), .B (n_17_73), .C1 (n_13_75), .C2 (n_11_78) );
AOI211_X1 g_24_72 (.ZN (n_24_72), .A (n_25_69), .B (n_19_72), .C1 (n_15_74), .C2 (n_13_77) );
AOI211_X1 g_22_73 (.ZN (n_22_73), .A (n_26_71), .B (n_21_71), .C1 (n_17_73), .C2 (n_11_76) );
AOI211_X1 g_20_74 (.ZN (n_20_74), .A (n_24_72), .B (n_23_70), .C1 (n_19_72), .C2 (n_13_75) );
AOI211_X1 g_18_75 (.ZN (n_18_75), .A (n_22_73), .B (n_25_69), .C1 (n_21_71), .C2 (n_15_74) );
AOI211_X1 g_16_76 (.ZN (n_16_76), .A (n_20_74), .B (n_26_71), .C1 (n_23_70), .C2 (n_17_73) );
AOI211_X1 g_14_77 (.ZN (n_14_77), .A (n_18_75), .B (n_24_72), .C1 (n_25_69), .C2 (n_19_72) );
AOI211_X1 g_12_78 (.ZN (n_12_78), .A (n_16_76), .B (n_22_73), .C1 (n_26_71), .C2 (n_21_71) );
AOI211_X1 g_10_79 (.ZN (n_10_79), .A (n_14_77), .B (n_20_74), .C1 (n_24_72), .C2 (n_23_70) );
AOI211_X1 g_11_77 (.ZN (n_11_77), .A (n_12_78), .B (n_18_75), .C1 (n_22_73), .C2 (n_25_69) );
AOI211_X1 g_9_78 (.ZN (n_9_78), .A (n_10_79), .B (n_16_76), .C1 (n_20_74), .C2 (n_26_71) );
AOI211_X1 g_7_79 (.ZN (n_7_79), .A (n_11_77), .B (n_14_77), .C1 (n_18_75), .C2 (n_24_72) );
AOI211_X1 g_5_80 (.ZN (n_5_80), .A (n_9_78), .B (n_12_78), .C1 (n_16_76), .C2 (n_22_73) );
AOI211_X1 g_4_82 (.ZN (n_4_82), .A (n_7_79), .B (n_10_79), .C1 (n_14_77), .C2 (n_20_74) );
AOI211_X1 g_6_81 (.ZN (n_6_81), .A (n_5_80), .B (n_11_77), .C1 (n_12_78), .C2 (n_18_75) );
AOI211_X1 g_8_80 (.ZN (n_8_80), .A (n_4_82), .B (n_9_78), .C1 (n_10_79), .C2 (n_16_76) );
AOI211_X1 g_7_82 (.ZN (n_7_82), .A (n_6_81), .B (n_7_79), .C1 (n_11_77), .C2 (n_14_77) );
AOI211_X1 g_5_83 (.ZN (n_5_83), .A (n_8_80), .B (n_5_80), .C1 (n_9_78), .C2 (n_12_78) );
AOI211_X1 g_3_84 (.ZN (n_3_84), .A (n_7_82), .B (n_4_82), .C1 (n_7_79), .C2 (n_10_79) );
AOI211_X1 g_2_86 (.ZN (n_2_86), .A (n_5_83), .B (n_6_81), .C1 (n_5_80), .C2 (n_11_77) );
AOI211_X1 g_1_88 (.ZN (n_1_88), .A (n_3_84), .B (n_8_80), .C1 (n_4_82), .C2 (n_9_78) );
AOI211_X1 g_3_87 (.ZN (n_3_87), .A (n_2_86), .B (n_7_82), .C1 (n_6_81), .C2 (n_7_79) );
AOI211_X1 g_4_85 (.ZN (n_4_85), .A (n_1_88), .B (n_5_83), .C1 (n_8_80), .C2 (n_5_80) );
AOI211_X1 g_6_84 (.ZN (n_6_84), .A (n_3_87), .B (n_3_84), .C1 (n_7_82), .C2 (n_4_82) );
AOI211_X1 g_4_83 (.ZN (n_4_83), .A (n_4_85), .B (n_2_86), .C1 (n_5_83), .C2 (n_6_81) );
AOI211_X1 g_3_85 (.ZN (n_3_85), .A (n_6_84), .B (n_1_88), .C1 (n_3_84), .C2 (n_8_80) );
AOI211_X1 g_5_86 (.ZN (n_5_86), .A (n_4_83), .B (n_3_87), .C1 (n_2_86), .C2 (n_7_82) );
AOI211_X1 g_7_85 (.ZN (n_7_85), .A (n_3_85), .B (n_4_85), .C1 (n_1_88), .C2 (n_5_83) );
AOI211_X1 g_6_83 (.ZN (n_6_83), .A (n_5_86), .B (n_6_84), .C1 (n_3_87), .C2 (n_3_84) );
AOI211_X1 g_7_81 (.ZN (n_7_81), .A (n_7_85), .B (n_4_83), .C1 (n_4_85), .C2 (n_2_86) );
AOI211_X1 g_8_79 (.ZN (n_8_79), .A (n_6_83), .B (n_3_85), .C1 (n_6_84), .C2 (n_1_88) );
AOI211_X1 g_10_78 (.ZN (n_10_78), .A (n_7_81), .B (n_5_86), .C1 (n_4_83), .C2 (n_3_87) );
AOI211_X1 g_12_77 (.ZN (n_12_77), .A (n_8_79), .B (n_7_85), .C1 (n_3_85), .C2 (n_4_85) );
AOI211_X1 g_14_76 (.ZN (n_14_76), .A (n_10_78), .B (n_6_83), .C1 (n_5_86), .C2 (n_6_84) );
AOI211_X1 g_16_75 (.ZN (n_16_75), .A (n_12_77), .B (n_7_81), .C1 (n_7_85), .C2 (n_4_83) );
AOI211_X1 g_18_74 (.ZN (n_18_74), .A (n_14_76), .B (n_8_79), .C1 (n_6_83), .C2 (n_3_85) );
AOI211_X1 g_20_73 (.ZN (n_20_73), .A (n_16_75), .B (n_10_78), .C1 (n_7_81), .C2 (n_5_86) );
AOI211_X1 g_22_72 (.ZN (n_22_72), .A (n_18_74), .B (n_12_77), .C1 (n_8_79), .C2 (n_7_85) );
AOI211_X1 g_24_71 (.ZN (n_24_71), .A (n_20_73), .B (n_14_76), .C1 (n_10_78), .C2 (n_6_83) );
AOI211_X1 g_26_70 (.ZN (n_26_70), .A (n_22_72), .B (n_16_75), .C1 (n_12_77), .C2 (n_7_81) );
AOI211_X1 g_28_69 (.ZN (n_28_69), .A (n_24_71), .B (n_18_74), .C1 (n_14_76), .C2 (n_8_79) );
AOI211_X1 g_30_68 (.ZN (n_30_68), .A (n_26_70), .B (n_20_73), .C1 (n_16_75), .C2 (n_10_78) );
AOI211_X1 g_32_67 (.ZN (n_32_67), .A (n_28_69), .B (n_22_72), .C1 (n_18_74), .C2 (n_12_77) );
AOI211_X1 g_34_66 (.ZN (n_34_66), .A (n_30_68), .B (n_24_71), .C1 (n_20_73), .C2 (n_14_76) );
AOI211_X1 g_36_65 (.ZN (n_36_65), .A (n_32_67), .B (n_26_70), .C1 (n_22_72), .C2 (n_16_75) );
AOI211_X1 g_38_64 (.ZN (n_38_64), .A (n_34_66), .B (n_28_69), .C1 (n_24_71), .C2 (n_18_74) );
AOI211_X1 g_40_63 (.ZN (n_40_63), .A (n_36_65), .B (n_30_68), .C1 (n_26_70), .C2 (n_20_73) );
AOI211_X1 g_42_62 (.ZN (n_42_62), .A (n_38_64), .B (n_32_67), .C1 (n_28_69), .C2 (n_22_72) );
AOI211_X1 g_44_61 (.ZN (n_44_61), .A (n_40_63), .B (n_34_66), .C1 (n_30_68), .C2 (n_24_71) );
AOI211_X1 g_46_60 (.ZN (n_46_60), .A (n_42_62), .B (n_36_65), .C1 (n_32_67), .C2 (n_26_70) );
AOI211_X1 g_48_59 (.ZN (n_48_59), .A (n_44_61), .B (n_38_64), .C1 (n_34_66), .C2 (n_28_69) );
AOI211_X1 g_50_58 (.ZN (n_50_58), .A (n_46_60), .B (n_40_63), .C1 (n_36_65), .C2 (n_30_68) );
AOI211_X1 g_52_57 (.ZN (n_52_57), .A (n_48_59), .B (n_42_62), .C1 (n_38_64), .C2 (n_32_67) );
AOI211_X1 g_54_56 (.ZN (n_54_56), .A (n_50_58), .B (n_44_61), .C1 (n_40_63), .C2 (n_34_66) );
AOI211_X1 g_56_55 (.ZN (n_56_55), .A (n_52_57), .B (n_46_60), .C1 (n_42_62), .C2 (n_36_65) );
AOI211_X1 g_58_54 (.ZN (n_58_54), .A (n_54_56), .B (n_48_59), .C1 (n_44_61), .C2 (n_38_64) );
AOI211_X1 g_60_53 (.ZN (n_60_53), .A (n_56_55), .B (n_50_58), .C1 (n_46_60), .C2 (n_40_63) );
AOI211_X1 g_62_52 (.ZN (n_62_52), .A (n_58_54), .B (n_52_57), .C1 (n_48_59), .C2 (n_42_62) );
AOI211_X1 g_64_51 (.ZN (n_64_51), .A (n_60_53), .B (n_54_56), .C1 (n_50_58), .C2 (n_44_61) );
AOI211_X1 g_66_50 (.ZN (n_66_50), .A (n_62_52), .B (n_56_55), .C1 (n_52_57), .C2 (n_46_60) );
AOI211_X1 g_68_49 (.ZN (n_68_49), .A (n_64_51), .B (n_58_54), .C1 (n_54_56), .C2 (n_48_59) );
AOI211_X1 g_70_48 (.ZN (n_70_48), .A (n_66_50), .B (n_60_53), .C1 (n_56_55), .C2 (n_50_58) );
AOI211_X1 g_72_47 (.ZN (n_72_47), .A (n_68_49), .B (n_62_52), .C1 (n_58_54), .C2 (n_52_57) );
AOI211_X1 g_74_46 (.ZN (n_74_46), .A (n_70_48), .B (n_64_51), .C1 (n_60_53), .C2 (n_54_56) );
AOI211_X1 g_76_45 (.ZN (n_76_45), .A (n_72_47), .B (n_66_50), .C1 (n_62_52), .C2 (n_56_55) );
AOI211_X1 g_78_44 (.ZN (n_78_44), .A (n_74_46), .B (n_68_49), .C1 (n_64_51), .C2 (n_58_54) );
AOI211_X1 g_80_43 (.ZN (n_80_43), .A (n_76_45), .B (n_70_48), .C1 (n_66_50), .C2 (n_60_53) );
AOI211_X1 g_82_42 (.ZN (n_82_42), .A (n_78_44), .B (n_72_47), .C1 (n_68_49), .C2 (n_62_52) );
AOI211_X1 g_84_41 (.ZN (n_84_41), .A (n_80_43), .B (n_74_46), .C1 (n_70_48), .C2 (n_64_51) );
AOI211_X1 g_86_40 (.ZN (n_86_40), .A (n_82_42), .B (n_76_45), .C1 (n_72_47), .C2 (n_66_50) );
AOI211_X1 g_88_39 (.ZN (n_88_39), .A (n_84_41), .B (n_78_44), .C1 (n_74_46), .C2 (n_68_49) );
AOI211_X1 g_90_38 (.ZN (n_90_38), .A (n_86_40), .B (n_80_43), .C1 (n_76_45), .C2 (n_70_48) );
AOI211_X1 g_92_37 (.ZN (n_92_37), .A (n_88_39), .B (n_82_42), .C1 (n_78_44), .C2 (n_72_47) );
AOI211_X1 g_94_36 (.ZN (n_94_36), .A (n_90_38), .B (n_84_41), .C1 (n_80_43), .C2 (n_74_46) );
AOI211_X1 g_96_35 (.ZN (n_96_35), .A (n_92_37), .B (n_86_40), .C1 (n_82_42), .C2 (n_76_45) );
AOI211_X1 g_98_34 (.ZN (n_98_34), .A (n_94_36), .B (n_88_39), .C1 (n_84_41), .C2 (n_78_44) );
AOI211_X1 g_100_33 (.ZN (n_100_33), .A (n_96_35), .B (n_90_38), .C1 (n_86_40), .C2 (n_80_43) );
AOI211_X1 g_102_32 (.ZN (n_102_32), .A (n_98_34), .B (n_92_37), .C1 (n_88_39), .C2 (n_82_42) );
AOI211_X1 g_104_31 (.ZN (n_104_31), .A (n_100_33), .B (n_94_36), .C1 (n_90_38), .C2 (n_84_41) );
AOI211_X1 g_106_30 (.ZN (n_106_30), .A (n_102_32), .B (n_96_35), .C1 (n_92_37), .C2 (n_86_40) );
AOI211_X1 g_108_29 (.ZN (n_108_29), .A (n_104_31), .B (n_98_34), .C1 (n_94_36), .C2 (n_88_39) );
AOI211_X1 g_110_28 (.ZN (n_110_28), .A (n_106_30), .B (n_100_33), .C1 (n_96_35), .C2 (n_90_38) );
AOI211_X1 g_112_27 (.ZN (n_112_27), .A (n_108_29), .B (n_102_32), .C1 (n_98_34), .C2 (n_92_37) );
AOI211_X1 g_114_26 (.ZN (n_114_26), .A (n_110_28), .B (n_104_31), .C1 (n_100_33), .C2 (n_94_36) );
AOI211_X1 g_116_25 (.ZN (n_116_25), .A (n_112_27), .B (n_106_30), .C1 (n_102_32), .C2 (n_96_35) );
AOI211_X1 g_118_24 (.ZN (n_118_24), .A (n_114_26), .B (n_108_29), .C1 (n_104_31), .C2 (n_98_34) );
AOI211_X1 g_120_23 (.ZN (n_120_23), .A (n_116_25), .B (n_110_28), .C1 (n_106_30), .C2 (n_100_33) );
AOI211_X1 g_122_22 (.ZN (n_122_22), .A (n_118_24), .B (n_112_27), .C1 (n_108_29), .C2 (n_102_32) );
AOI211_X1 g_121_24 (.ZN (n_121_24), .A (n_120_23), .B (n_114_26), .C1 (n_110_28), .C2 (n_104_31) );
AOI211_X1 g_123_23 (.ZN (n_123_23), .A (n_122_22), .B (n_116_25), .C1 (n_112_27), .C2 (n_106_30) );
AOI211_X1 g_125_22 (.ZN (n_125_22), .A (n_121_24), .B (n_118_24), .C1 (n_114_26), .C2 (n_108_29) );
AOI211_X1 g_127_21 (.ZN (n_127_21), .A (n_123_23), .B (n_120_23), .C1 (n_116_25), .C2 (n_110_28) );
AOI211_X1 g_129_22 (.ZN (n_129_22), .A (n_125_22), .B (n_122_22), .C1 (n_118_24), .C2 (n_112_27) );
AOI211_X1 g_130_20 (.ZN (n_130_20), .A (n_127_21), .B (n_121_24), .C1 (n_120_23), .C2 (n_114_26) );
AOI211_X1 g_132_19 (.ZN (n_132_19), .A (n_129_22), .B (n_123_23), .C1 (n_122_22), .C2 (n_116_25) );
AOI211_X1 g_134_18 (.ZN (n_134_18), .A (n_130_20), .B (n_125_22), .C1 (n_121_24), .C2 (n_118_24) );
AOI211_X1 g_136_17 (.ZN (n_136_17), .A (n_132_19), .B (n_127_21), .C1 (n_123_23), .C2 (n_120_23) );
AOI211_X1 g_138_18 (.ZN (n_138_18), .A (n_134_18), .B (n_129_22), .C1 (n_125_22), .C2 (n_122_22) );
AOI211_X1 g_136_19 (.ZN (n_136_19), .A (n_136_17), .B (n_130_20), .C1 (n_127_21), .C2 (n_121_24) );
AOI211_X1 g_134_20 (.ZN (n_134_20), .A (n_138_18), .B (n_132_19), .C1 (n_129_22), .C2 (n_123_23) );
AOI211_X1 g_135_18 (.ZN (n_135_18), .A (n_136_19), .B (n_134_18), .C1 (n_130_20), .C2 (n_125_22) );
AOI211_X1 g_133_19 (.ZN (n_133_19), .A (n_134_20), .B (n_136_17), .C1 (n_132_19), .C2 (n_127_21) );
AOI211_X1 g_131_20 (.ZN (n_131_20), .A (n_135_18), .B (n_138_18), .C1 (n_134_18), .C2 (n_129_22) );
AOI211_X1 g_129_21 (.ZN (n_129_21), .A (n_133_19), .B (n_136_19), .C1 (n_136_17), .C2 (n_130_20) );
AOI211_X1 g_127_20 (.ZN (n_127_20), .A (n_131_20), .B (n_134_20), .C1 (n_138_18), .C2 (n_132_19) );
AOI211_X1 g_125_21 (.ZN (n_125_21), .A (n_129_21), .B (n_135_18), .C1 (n_136_19), .C2 (n_134_18) );
AOI211_X1 g_123_22 (.ZN (n_123_22), .A (n_127_20), .B (n_133_19), .C1 (n_134_20), .C2 (n_136_17) );
AOI211_X1 g_121_23 (.ZN (n_121_23), .A (n_125_21), .B (n_131_20), .C1 (n_135_18), .C2 (n_138_18) );
AOI211_X1 g_119_24 (.ZN (n_119_24), .A (n_123_22), .B (n_129_21), .C1 (n_133_19), .C2 (n_136_19) );
AOI211_X1 g_117_25 (.ZN (n_117_25), .A (n_121_23), .B (n_127_20), .C1 (n_131_20), .C2 (n_134_20) );
AOI211_X1 g_115_26 (.ZN (n_115_26), .A (n_119_24), .B (n_125_21), .C1 (n_129_21), .C2 (n_135_18) );
AOI211_X1 g_113_27 (.ZN (n_113_27), .A (n_117_25), .B (n_123_22), .C1 (n_127_20), .C2 (n_133_19) );
AOI211_X1 g_111_28 (.ZN (n_111_28), .A (n_115_26), .B (n_121_23), .C1 (n_125_21), .C2 (n_131_20) );
AOI211_X1 g_113_29 (.ZN (n_113_29), .A (n_113_27), .B (n_119_24), .C1 (n_123_22), .C2 (n_129_21) );
AOI211_X1 g_115_28 (.ZN (n_115_28), .A (n_111_28), .B (n_117_25), .C1 (n_121_23), .C2 (n_127_20) );
AOI211_X1 g_117_27 (.ZN (n_117_27), .A (n_113_29), .B (n_115_26), .C1 (n_119_24), .C2 (n_125_21) );
AOI211_X1 g_119_26 (.ZN (n_119_26), .A (n_115_28), .B (n_113_27), .C1 (n_117_25), .C2 (n_123_22) );
AOI211_X1 g_120_24 (.ZN (n_120_24), .A (n_117_27), .B (n_111_28), .C1 (n_115_26), .C2 (n_121_23) );
AOI211_X1 g_122_23 (.ZN (n_122_23), .A (n_119_26), .B (n_113_29), .C1 (n_113_27), .C2 (n_119_24) );
AOI211_X1 g_124_22 (.ZN (n_124_22), .A (n_120_24), .B (n_115_28), .C1 (n_111_28), .C2 (n_117_25) );
AOI211_X1 g_126_21 (.ZN (n_126_21), .A (n_122_23), .B (n_117_27), .C1 (n_113_29), .C2 (n_115_26) );
AOI211_X1 g_128_22 (.ZN (n_128_22), .A (n_124_22), .B (n_119_26), .C1 (n_115_28), .C2 (n_113_27) );
AOI211_X1 g_126_23 (.ZN (n_126_23), .A (n_126_21), .B (n_120_24), .C1 (n_117_27), .C2 (n_111_28) );
AOI211_X1 g_124_24 (.ZN (n_124_24), .A (n_128_22), .B (n_122_23), .C1 (n_119_26), .C2 (n_113_29) );
AOI211_X1 g_122_25 (.ZN (n_122_25), .A (n_126_23), .B (n_124_22), .C1 (n_120_24), .C2 (n_115_28) );
AOI211_X1 g_120_26 (.ZN (n_120_26), .A (n_124_24), .B (n_126_21), .C1 (n_122_23), .C2 (n_117_27) );
AOI211_X1 g_118_27 (.ZN (n_118_27), .A (n_122_25), .B (n_128_22), .C1 (n_124_22), .C2 (n_119_26) );
AOI211_X1 g_119_25 (.ZN (n_119_25), .A (n_120_26), .B (n_126_23), .C1 (n_126_21), .C2 (n_120_24) );
AOI211_X1 g_117_26 (.ZN (n_117_26), .A (n_118_27), .B (n_124_24), .C1 (n_128_22), .C2 (n_122_23) );
AOI211_X1 g_115_27 (.ZN (n_115_27), .A (n_119_25), .B (n_122_25), .C1 (n_126_23), .C2 (n_124_22) );
AOI211_X1 g_113_28 (.ZN (n_113_28), .A (n_117_26), .B (n_120_26), .C1 (n_124_24), .C2 (n_126_21) );
AOI211_X1 g_111_29 (.ZN (n_111_29), .A (n_115_27), .B (n_118_27), .C1 (n_122_25), .C2 (n_128_22) );
AOI211_X1 g_109_28 (.ZN (n_109_28), .A (n_113_28), .B (n_119_25), .C1 (n_120_26), .C2 (n_126_23) );
AOI211_X1 g_107_29 (.ZN (n_107_29), .A (n_111_29), .B (n_117_26), .C1 (n_118_27), .C2 (n_124_24) );
AOI211_X1 g_105_30 (.ZN (n_105_30), .A (n_109_28), .B (n_115_27), .C1 (n_119_25), .C2 (n_122_25) );
AOI211_X1 g_103_31 (.ZN (n_103_31), .A (n_107_29), .B (n_113_28), .C1 (n_117_26), .C2 (n_120_26) );
AOI211_X1 g_101_32 (.ZN (n_101_32), .A (n_105_30), .B (n_111_29), .C1 (n_115_27), .C2 (n_118_27) );
AOI211_X1 g_99_33 (.ZN (n_99_33), .A (n_103_31), .B (n_109_28), .C1 (n_113_28), .C2 (n_119_25) );
AOI211_X1 g_97_34 (.ZN (n_97_34), .A (n_101_32), .B (n_107_29), .C1 (n_111_29), .C2 (n_117_26) );
AOI211_X1 g_95_35 (.ZN (n_95_35), .A (n_99_33), .B (n_105_30), .C1 (n_109_28), .C2 (n_115_27) );
AOI211_X1 g_93_36 (.ZN (n_93_36), .A (n_97_34), .B (n_103_31), .C1 (n_107_29), .C2 (n_113_28) );
AOI211_X1 g_91_37 (.ZN (n_91_37), .A (n_95_35), .B (n_101_32), .C1 (n_105_30), .C2 (n_111_29) );
AOI211_X1 g_89_38 (.ZN (n_89_38), .A (n_93_36), .B (n_99_33), .C1 (n_103_31), .C2 (n_109_28) );
AOI211_X1 g_87_39 (.ZN (n_87_39), .A (n_91_37), .B (n_97_34), .C1 (n_101_32), .C2 (n_107_29) );
AOI211_X1 g_85_40 (.ZN (n_85_40), .A (n_89_38), .B (n_95_35), .C1 (n_99_33), .C2 (n_105_30) );
AOI211_X1 g_83_41 (.ZN (n_83_41), .A (n_87_39), .B (n_93_36), .C1 (n_97_34), .C2 (n_103_31) );
AOI211_X1 g_81_42 (.ZN (n_81_42), .A (n_85_40), .B (n_91_37), .C1 (n_95_35), .C2 (n_101_32) );
AOI211_X1 g_79_43 (.ZN (n_79_43), .A (n_83_41), .B (n_89_38), .C1 (n_93_36), .C2 (n_99_33) );
AOI211_X1 g_77_44 (.ZN (n_77_44), .A (n_81_42), .B (n_87_39), .C1 (n_91_37), .C2 (n_97_34) );
AOI211_X1 g_75_45 (.ZN (n_75_45), .A (n_79_43), .B (n_85_40), .C1 (n_89_38), .C2 (n_95_35) );
AOI211_X1 g_73_46 (.ZN (n_73_46), .A (n_77_44), .B (n_83_41), .C1 (n_87_39), .C2 (n_93_36) );
AOI211_X1 g_71_47 (.ZN (n_71_47), .A (n_75_45), .B (n_81_42), .C1 (n_85_40), .C2 (n_91_37) );
AOI211_X1 g_70_49 (.ZN (n_70_49), .A (n_73_46), .B (n_79_43), .C1 (n_83_41), .C2 (n_89_38) );
AOI211_X1 g_68_50 (.ZN (n_68_50), .A (n_71_47), .B (n_77_44), .C1 (n_81_42), .C2 (n_87_39) );
AOI211_X1 g_67_52 (.ZN (n_67_52), .A (n_70_49), .B (n_75_45), .C1 (n_79_43), .C2 (n_85_40) );
AOI211_X1 g_69_51 (.ZN (n_69_51), .A (n_68_50), .B (n_73_46), .C1 (n_77_44), .C2 (n_83_41) );
AOI211_X1 g_71_50 (.ZN (n_71_50), .A (n_67_52), .B (n_71_47), .C1 (n_75_45), .C2 (n_81_42) );
AOI211_X1 g_72_48 (.ZN (n_72_48), .A (n_69_51), .B (n_70_49), .C1 (n_73_46), .C2 (n_79_43) );
AOI211_X1 g_74_47 (.ZN (n_74_47), .A (n_71_50), .B (n_68_50), .C1 (n_71_47), .C2 (n_77_44) );
AOI211_X1 g_76_46 (.ZN (n_76_46), .A (n_72_48), .B (n_67_52), .C1 (n_70_49), .C2 (n_75_45) );
AOI211_X1 g_78_45 (.ZN (n_78_45), .A (n_74_47), .B (n_69_51), .C1 (n_68_50), .C2 (n_73_46) );
AOI211_X1 g_80_44 (.ZN (n_80_44), .A (n_76_46), .B (n_71_50), .C1 (n_67_52), .C2 (n_71_47) );
AOI211_X1 g_82_43 (.ZN (n_82_43), .A (n_78_45), .B (n_72_48), .C1 (n_69_51), .C2 (n_70_49) );
AOI211_X1 g_84_42 (.ZN (n_84_42), .A (n_80_44), .B (n_74_47), .C1 (n_71_50), .C2 (n_68_50) );
AOI211_X1 g_86_41 (.ZN (n_86_41), .A (n_82_43), .B (n_76_46), .C1 (n_72_48), .C2 (n_67_52) );
AOI211_X1 g_88_40 (.ZN (n_88_40), .A (n_84_42), .B (n_78_45), .C1 (n_74_47), .C2 (n_69_51) );
AOI211_X1 g_90_39 (.ZN (n_90_39), .A (n_86_41), .B (n_80_44), .C1 (n_76_46), .C2 (n_71_50) );
AOI211_X1 g_92_38 (.ZN (n_92_38), .A (n_88_40), .B (n_82_43), .C1 (n_78_45), .C2 (n_72_48) );
AOI211_X1 g_94_37 (.ZN (n_94_37), .A (n_90_39), .B (n_84_42), .C1 (n_80_44), .C2 (n_74_47) );
AOI211_X1 g_96_36 (.ZN (n_96_36), .A (n_92_38), .B (n_86_41), .C1 (n_82_43), .C2 (n_76_46) );
AOI211_X1 g_98_35 (.ZN (n_98_35), .A (n_94_37), .B (n_88_40), .C1 (n_84_42), .C2 (n_78_45) );
AOI211_X1 g_100_34 (.ZN (n_100_34), .A (n_96_36), .B (n_90_39), .C1 (n_86_41), .C2 (n_80_44) );
AOI211_X1 g_102_33 (.ZN (n_102_33), .A (n_98_35), .B (n_92_38), .C1 (n_88_40), .C2 (n_82_43) );
AOI211_X1 g_104_32 (.ZN (n_104_32), .A (n_100_34), .B (n_94_37), .C1 (n_90_39), .C2 (n_84_42) );
AOI211_X1 g_106_31 (.ZN (n_106_31), .A (n_102_33), .B (n_96_36), .C1 (n_92_38), .C2 (n_86_41) );
AOI211_X1 g_108_30 (.ZN (n_108_30), .A (n_104_32), .B (n_98_35), .C1 (n_94_37), .C2 (n_88_40) );
AOI211_X1 g_107_32 (.ZN (n_107_32), .A (n_106_31), .B (n_100_34), .C1 (n_96_36), .C2 (n_90_39) );
AOI211_X1 g_109_31 (.ZN (n_109_31), .A (n_108_30), .B (n_102_33), .C1 (n_98_35), .C2 (n_92_38) );
AOI211_X1 g_111_30 (.ZN (n_111_30), .A (n_107_32), .B (n_104_32), .C1 (n_100_34), .C2 (n_94_37) );
AOI211_X1 g_110_32 (.ZN (n_110_32), .A (n_109_31), .B (n_106_31), .C1 (n_102_33), .C2 (n_96_36) );
AOI211_X1 g_109_30 (.ZN (n_109_30), .A (n_111_30), .B (n_108_30), .C1 (n_104_32), .C2 (n_98_35) );
AOI211_X1 g_107_31 (.ZN (n_107_31), .A (n_110_32), .B (n_107_32), .C1 (n_106_31), .C2 (n_100_34) );
AOI211_X1 g_105_32 (.ZN (n_105_32), .A (n_109_30), .B (n_109_31), .C1 (n_108_30), .C2 (n_102_33) );
AOI211_X1 g_103_33 (.ZN (n_103_33), .A (n_107_31), .B (n_111_30), .C1 (n_107_32), .C2 (n_104_32) );
AOI211_X1 g_101_34 (.ZN (n_101_34), .A (n_105_32), .B (n_110_32), .C1 (n_109_31), .C2 (n_106_31) );
AOI211_X1 g_99_35 (.ZN (n_99_35), .A (n_103_33), .B (n_109_30), .C1 (n_111_30), .C2 (n_108_30) );
AOI211_X1 g_97_36 (.ZN (n_97_36), .A (n_101_34), .B (n_107_31), .C1 (n_110_32), .C2 (n_107_32) );
AOI211_X1 g_95_37 (.ZN (n_95_37), .A (n_99_35), .B (n_105_32), .C1 (n_109_30), .C2 (n_109_31) );
AOI211_X1 g_93_38 (.ZN (n_93_38), .A (n_97_36), .B (n_103_33), .C1 (n_107_31), .C2 (n_111_30) );
AOI211_X1 g_91_39 (.ZN (n_91_39), .A (n_95_37), .B (n_101_34), .C1 (n_105_32), .C2 (n_110_32) );
AOI211_X1 g_89_40 (.ZN (n_89_40), .A (n_93_38), .B (n_99_35), .C1 (n_103_33), .C2 (n_109_30) );
AOI211_X1 g_87_41 (.ZN (n_87_41), .A (n_91_39), .B (n_97_36), .C1 (n_101_34), .C2 (n_107_31) );
AOI211_X1 g_85_42 (.ZN (n_85_42), .A (n_89_40), .B (n_95_37), .C1 (n_99_35), .C2 (n_105_32) );
AOI211_X1 g_83_43 (.ZN (n_83_43), .A (n_87_41), .B (n_93_38), .C1 (n_97_36), .C2 (n_103_33) );
AOI211_X1 g_81_44 (.ZN (n_81_44), .A (n_85_42), .B (n_91_39), .C1 (n_95_37), .C2 (n_101_34) );
AOI211_X1 g_79_45 (.ZN (n_79_45), .A (n_83_43), .B (n_89_40), .C1 (n_93_38), .C2 (n_99_35) );
AOI211_X1 g_77_46 (.ZN (n_77_46), .A (n_81_44), .B (n_87_41), .C1 (n_91_39), .C2 (n_97_36) );
AOI211_X1 g_75_47 (.ZN (n_75_47), .A (n_79_45), .B (n_85_42), .C1 (n_89_40), .C2 (n_95_37) );
AOI211_X1 g_73_48 (.ZN (n_73_48), .A (n_77_46), .B (n_83_43), .C1 (n_87_41), .C2 (n_93_38) );
AOI211_X1 g_71_49 (.ZN (n_71_49), .A (n_75_47), .B (n_81_44), .C1 (n_85_42), .C2 (n_91_39) );
AOI211_X1 g_69_50 (.ZN (n_69_50), .A (n_73_48), .B (n_79_45), .C1 (n_83_43), .C2 (n_89_40) );
AOI211_X1 g_67_51 (.ZN (n_67_51), .A (n_71_49), .B (n_77_46), .C1 (n_81_44), .C2 (n_87_41) );
AOI211_X1 g_65_52 (.ZN (n_65_52), .A (n_69_50), .B (n_75_47), .C1 (n_79_45), .C2 (n_85_42) );
AOI211_X1 g_63_53 (.ZN (n_63_53), .A (n_67_51), .B (n_73_48), .C1 (n_77_46), .C2 (n_83_43) );
AOI211_X1 g_61_54 (.ZN (n_61_54), .A (n_65_52), .B (n_71_49), .C1 (n_75_47), .C2 (n_81_44) );
AOI211_X1 g_59_55 (.ZN (n_59_55), .A (n_63_53), .B (n_69_50), .C1 (n_73_48), .C2 (n_79_45) );
AOI211_X1 g_57_56 (.ZN (n_57_56), .A (n_61_54), .B (n_67_51), .C1 (n_71_49), .C2 (n_77_46) );
AOI211_X1 g_55_57 (.ZN (n_55_57), .A (n_59_55), .B (n_65_52), .C1 (n_69_50), .C2 (n_75_47) );
AOI211_X1 g_53_58 (.ZN (n_53_58), .A (n_57_56), .B (n_63_53), .C1 (n_67_51), .C2 (n_73_48) );
AOI211_X1 g_51_59 (.ZN (n_51_59), .A (n_55_57), .B (n_61_54), .C1 (n_65_52), .C2 (n_71_49) );
AOI211_X1 g_49_60 (.ZN (n_49_60), .A (n_53_58), .B (n_59_55), .C1 (n_63_53), .C2 (n_69_50) );
AOI211_X1 g_47_61 (.ZN (n_47_61), .A (n_51_59), .B (n_57_56), .C1 (n_61_54), .C2 (n_67_51) );
AOI211_X1 g_45_62 (.ZN (n_45_62), .A (n_49_60), .B (n_55_57), .C1 (n_59_55), .C2 (n_65_52) );
AOI211_X1 g_43_63 (.ZN (n_43_63), .A (n_47_61), .B (n_53_58), .C1 (n_57_56), .C2 (n_63_53) );
AOI211_X1 g_41_64 (.ZN (n_41_64), .A (n_45_62), .B (n_51_59), .C1 (n_55_57), .C2 (n_61_54) );
AOI211_X1 g_39_65 (.ZN (n_39_65), .A (n_43_63), .B (n_49_60), .C1 (n_53_58), .C2 (n_59_55) );
AOI211_X1 g_37_66 (.ZN (n_37_66), .A (n_41_64), .B (n_47_61), .C1 (n_51_59), .C2 (n_57_56) );
AOI211_X1 g_35_67 (.ZN (n_35_67), .A (n_39_65), .B (n_45_62), .C1 (n_49_60), .C2 (n_55_57) );
AOI211_X1 g_33_68 (.ZN (n_33_68), .A (n_37_66), .B (n_43_63), .C1 (n_47_61), .C2 (n_53_58) );
AOI211_X1 g_31_69 (.ZN (n_31_69), .A (n_35_67), .B (n_41_64), .C1 (n_45_62), .C2 (n_51_59) );
AOI211_X1 g_29_70 (.ZN (n_29_70), .A (n_33_68), .B (n_39_65), .C1 (n_43_63), .C2 (n_49_60) );
AOI211_X1 g_27_71 (.ZN (n_27_71), .A (n_31_69), .B (n_37_66), .C1 (n_41_64), .C2 (n_47_61) );
AOI211_X1 g_25_72 (.ZN (n_25_72), .A (n_29_70), .B (n_35_67), .C1 (n_39_65), .C2 (n_45_62) );
AOI211_X1 g_23_73 (.ZN (n_23_73), .A (n_27_71), .B (n_33_68), .C1 (n_37_66), .C2 (n_43_63) );
AOI211_X1 g_21_74 (.ZN (n_21_74), .A (n_25_72), .B (n_31_69), .C1 (n_35_67), .C2 (n_41_64) );
AOI211_X1 g_19_75 (.ZN (n_19_75), .A (n_23_73), .B (n_29_70), .C1 (n_33_68), .C2 (n_39_65) );
AOI211_X1 g_17_76 (.ZN (n_17_76), .A (n_21_74), .B (n_27_71), .C1 (n_31_69), .C2 (n_37_66) );
AOI211_X1 g_15_77 (.ZN (n_15_77), .A (n_19_75), .B (n_25_72), .C1 (n_29_70), .C2 (n_35_67) );
AOI211_X1 g_13_78 (.ZN (n_13_78), .A (n_17_76), .B (n_23_73), .C1 (n_27_71), .C2 (n_33_68) );
AOI211_X1 g_11_79 (.ZN (n_11_79), .A (n_15_77), .B (n_21_74), .C1 (n_25_72), .C2 (n_31_69) );
AOI211_X1 g_9_80 (.ZN (n_9_80), .A (n_13_78), .B (n_19_75), .C1 (n_23_73), .C2 (n_29_70) );
AOI211_X1 g_8_82 (.ZN (n_8_82), .A (n_11_79), .B (n_17_76), .C1 (n_21_74), .C2 (n_27_71) );
AOI211_X1 g_10_81 (.ZN (n_10_81), .A (n_9_80), .B (n_15_77), .C1 (n_19_75), .C2 (n_25_72) );
AOI211_X1 g_12_80 (.ZN (n_12_80), .A (n_8_82), .B (n_13_78), .C1 (n_17_76), .C2 (n_23_73) );
AOI211_X1 g_14_79 (.ZN (n_14_79), .A (n_10_81), .B (n_11_79), .C1 (n_15_77), .C2 (n_21_74) );
AOI211_X1 g_16_78 (.ZN (n_16_78), .A (n_12_80), .B (n_9_80), .C1 (n_13_78), .C2 (n_19_75) );
AOI211_X1 g_15_76 (.ZN (n_15_76), .A (n_14_79), .B (n_8_82), .C1 (n_11_79), .C2 (n_17_76) );
AOI211_X1 g_17_75 (.ZN (n_17_75), .A (n_16_78), .B (n_10_81), .C1 (n_9_80), .C2 (n_15_77) );
AOI211_X1 g_19_74 (.ZN (n_19_74), .A (n_15_76), .B (n_12_80), .C1 (n_8_82), .C2 (n_13_78) );
AOI211_X1 g_21_73 (.ZN (n_21_73), .A (n_17_75), .B (n_14_79), .C1 (n_10_81), .C2 (n_11_79) );
AOI211_X1 g_23_72 (.ZN (n_23_72), .A (n_19_74), .B (n_16_78), .C1 (n_12_80), .C2 (n_9_80) );
AOI211_X1 g_25_71 (.ZN (n_25_71), .A (n_21_73), .B (n_15_76), .C1 (n_14_79), .C2 (n_8_82) );
AOI211_X1 g_27_70 (.ZN (n_27_70), .A (n_23_72), .B (n_17_75), .C1 (n_16_78), .C2 (n_10_81) );
AOI211_X1 g_26_72 (.ZN (n_26_72), .A (n_25_71), .B (n_19_74), .C1 (n_15_76), .C2 (n_12_80) );
AOI211_X1 g_28_71 (.ZN (n_28_71), .A (n_27_70), .B (n_21_73), .C1 (n_17_75), .C2 (n_14_79) );
AOI211_X1 g_30_70 (.ZN (n_30_70), .A (n_26_72), .B (n_23_72), .C1 (n_19_74), .C2 (n_16_78) );
AOI211_X1 g_32_69 (.ZN (n_32_69), .A (n_28_71), .B (n_25_71), .C1 (n_21_73), .C2 (n_15_76) );
AOI211_X1 g_34_68 (.ZN (n_34_68), .A (n_30_70), .B (n_27_70), .C1 (n_23_72), .C2 (n_17_75) );
AOI211_X1 g_36_67 (.ZN (n_36_67), .A (n_32_69), .B (n_26_72), .C1 (n_25_71), .C2 (n_19_74) );
AOI211_X1 g_38_66 (.ZN (n_38_66), .A (n_34_68), .B (n_28_71), .C1 (n_27_70), .C2 (n_21_73) );
AOI211_X1 g_40_65 (.ZN (n_40_65), .A (n_36_67), .B (n_30_70), .C1 (n_26_72), .C2 (n_23_72) );
AOI211_X1 g_42_64 (.ZN (n_42_64), .A (n_38_66), .B (n_32_69), .C1 (n_28_71), .C2 (n_25_71) );
AOI211_X1 g_44_63 (.ZN (n_44_63), .A (n_40_65), .B (n_34_68), .C1 (n_30_70), .C2 (n_27_70) );
AOI211_X1 g_46_62 (.ZN (n_46_62), .A (n_42_64), .B (n_36_67), .C1 (n_32_69), .C2 (n_26_72) );
AOI211_X1 g_48_61 (.ZN (n_48_61), .A (n_44_63), .B (n_38_66), .C1 (n_34_68), .C2 (n_28_71) );
AOI211_X1 g_50_60 (.ZN (n_50_60), .A (n_46_62), .B (n_40_65), .C1 (n_36_67), .C2 (n_30_70) );
AOI211_X1 g_51_58 (.ZN (n_51_58), .A (n_48_61), .B (n_42_64), .C1 (n_38_66), .C2 (n_32_69) );
AOI211_X1 g_53_57 (.ZN (n_53_57), .A (n_50_60), .B (n_44_63), .C1 (n_40_65), .C2 (n_34_68) );
AOI211_X1 g_55_56 (.ZN (n_55_56), .A (n_51_58), .B (n_46_62), .C1 (n_42_64), .C2 (n_36_67) );
AOI211_X1 g_57_55 (.ZN (n_57_55), .A (n_53_57), .B (n_48_61), .C1 (n_44_63), .C2 (n_38_66) );
AOI211_X1 g_59_54 (.ZN (n_59_54), .A (n_55_56), .B (n_50_60), .C1 (n_46_62), .C2 (n_40_65) );
AOI211_X1 g_61_53 (.ZN (n_61_53), .A (n_57_55), .B (n_51_58), .C1 (n_48_61), .C2 (n_42_64) );
AOI211_X1 g_63_52 (.ZN (n_63_52), .A (n_59_54), .B (n_53_57), .C1 (n_50_60), .C2 (n_44_63) );
AOI211_X1 g_65_53 (.ZN (n_65_53), .A (n_61_53), .B (n_55_56), .C1 (n_51_58), .C2 (n_46_62) );
AOI211_X1 g_63_54 (.ZN (n_63_54), .A (n_63_52), .B (n_57_55), .C1 (n_53_57), .C2 (n_48_61) );
AOI211_X1 g_61_55 (.ZN (n_61_55), .A (n_65_53), .B (n_59_54), .C1 (n_55_56), .C2 (n_50_60) );
AOI211_X1 g_59_56 (.ZN (n_59_56), .A (n_63_54), .B (n_61_53), .C1 (n_57_55), .C2 (n_51_58) );
AOI211_X1 g_57_57 (.ZN (n_57_57), .A (n_61_55), .B (n_63_52), .C1 (n_59_54), .C2 (n_53_57) );
AOI211_X1 g_55_58 (.ZN (n_55_58), .A (n_59_56), .B (n_65_53), .C1 (n_61_53), .C2 (n_55_56) );
AOI211_X1 g_53_59 (.ZN (n_53_59), .A (n_57_57), .B (n_63_54), .C1 (n_63_52), .C2 (n_57_55) );
AOI211_X1 g_51_60 (.ZN (n_51_60), .A (n_55_58), .B (n_61_55), .C1 (n_65_53), .C2 (n_59_54) );
AOI211_X1 g_49_61 (.ZN (n_49_61), .A (n_53_59), .B (n_59_56), .C1 (n_63_54), .C2 (n_61_53) );
AOI211_X1 g_47_62 (.ZN (n_47_62), .A (n_51_60), .B (n_57_57), .C1 (n_61_55), .C2 (n_63_52) );
AOI211_X1 g_48_60 (.ZN (n_48_60), .A (n_49_61), .B (n_55_58), .C1 (n_59_56), .C2 (n_65_53) );
AOI211_X1 g_46_61 (.ZN (n_46_61), .A (n_47_62), .B (n_53_59), .C1 (n_57_57), .C2 (n_63_54) );
AOI211_X1 g_44_62 (.ZN (n_44_62), .A (n_48_60), .B (n_51_60), .C1 (n_55_58), .C2 (n_61_55) );
AOI211_X1 g_42_63 (.ZN (n_42_63), .A (n_46_61), .B (n_49_61), .C1 (n_53_59), .C2 (n_59_56) );
AOI211_X1 g_40_64 (.ZN (n_40_64), .A (n_44_62), .B (n_47_62), .C1 (n_51_60), .C2 (n_57_57) );
AOI211_X1 g_38_65 (.ZN (n_38_65), .A (n_42_63), .B (n_48_60), .C1 (n_49_61), .C2 (n_55_58) );
AOI211_X1 g_36_66 (.ZN (n_36_66), .A (n_40_64), .B (n_46_61), .C1 (n_47_62), .C2 (n_53_59) );
AOI211_X1 g_34_67 (.ZN (n_34_67), .A (n_38_65), .B (n_44_62), .C1 (n_48_60), .C2 (n_51_60) );
AOI211_X1 g_32_68 (.ZN (n_32_68), .A (n_36_66), .B (n_42_63), .C1 (n_46_61), .C2 (n_49_61) );
AOI211_X1 g_30_69 (.ZN (n_30_69), .A (n_34_67), .B (n_40_64), .C1 (n_44_62), .C2 (n_47_62) );
AOI211_X1 g_29_71 (.ZN (n_29_71), .A (n_32_68), .B (n_38_65), .C1 (n_42_63), .C2 (n_48_60) );
AOI211_X1 g_31_70 (.ZN (n_31_70), .A (n_30_69), .B (n_36_66), .C1 (n_40_64), .C2 (n_46_61) );
AOI211_X1 g_33_69 (.ZN (n_33_69), .A (n_29_71), .B (n_34_67), .C1 (n_38_65), .C2 (n_44_62) );
AOI211_X1 g_35_68 (.ZN (n_35_68), .A (n_31_70), .B (n_32_68), .C1 (n_36_66), .C2 (n_42_63) );
AOI211_X1 g_37_67 (.ZN (n_37_67), .A (n_33_69), .B (n_30_69), .C1 (n_34_67), .C2 (n_40_64) );
AOI211_X1 g_39_66 (.ZN (n_39_66), .A (n_35_68), .B (n_29_71), .C1 (n_32_68), .C2 (n_38_65) );
AOI211_X1 g_41_65 (.ZN (n_41_65), .A (n_37_67), .B (n_31_70), .C1 (n_30_69), .C2 (n_36_66) );
AOI211_X1 g_43_64 (.ZN (n_43_64), .A (n_39_66), .B (n_33_69), .C1 (n_29_71), .C2 (n_34_67) );
AOI211_X1 g_45_63 (.ZN (n_45_63), .A (n_41_65), .B (n_35_68), .C1 (n_31_70), .C2 (n_32_68) );
AOI211_X1 g_44_65 (.ZN (n_44_65), .A (n_43_64), .B (n_37_67), .C1 (n_33_69), .C2 (n_30_69) );
AOI211_X1 g_46_64 (.ZN (n_46_64), .A (n_45_63), .B (n_39_66), .C1 (n_35_68), .C2 (n_29_71) );
AOI211_X1 g_48_63 (.ZN (n_48_63), .A (n_44_65), .B (n_41_65), .C1 (n_37_67), .C2 (n_31_70) );
AOI211_X1 g_50_62 (.ZN (n_50_62), .A (n_46_64), .B (n_43_64), .C1 (n_39_66), .C2 (n_33_69) );
AOI211_X1 g_52_61 (.ZN (n_52_61), .A (n_48_63), .B (n_45_63), .C1 (n_41_65), .C2 (n_35_68) );
AOI211_X1 g_54_60 (.ZN (n_54_60), .A (n_50_62), .B (n_44_65), .C1 (n_43_64), .C2 (n_37_67) );
AOI211_X1 g_52_59 (.ZN (n_52_59), .A (n_52_61), .B (n_46_64), .C1 (n_45_63), .C2 (n_39_66) );
AOI211_X1 g_54_58 (.ZN (n_54_58), .A (n_54_60), .B (n_48_63), .C1 (n_44_65), .C2 (n_41_65) );
AOI211_X1 g_56_57 (.ZN (n_56_57), .A (n_52_59), .B (n_50_62), .C1 (n_46_64), .C2 (n_43_64) );
AOI211_X1 g_58_56 (.ZN (n_58_56), .A (n_54_58), .B (n_52_61), .C1 (n_48_63), .C2 (n_45_63) );
AOI211_X1 g_60_55 (.ZN (n_60_55), .A (n_56_57), .B (n_54_60), .C1 (n_50_62), .C2 (n_44_65) );
AOI211_X1 g_62_54 (.ZN (n_62_54), .A (n_58_56), .B (n_52_59), .C1 (n_52_61), .C2 (n_46_64) );
AOI211_X1 g_64_53 (.ZN (n_64_53), .A (n_60_55), .B (n_54_58), .C1 (n_54_60), .C2 (n_48_63) );
AOI211_X1 g_66_52 (.ZN (n_66_52), .A (n_62_54), .B (n_56_57), .C1 (n_52_59), .C2 (n_50_62) );
AOI211_X1 g_68_51 (.ZN (n_68_51), .A (n_64_53), .B (n_58_56), .C1 (n_54_58), .C2 (n_52_61) );
AOI211_X1 g_70_50 (.ZN (n_70_50), .A (n_66_52), .B (n_60_55), .C1 (n_56_57), .C2 (n_54_60) );
AOI211_X1 g_72_49 (.ZN (n_72_49), .A (n_68_51), .B (n_62_54), .C1 (n_58_56), .C2 (n_52_59) );
AOI211_X1 g_74_48 (.ZN (n_74_48), .A (n_70_50), .B (n_64_53), .C1 (n_60_55), .C2 (n_54_58) );
AOI211_X1 g_76_47 (.ZN (n_76_47), .A (n_72_49), .B (n_66_52), .C1 (n_62_54), .C2 (n_56_57) );
AOI211_X1 g_78_46 (.ZN (n_78_46), .A (n_74_48), .B (n_68_51), .C1 (n_64_53), .C2 (n_58_56) );
AOI211_X1 g_80_45 (.ZN (n_80_45), .A (n_76_47), .B (n_70_50), .C1 (n_66_52), .C2 (n_60_55) );
AOI211_X1 g_82_44 (.ZN (n_82_44), .A (n_78_46), .B (n_72_49), .C1 (n_68_51), .C2 (n_62_54) );
AOI211_X1 g_84_43 (.ZN (n_84_43), .A (n_80_45), .B (n_74_48), .C1 (n_70_50), .C2 (n_64_53) );
AOI211_X1 g_86_42 (.ZN (n_86_42), .A (n_82_44), .B (n_76_47), .C1 (n_72_49), .C2 (n_66_52) );
AOI211_X1 g_88_41 (.ZN (n_88_41), .A (n_84_43), .B (n_78_46), .C1 (n_74_48), .C2 (n_68_51) );
AOI211_X1 g_90_40 (.ZN (n_90_40), .A (n_86_42), .B (n_80_45), .C1 (n_76_47), .C2 (n_70_50) );
AOI211_X1 g_92_39 (.ZN (n_92_39), .A (n_88_41), .B (n_82_44), .C1 (n_78_46), .C2 (n_72_49) );
AOI211_X1 g_94_38 (.ZN (n_94_38), .A (n_90_40), .B (n_84_43), .C1 (n_80_45), .C2 (n_74_48) );
AOI211_X1 g_96_37 (.ZN (n_96_37), .A (n_92_39), .B (n_86_42), .C1 (n_82_44), .C2 (n_76_47) );
AOI211_X1 g_98_36 (.ZN (n_98_36), .A (n_94_38), .B (n_88_41), .C1 (n_84_43), .C2 (n_78_46) );
AOI211_X1 g_100_35 (.ZN (n_100_35), .A (n_96_37), .B (n_90_40), .C1 (n_86_42), .C2 (n_80_45) );
AOI211_X1 g_102_34 (.ZN (n_102_34), .A (n_98_36), .B (n_92_39), .C1 (n_88_41), .C2 (n_82_44) );
AOI211_X1 g_104_33 (.ZN (n_104_33), .A (n_100_35), .B (n_94_38), .C1 (n_90_40), .C2 (n_84_43) );
AOI211_X1 g_106_32 (.ZN (n_106_32), .A (n_102_34), .B (n_96_37), .C1 (n_92_39), .C2 (n_86_42) );
AOI211_X1 g_108_31 (.ZN (n_108_31), .A (n_104_33), .B (n_98_36), .C1 (n_94_38), .C2 (n_88_41) );
AOI211_X1 g_110_30 (.ZN (n_110_30), .A (n_106_32), .B (n_100_35), .C1 (n_96_37), .C2 (n_90_40) );
AOI211_X1 g_112_29 (.ZN (n_112_29), .A (n_108_31), .B (n_102_34), .C1 (n_98_36), .C2 (n_92_39) );
AOI211_X1 g_114_28 (.ZN (n_114_28), .A (n_110_30), .B (n_104_33), .C1 (n_100_35), .C2 (n_94_38) );
AOI211_X1 g_116_27 (.ZN (n_116_27), .A (n_112_29), .B (n_106_32), .C1 (n_102_34), .C2 (n_96_37) );
AOI211_X1 g_118_26 (.ZN (n_118_26), .A (n_114_28), .B (n_108_31), .C1 (n_104_33), .C2 (n_98_36) );
AOI211_X1 g_120_25 (.ZN (n_120_25), .A (n_116_27), .B (n_110_30), .C1 (n_106_32), .C2 (n_100_35) );
AOI211_X1 g_122_24 (.ZN (n_122_24), .A (n_118_26), .B (n_112_29), .C1 (n_108_31), .C2 (n_102_34) );
AOI211_X1 g_124_23 (.ZN (n_124_23), .A (n_120_25), .B (n_114_28), .C1 (n_110_30), .C2 (n_104_33) );
AOI211_X1 g_126_22 (.ZN (n_126_22), .A (n_122_24), .B (n_116_27), .C1 (n_112_29), .C2 (n_106_32) );
AOI211_X1 g_128_21 (.ZN (n_128_21), .A (n_124_23), .B (n_118_26), .C1 (n_114_28), .C2 (n_108_31) );
AOI211_X1 g_127_23 (.ZN (n_127_23), .A (n_126_22), .B (n_120_25), .C1 (n_116_27), .C2 (n_110_30) );
AOI211_X1 g_125_24 (.ZN (n_125_24), .A (n_128_21), .B (n_122_24), .C1 (n_118_26), .C2 (n_112_29) );
AOI211_X1 g_123_25 (.ZN (n_123_25), .A (n_127_23), .B (n_124_23), .C1 (n_120_25), .C2 (n_114_28) );
AOI211_X1 g_121_26 (.ZN (n_121_26), .A (n_125_24), .B (n_126_22), .C1 (n_122_24), .C2 (n_116_27) );
AOI211_X1 g_119_27 (.ZN (n_119_27), .A (n_123_25), .B (n_128_21), .C1 (n_124_23), .C2 (n_118_26) );
AOI211_X1 g_117_28 (.ZN (n_117_28), .A (n_121_26), .B (n_127_23), .C1 (n_126_22), .C2 (n_120_25) );
AOI211_X1 g_115_29 (.ZN (n_115_29), .A (n_119_27), .B (n_125_24), .C1 (n_128_21), .C2 (n_122_24) );
AOI211_X1 g_113_30 (.ZN (n_113_30), .A (n_117_28), .B (n_123_25), .C1 (n_127_23), .C2 (n_124_23) );
AOI211_X1 g_111_31 (.ZN (n_111_31), .A (n_115_29), .B (n_121_26), .C1 (n_125_24), .C2 (n_126_22) );
AOI211_X1 g_109_32 (.ZN (n_109_32), .A (n_113_30), .B (n_119_27), .C1 (n_123_25), .C2 (n_128_21) );
AOI211_X1 g_107_33 (.ZN (n_107_33), .A (n_111_31), .B (n_117_28), .C1 (n_121_26), .C2 (n_127_23) );
AOI211_X1 g_105_34 (.ZN (n_105_34), .A (n_109_32), .B (n_115_29), .C1 (n_119_27), .C2 (n_125_24) );
AOI211_X1 g_103_35 (.ZN (n_103_35), .A (n_107_33), .B (n_113_30), .C1 (n_117_28), .C2 (n_123_25) );
AOI211_X1 g_101_36 (.ZN (n_101_36), .A (n_105_34), .B (n_111_31), .C1 (n_115_29), .C2 (n_121_26) );
AOI211_X1 g_99_37 (.ZN (n_99_37), .A (n_103_35), .B (n_109_32), .C1 (n_113_30), .C2 (n_119_27) );
AOI211_X1 g_97_38 (.ZN (n_97_38), .A (n_101_36), .B (n_107_33), .C1 (n_111_31), .C2 (n_117_28) );
AOI211_X1 g_95_39 (.ZN (n_95_39), .A (n_99_37), .B (n_105_34), .C1 (n_109_32), .C2 (n_115_29) );
AOI211_X1 g_93_40 (.ZN (n_93_40), .A (n_97_38), .B (n_103_35), .C1 (n_107_33), .C2 (n_113_30) );
AOI211_X1 g_91_41 (.ZN (n_91_41), .A (n_95_39), .B (n_101_36), .C1 (n_105_34), .C2 (n_111_31) );
AOI211_X1 g_89_42 (.ZN (n_89_42), .A (n_93_40), .B (n_99_37), .C1 (n_103_35), .C2 (n_109_32) );
AOI211_X1 g_87_43 (.ZN (n_87_43), .A (n_91_41), .B (n_97_38), .C1 (n_101_36), .C2 (n_107_33) );
AOI211_X1 g_85_44 (.ZN (n_85_44), .A (n_89_42), .B (n_95_39), .C1 (n_99_37), .C2 (n_105_34) );
AOI211_X1 g_83_45 (.ZN (n_83_45), .A (n_87_43), .B (n_93_40), .C1 (n_97_38), .C2 (n_103_35) );
AOI211_X1 g_81_46 (.ZN (n_81_46), .A (n_85_44), .B (n_91_41), .C1 (n_95_39), .C2 (n_101_36) );
AOI211_X1 g_79_47 (.ZN (n_79_47), .A (n_83_45), .B (n_89_42), .C1 (n_93_40), .C2 (n_99_37) );
AOI211_X1 g_77_48 (.ZN (n_77_48), .A (n_81_46), .B (n_87_43), .C1 (n_91_41), .C2 (n_97_38) );
AOI211_X1 g_75_49 (.ZN (n_75_49), .A (n_79_47), .B (n_85_44), .C1 (n_89_42), .C2 (n_95_39) );
AOI211_X1 g_73_50 (.ZN (n_73_50), .A (n_77_48), .B (n_83_45), .C1 (n_87_43), .C2 (n_93_40) );
AOI211_X1 g_71_51 (.ZN (n_71_51), .A (n_75_49), .B (n_81_46), .C1 (n_85_44), .C2 (n_91_41) );
AOI211_X1 g_69_52 (.ZN (n_69_52), .A (n_73_50), .B (n_79_47), .C1 (n_83_45), .C2 (n_89_42) );
AOI211_X1 g_67_53 (.ZN (n_67_53), .A (n_71_51), .B (n_77_48), .C1 (n_81_46), .C2 (n_87_43) );
AOI211_X1 g_65_54 (.ZN (n_65_54), .A (n_69_52), .B (n_75_49), .C1 (n_79_47), .C2 (n_85_44) );
AOI211_X1 g_63_55 (.ZN (n_63_55), .A (n_67_53), .B (n_73_50), .C1 (n_77_48), .C2 (n_83_45) );
AOI211_X1 g_61_56 (.ZN (n_61_56), .A (n_65_54), .B (n_71_51), .C1 (n_75_49), .C2 (n_81_46) );
AOI211_X1 g_59_57 (.ZN (n_59_57), .A (n_63_55), .B (n_69_52), .C1 (n_73_50), .C2 (n_79_47) );
AOI211_X1 g_57_58 (.ZN (n_57_58), .A (n_61_56), .B (n_67_53), .C1 (n_71_51), .C2 (n_77_48) );
AOI211_X1 g_55_59 (.ZN (n_55_59), .A (n_59_57), .B (n_65_54), .C1 (n_69_52), .C2 (n_75_49) );
AOI211_X1 g_53_60 (.ZN (n_53_60), .A (n_57_58), .B (n_63_55), .C1 (n_67_53), .C2 (n_73_50) );
AOI211_X1 g_51_61 (.ZN (n_51_61), .A (n_55_59), .B (n_61_56), .C1 (n_65_54), .C2 (n_71_51) );
AOI211_X1 g_49_62 (.ZN (n_49_62), .A (n_53_60), .B (n_59_57), .C1 (n_63_55), .C2 (n_69_52) );
AOI211_X1 g_47_63 (.ZN (n_47_63), .A (n_51_61), .B (n_57_58), .C1 (n_61_56), .C2 (n_67_53) );
AOI211_X1 g_45_64 (.ZN (n_45_64), .A (n_49_62), .B (n_55_59), .C1 (n_59_57), .C2 (n_65_54) );
AOI211_X1 g_43_65 (.ZN (n_43_65), .A (n_47_63), .B (n_53_60), .C1 (n_57_58), .C2 (n_63_55) );
AOI211_X1 g_41_66 (.ZN (n_41_66), .A (n_45_64), .B (n_51_61), .C1 (n_55_59), .C2 (n_61_56) );
AOI211_X1 g_39_67 (.ZN (n_39_67), .A (n_43_65), .B (n_49_62), .C1 (n_53_60), .C2 (n_59_57) );
AOI211_X1 g_37_68 (.ZN (n_37_68), .A (n_41_66), .B (n_47_63), .C1 (n_51_61), .C2 (n_57_58) );
AOI211_X1 g_35_69 (.ZN (n_35_69), .A (n_39_67), .B (n_45_64), .C1 (n_49_62), .C2 (n_55_59) );
AOI211_X1 g_33_70 (.ZN (n_33_70), .A (n_37_68), .B (n_43_65), .C1 (n_47_63), .C2 (n_53_60) );
AOI211_X1 g_31_71 (.ZN (n_31_71), .A (n_35_69), .B (n_41_66), .C1 (n_45_64), .C2 (n_51_61) );
AOI211_X1 g_29_72 (.ZN (n_29_72), .A (n_33_70), .B (n_39_67), .C1 (n_43_65), .C2 (n_49_62) );
AOI211_X1 g_27_73 (.ZN (n_27_73), .A (n_31_71), .B (n_37_68), .C1 (n_41_66), .C2 (n_47_63) );
AOI211_X1 g_25_74 (.ZN (n_25_74), .A (n_29_72), .B (n_35_69), .C1 (n_39_67), .C2 (n_45_64) );
AOI211_X1 g_23_75 (.ZN (n_23_75), .A (n_27_73), .B (n_33_70), .C1 (n_37_68), .C2 (n_43_65) );
AOI211_X1 g_24_73 (.ZN (n_24_73), .A (n_25_74), .B (n_31_71), .C1 (n_35_69), .C2 (n_41_66) );
AOI211_X1 g_22_74 (.ZN (n_22_74), .A (n_23_75), .B (n_29_72), .C1 (n_33_70), .C2 (n_39_67) );
AOI211_X1 g_20_75 (.ZN (n_20_75), .A (n_24_73), .B (n_27_73), .C1 (n_31_71), .C2 (n_37_68) );
AOI211_X1 g_18_76 (.ZN (n_18_76), .A (n_22_74), .B (n_25_74), .C1 (n_29_72), .C2 (n_35_69) );
AOI211_X1 g_16_77 (.ZN (n_16_77), .A (n_20_75), .B (n_23_75), .C1 (n_27_73), .C2 (n_33_70) );
AOI211_X1 g_14_78 (.ZN (n_14_78), .A (n_18_76), .B (n_24_73), .C1 (n_25_74), .C2 (n_31_71) );
AOI211_X1 g_12_79 (.ZN (n_12_79), .A (n_16_77), .B (n_22_74), .C1 (n_23_75), .C2 (n_29_72) );
AOI211_X1 g_10_80 (.ZN (n_10_80), .A (n_14_78), .B (n_20_75), .C1 (n_24_73), .C2 (n_27_73) );
AOI211_X1 g_8_81 (.ZN (n_8_81), .A (n_12_79), .B (n_18_76), .C1 (n_22_74), .C2 (n_25_74) );
AOI211_X1 g_6_82 (.ZN (n_6_82), .A (n_10_80), .B (n_16_77), .C1 (n_20_75), .C2 (n_23_75) );
AOI211_X1 g_5_84 (.ZN (n_5_84), .A (n_8_81), .B (n_14_78), .C1 (n_18_76), .C2 (n_24_73) );
AOI211_X1 g_7_83 (.ZN (n_7_83), .A (n_6_82), .B (n_12_79), .C1 (n_16_77), .C2 (n_22_74) );
AOI211_X1 g_9_82 (.ZN (n_9_82), .A (n_5_84), .B (n_10_80), .C1 (n_14_78), .C2 (n_20_75) );
AOI211_X1 g_11_81 (.ZN (n_11_81), .A (n_7_83), .B (n_8_81), .C1 (n_12_79), .C2 (n_18_76) );
AOI211_X1 g_13_80 (.ZN (n_13_80), .A (n_9_82), .B (n_6_82), .C1 (n_10_80), .C2 (n_16_77) );
AOI211_X1 g_15_79 (.ZN (n_15_79), .A (n_11_81), .B (n_5_84), .C1 (n_8_81), .C2 (n_14_78) );
AOI211_X1 g_17_78 (.ZN (n_17_78), .A (n_13_80), .B (n_7_83), .C1 (n_6_82), .C2 (n_12_79) );
AOI211_X1 g_19_77 (.ZN (n_19_77), .A (n_15_79), .B (n_9_82), .C1 (n_5_84), .C2 (n_10_80) );
AOI211_X1 g_21_76 (.ZN (n_21_76), .A (n_17_78), .B (n_11_81), .C1 (n_7_83), .C2 (n_8_81) );
AOI211_X1 g_20_78 (.ZN (n_20_78), .A (n_19_77), .B (n_13_80), .C1 (n_9_82), .C2 (n_6_82) );
AOI211_X1 g_18_77 (.ZN (n_18_77), .A (n_21_76), .B (n_15_79), .C1 (n_11_81), .C2 (n_5_84) );
AOI211_X1 g_20_76 (.ZN (n_20_76), .A (n_20_78), .B (n_17_78), .C1 (n_13_80), .C2 (n_7_83) );
AOI211_X1 g_22_75 (.ZN (n_22_75), .A (n_18_77), .B (n_19_77), .C1 (n_15_79), .C2 (n_9_82) );
AOI211_X1 g_24_74 (.ZN (n_24_74), .A (n_20_76), .B (n_21_76), .C1 (n_17_78), .C2 (n_11_81) );
AOI211_X1 g_26_73 (.ZN (n_26_73), .A (n_22_75), .B (n_20_78), .C1 (n_19_77), .C2 (n_13_80) );
AOI211_X1 g_28_72 (.ZN (n_28_72), .A (n_24_74), .B (n_18_77), .C1 (n_21_76), .C2 (n_15_79) );
AOI211_X1 g_30_71 (.ZN (n_30_71), .A (n_26_73), .B (n_20_76), .C1 (n_20_78), .C2 (n_17_78) );
AOI211_X1 g_32_70 (.ZN (n_32_70), .A (n_28_72), .B (n_22_75), .C1 (n_18_77), .C2 (n_19_77) );
AOI211_X1 g_34_69 (.ZN (n_34_69), .A (n_30_71), .B (n_24_74), .C1 (n_20_76), .C2 (n_21_76) );
AOI211_X1 g_36_68 (.ZN (n_36_68), .A (n_32_70), .B (n_26_73), .C1 (n_22_75), .C2 (n_20_78) );
AOI211_X1 g_38_67 (.ZN (n_38_67), .A (n_34_69), .B (n_28_72), .C1 (n_24_74), .C2 (n_18_77) );
AOI211_X1 g_40_66 (.ZN (n_40_66), .A (n_36_68), .B (n_30_71), .C1 (n_26_73), .C2 (n_20_76) );
AOI211_X1 g_42_65 (.ZN (n_42_65), .A (n_38_67), .B (n_32_70), .C1 (n_28_72), .C2 (n_22_75) );
AOI211_X1 g_44_64 (.ZN (n_44_64), .A (n_40_66), .B (n_34_69), .C1 (n_30_71), .C2 (n_24_74) );
AOI211_X1 g_46_63 (.ZN (n_46_63), .A (n_42_65), .B (n_36_68), .C1 (n_32_70), .C2 (n_26_73) );
AOI211_X1 g_48_62 (.ZN (n_48_62), .A (n_44_64), .B (n_38_67), .C1 (n_34_69), .C2 (n_28_72) );
AOI211_X1 g_50_61 (.ZN (n_50_61), .A (n_46_63), .B (n_40_66), .C1 (n_36_68), .C2 (n_30_71) );
AOI211_X1 g_52_60 (.ZN (n_52_60), .A (n_48_62), .B (n_42_65), .C1 (n_38_67), .C2 (n_32_70) );
AOI211_X1 g_54_59 (.ZN (n_54_59), .A (n_50_61), .B (n_44_64), .C1 (n_40_66), .C2 (n_34_69) );
AOI211_X1 g_56_58 (.ZN (n_56_58), .A (n_52_60), .B (n_46_63), .C1 (n_42_65), .C2 (n_36_68) );
AOI211_X1 g_58_57 (.ZN (n_58_57), .A (n_54_59), .B (n_48_62), .C1 (n_44_64), .C2 (n_38_67) );
AOI211_X1 g_60_56 (.ZN (n_60_56), .A (n_56_58), .B (n_50_61), .C1 (n_46_63), .C2 (n_40_66) );
AOI211_X1 g_62_55 (.ZN (n_62_55), .A (n_58_57), .B (n_52_60), .C1 (n_48_62), .C2 (n_42_65) );
AOI211_X1 g_64_54 (.ZN (n_64_54), .A (n_60_56), .B (n_54_59), .C1 (n_50_61), .C2 (n_44_64) );
AOI211_X1 g_66_53 (.ZN (n_66_53), .A (n_62_55), .B (n_56_58), .C1 (n_52_60), .C2 (n_46_63) );
AOI211_X1 g_68_52 (.ZN (n_68_52), .A (n_64_54), .B (n_58_57), .C1 (n_54_59), .C2 (n_48_62) );
AOI211_X1 g_70_51 (.ZN (n_70_51), .A (n_66_53), .B (n_60_56), .C1 (n_56_58), .C2 (n_50_61) );
AOI211_X1 g_72_50 (.ZN (n_72_50), .A (n_68_52), .B (n_62_55), .C1 (n_58_57), .C2 (n_52_60) );
AOI211_X1 g_74_49 (.ZN (n_74_49), .A (n_70_51), .B (n_64_54), .C1 (n_60_56), .C2 (n_54_59) );
AOI211_X1 g_76_48 (.ZN (n_76_48), .A (n_72_50), .B (n_66_53), .C1 (n_62_55), .C2 (n_56_58) );
AOI211_X1 g_78_47 (.ZN (n_78_47), .A (n_74_49), .B (n_68_52), .C1 (n_64_54), .C2 (n_58_57) );
AOI211_X1 g_80_46 (.ZN (n_80_46), .A (n_76_48), .B (n_70_51), .C1 (n_66_53), .C2 (n_60_56) );
AOI211_X1 g_82_45 (.ZN (n_82_45), .A (n_78_47), .B (n_72_50), .C1 (n_68_52), .C2 (n_62_55) );
AOI211_X1 g_84_44 (.ZN (n_84_44), .A (n_80_46), .B (n_74_49), .C1 (n_70_51), .C2 (n_64_54) );
AOI211_X1 g_86_43 (.ZN (n_86_43), .A (n_82_45), .B (n_76_48), .C1 (n_72_50), .C2 (n_66_53) );
AOI211_X1 g_88_42 (.ZN (n_88_42), .A (n_84_44), .B (n_78_47), .C1 (n_74_49), .C2 (n_68_52) );
AOI211_X1 g_90_41 (.ZN (n_90_41), .A (n_86_43), .B (n_80_46), .C1 (n_76_48), .C2 (n_70_51) );
AOI211_X1 g_92_40 (.ZN (n_92_40), .A (n_88_42), .B (n_82_45), .C1 (n_78_47), .C2 (n_72_50) );
AOI211_X1 g_94_39 (.ZN (n_94_39), .A (n_90_41), .B (n_84_44), .C1 (n_80_46), .C2 (n_74_49) );
AOI211_X1 g_96_38 (.ZN (n_96_38), .A (n_92_40), .B (n_86_43), .C1 (n_82_45), .C2 (n_76_48) );
AOI211_X1 g_98_37 (.ZN (n_98_37), .A (n_94_39), .B (n_88_42), .C1 (n_84_44), .C2 (n_78_47) );
AOI211_X1 g_100_36 (.ZN (n_100_36), .A (n_96_38), .B (n_90_41), .C1 (n_86_43), .C2 (n_80_46) );
AOI211_X1 g_102_35 (.ZN (n_102_35), .A (n_98_37), .B (n_92_40), .C1 (n_88_42), .C2 (n_82_45) );
AOI211_X1 g_104_34 (.ZN (n_104_34), .A (n_100_36), .B (n_94_39), .C1 (n_90_41), .C2 (n_84_44) );
AOI211_X1 g_106_33 (.ZN (n_106_33), .A (n_102_35), .B (n_96_38), .C1 (n_92_40), .C2 (n_86_43) );
AOI211_X1 g_108_32 (.ZN (n_108_32), .A (n_104_34), .B (n_98_37), .C1 (n_94_39), .C2 (n_88_42) );
AOI211_X1 g_110_31 (.ZN (n_110_31), .A (n_106_33), .B (n_100_36), .C1 (n_96_38), .C2 (n_90_41) );
AOI211_X1 g_112_30 (.ZN (n_112_30), .A (n_108_32), .B (n_102_35), .C1 (n_98_37), .C2 (n_92_40) );
AOI211_X1 g_114_29 (.ZN (n_114_29), .A (n_110_31), .B (n_104_34), .C1 (n_100_36), .C2 (n_94_39) );
AOI211_X1 g_116_28 (.ZN (n_116_28), .A (n_112_30), .B (n_106_33), .C1 (n_102_35), .C2 (n_96_38) );
AOI211_X1 g_115_30 (.ZN (n_115_30), .A (n_114_29), .B (n_108_32), .C1 (n_104_34), .C2 (n_98_37) );
AOI211_X1 g_117_29 (.ZN (n_117_29), .A (n_116_28), .B (n_110_31), .C1 (n_106_33), .C2 (n_100_36) );
AOI211_X1 g_119_28 (.ZN (n_119_28), .A (n_115_30), .B (n_112_30), .C1 (n_108_32), .C2 (n_102_35) );
AOI211_X1 g_121_27 (.ZN (n_121_27), .A (n_117_29), .B (n_114_29), .C1 (n_110_31), .C2 (n_104_34) );
AOI211_X1 g_123_26 (.ZN (n_123_26), .A (n_119_28), .B (n_116_28), .C1 (n_112_30), .C2 (n_106_33) );
AOI211_X1 g_121_25 (.ZN (n_121_25), .A (n_121_27), .B (n_115_30), .C1 (n_114_29), .C2 (n_108_32) );
AOI211_X1 g_123_24 (.ZN (n_123_24), .A (n_123_26), .B (n_117_29), .C1 (n_116_28), .C2 (n_110_31) );
AOI211_X1 g_125_23 (.ZN (n_125_23), .A (n_121_25), .B (n_119_28), .C1 (n_115_30), .C2 (n_112_30) );
AOI211_X1 g_127_22 (.ZN (n_127_22), .A (n_123_24), .B (n_121_27), .C1 (n_117_29), .C2 (n_114_29) );
AOI211_X1 g_126_24 (.ZN (n_126_24), .A (n_125_23), .B (n_123_26), .C1 (n_119_28), .C2 (n_116_28) );
AOI211_X1 g_128_23 (.ZN (n_128_23), .A (n_127_22), .B (n_121_25), .C1 (n_121_27), .C2 (n_115_30) );
AOI211_X1 g_130_22 (.ZN (n_130_22), .A (n_126_24), .B (n_123_24), .C1 (n_123_26), .C2 (n_117_29) );
AOI211_X1 g_132_21 (.ZN (n_132_21), .A (n_128_23), .B (n_125_23), .C1 (n_121_25), .C2 (n_119_28) );
AOI211_X1 g_131_23 (.ZN (n_131_23), .A (n_130_22), .B (n_127_22), .C1 (n_123_24), .C2 (n_121_27) );
AOI211_X1 g_129_24 (.ZN (n_129_24), .A (n_132_21), .B (n_126_24), .C1 (n_125_23), .C2 (n_123_26) );
AOI211_X1 g_127_25 (.ZN (n_127_25), .A (n_131_23), .B (n_128_23), .C1 (n_127_22), .C2 (n_121_25) );
AOI211_X1 g_125_26 (.ZN (n_125_26), .A (n_129_24), .B (n_130_22), .C1 (n_126_24), .C2 (n_123_24) );
AOI211_X1 g_123_27 (.ZN (n_123_27), .A (n_127_25), .B (n_132_21), .C1 (n_128_23), .C2 (n_125_23) );
AOI211_X1 g_124_25 (.ZN (n_124_25), .A (n_125_26), .B (n_131_23), .C1 (n_130_22), .C2 (n_127_22) );
AOI211_X1 g_122_26 (.ZN (n_122_26), .A (n_123_27), .B (n_129_24), .C1 (n_132_21), .C2 (n_126_24) );
AOI211_X1 g_120_27 (.ZN (n_120_27), .A (n_124_25), .B (n_127_25), .C1 (n_131_23), .C2 (n_128_23) );
AOI211_X1 g_118_28 (.ZN (n_118_28), .A (n_122_26), .B (n_125_26), .C1 (n_129_24), .C2 (n_130_22) );
AOI211_X1 g_116_29 (.ZN (n_116_29), .A (n_120_27), .B (n_123_27), .C1 (n_127_25), .C2 (n_132_21) );
AOI211_X1 g_114_30 (.ZN (n_114_30), .A (n_118_28), .B (n_124_25), .C1 (n_125_26), .C2 (n_131_23) );
AOI211_X1 g_112_31 (.ZN (n_112_31), .A (n_116_29), .B (n_122_26), .C1 (n_123_27), .C2 (n_129_24) );
AOI211_X1 g_111_33 (.ZN (n_111_33), .A (n_114_30), .B (n_120_27), .C1 (n_124_25), .C2 (n_127_25) );
AOI211_X1 g_113_32 (.ZN (n_113_32), .A (n_112_31), .B (n_118_28), .C1 (n_122_26), .C2 (n_125_26) );
AOI211_X1 g_115_31 (.ZN (n_115_31), .A (n_111_33), .B (n_116_29), .C1 (n_120_27), .C2 (n_123_27) );
AOI211_X1 g_117_30 (.ZN (n_117_30), .A (n_113_32), .B (n_114_30), .C1 (n_118_28), .C2 (n_124_25) );
AOI211_X1 g_119_29 (.ZN (n_119_29), .A (n_115_31), .B (n_112_31), .C1 (n_116_29), .C2 (n_122_26) );
AOI211_X1 g_121_28 (.ZN (n_121_28), .A (n_117_30), .B (n_111_33), .C1 (n_114_30), .C2 (n_120_27) );
AOI211_X1 g_120_30 (.ZN (n_120_30), .A (n_119_29), .B (n_113_32), .C1 (n_112_31), .C2 (n_118_28) );
AOI211_X1 g_118_29 (.ZN (n_118_29), .A (n_121_28), .B (n_115_31), .C1 (n_111_33), .C2 (n_116_29) );
AOI211_X1 g_120_28 (.ZN (n_120_28), .A (n_120_30), .B (n_117_30), .C1 (n_113_32), .C2 (n_114_30) );
AOI211_X1 g_122_27 (.ZN (n_122_27), .A (n_118_29), .B (n_119_29), .C1 (n_115_31), .C2 (n_112_31) );
AOI211_X1 g_124_26 (.ZN (n_124_26), .A (n_120_28), .B (n_121_28), .C1 (n_117_30), .C2 (n_111_33) );
AOI211_X1 g_126_25 (.ZN (n_126_25), .A (n_122_27), .B (n_120_30), .C1 (n_119_29), .C2 (n_113_32) );
AOI211_X1 g_128_24 (.ZN (n_128_24), .A (n_124_26), .B (n_118_29), .C1 (n_121_28), .C2 (n_115_31) );
AOI211_X1 g_130_23 (.ZN (n_130_23), .A (n_126_25), .B (n_120_28), .C1 (n_120_30), .C2 (n_117_30) );
AOI211_X1 g_131_21 (.ZN (n_131_21), .A (n_128_24), .B (n_122_27), .C1 (n_118_29), .C2 (n_119_29) );
AOI211_X1 g_133_20 (.ZN (n_133_20), .A (n_130_23), .B (n_124_26), .C1 (n_120_28), .C2 (n_121_28) );
AOI211_X1 g_135_19 (.ZN (n_135_19), .A (n_131_21), .B (n_126_25), .C1 (n_122_27), .C2 (n_120_30) );
AOI211_X1 g_137_18 (.ZN (n_137_18), .A (n_133_20), .B (n_128_24), .C1 (n_124_26), .C2 (n_118_29) );
AOI211_X1 g_139_19 (.ZN (n_139_19), .A (n_135_19), .B (n_130_23), .C1 (n_126_25), .C2 (n_120_28) );
AOI211_X1 g_137_20 (.ZN (n_137_20), .A (n_137_18), .B (n_131_21), .C1 (n_128_24), .C2 (n_122_27) );
AOI211_X1 g_136_18 (.ZN (n_136_18), .A (n_139_19), .B (n_133_20), .C1 (n_130_23), .C2 (n_124_26) );
AOI211_X1 g_134_19 (.ZN (n_134_19), .A (n_137_20), .B (n_135_19), .C1 (n_131_21), .C2 (n_126_25) );
AOI211_X1 g_132_20 (.ZN (n_132_20), .A (n_136_18), .B (n_137_18), .C1 (n_133_20), .C2 (n_128_24) );
AOI211_X1 g_133_22 (.ZN (n_133_22), .A (n_134_19), .B (n_139_19), .C1 (n_135_19), .C2 (n_130_23) );
AOI211_X1 g_135_21 (.ZN (n_135_21), .A (n_132_20), .B (n_137_20), .C1 (n_137_18), .C2 (n_131_21) );
AOI211_X1 g_134_23 (.ZN (n_134_23), .A (n_133_22), .B (n_136_18), .C1 (n_139_19), .C2 (n_133_20) );
AOI211_X1 g_132_22 (.ZN (n_132_22), .A (n_135_21), .B (n_134_19), .C1 (n_137_20), .C2 (n_135_19) );
AOI211_X1 g_134_21 (.ZN (n_134_21), .A (n_134_23), .B (n_132_20), .C1 (n_136_18), .C2 (n_137_18) );
AOI211_X1 g_136_20 (.ZN (n_136_20), .A (n_132_22), .B (n_133_22), .C1 (n_134_19), .C2 (n_139_19) );
AOI211_X1 g_138_19 (.ZN (n_138_19), .A (n_134_21), .B (n_135_21), .C1 (n_132_20), .C2 (n_137_20) );
AOI211_X1 g_139_21 (.ZN (n_139_21), .A (n_136_20), .B (n_134_23), .C1 (n_133_22), .C2 (n_136_18) );
AOI211_X1 g_137_22 (.ZN (n_137_22), .A (n_138_19), .B (n_132_22), .C1 (n_135_21), .C2 (n_134_19) );
AOI211_X1 g_138_20 (.ZN (n_138_20), .A (n_139_21), .B (n_134_21), .C1 (n_134_23), .C2 (n_132_20) );
AOI211_X1 g_136_21 (.ZN (n_136_21), .A (n_137_22), .B (n_136_20), .C1 (n_132_22), .C2 (n_133_22) );
AOI211_X1 g_137_19 (.ZN (n_137_19), .A (n_138_20), .B (n_138_19), .C1 (n_134_21), .C2 (n_135_21) );
AOI211_X1 g_135_20 (.ZN (n_135_20), .A (n_136_21), .B (n_139_21), .C1 (n_136_20), .C2 (n_134_23) );
AOI211_X1 g_133_21 (.ZN (n_133_21), .A (n_137_19), .B (n_137_22), .C1 (n_138_19), .C2 (n_132_22) );
AOI211_X1 g_131_22 (.ZN (n_131_22), .A (n_135_20), .B (n_138_20), .C1 (n_139_21), .C2 (n_134_21) );
AOI211_X1 g_129_23 (.ZN (n_129_23), .A (n_133_21), .B (n_136_21), .C1 (n_137_22), .C2 (n_136_20) );
AOI211_X1 g_127_24 (.ZN (n_127_24), .A (n_131_22), .B (n_137_19), .C1 (n_138_20), .C2 (n_138_19) );
AOI211_X1 g_125_25 (.ZN (n_125_25), .A (n_129_23), .B (n_135_20), .C1 (n_136_21), .C2 (n_139_21) );
AOI211_X1 g_124_27 (.ZN (n_124_27), .A (n_127_24), .B (n_133_21), .C1 (n_137_19), .C2 (n_137_22) );
AOI211_X1 g_126_26 (.ZN (n_126_26), .A (n_125_25), .B (n_131_22), .C1 (n_135_20), .C2 (n_138_20) );
AOI211_X1 g_128_25 (.ZN (n_128_25), .A (n_124_27), .B (n_129_23), .C1 (n_133_21), .C2 (n_136_21) );
AOI211_X1 g_130_24 (.ZN (n_130_24), .A (n_126_26), .B (n_127_24), .C1 (n_131_22), .C2 (n_137_19) );
AOI211_X1 g_132_23 (.ZN (n_132_23), .A (n_128_25), .B (n_125_25), .C1 (n_129_23), .C2 (n_135_20) );
AOI211_X1 g_134_22 (.ZN (n_134_22), .A (n_130_24), .B (n_124_27), .C1 (n_127_24), .C2 (n_133_21) );
AOI211_X1 g_133_24 (.ZN (n_133_24), .A (n_132_23), .B (n_126_26), .C1 (n_125_25), .C2 (n_131_22) );
AOI211_X1 g_135_23 (.ZN (n_135_23), .A (n_134_22), .B (n_128_25), .C1 (n_124_27), .C2 (n_129_23) );
AOI211_X1 g_134_25 (.ZN (n_134_25), .A (n_133_24), .B (n_130_24), .C1 (n_126_26), .C2 (n_127_24) );
AOI211_X1 g_132_24 (.ZN (n_132_24), .A (n_135_23), .B (n_132_23), .C1 (n_128_25), .C2 (n_125_25) );
AOI211_X1 g_130_25 (.ZN (n_130_25), .A (n_134_25), .B (n_134_22), .C1 (n_130_24), .C2 (n_124_27) );
AOI211_X1 g_128_26 (.ZN (n_128_26), .A (n_132_24), .B (n_133_24), .C1 (n_132_23), .C2 (n_126_26) );
AOI211_X1 g_126_27 (.ZN (n_126_27), .A (n_130_25), .B (n_135_23), .C1 (n_134_22), .C2 (n_128_25) );
AOI211_X1 g_124_28 (.ZN (n_124_28), .A (n_128_26), .B (n_134_25), .C1 (n_133_24), .C2 (n_130_24) );
AOI211_X1 g_122_29 (.ZN (n_122_29), .A (n_126_27), .B (n_132_24), .C1 (n_135_23), .C2 (n_132_23) );
AOI211_X1 g_121_31 (.ZN (n_121_31), .A (n_124_28), .B (n_130_25), .C1 (n_134_25), .C2 (n_134_22) );
AOI211_X1 g_120_29 (.ZN (n_120_29), .A (n_122_29), .B (n_128_26), .C1 (n_132_24), .C2 (n_133_24) );
AOI211_X1 g_122_28 (.ZN (n_122_28), .A (n_121_31), .B (n_126_27), .C1 (n_130_25), .C2 (n_135_23) );
AOI211_X1 g_121_30 (.ZN (n_121_30), .A (n_120_29), .B (n_124_28), .C1 (n_128_26), .C2 (n_134_25) );
AOI211_X1 g_123_29 (.ZN (n_123_29), .A (n_122_28), .B (n_122_29), .C1 (n_126_27), .C2 (n_132_24) );
AOI211_X1 g_125_28 (.ZN (n_125_28), .A (n_121_30), .B (n_121_31), .C1 (n_124_28), .C2 (n_130_25) );
AOI211_X1 g_127_27 (.ZN (n_127_27), .A (n_123_29), .B (n_120_29), .C1 (n_122_29), .C2 (n_128_26) );
AOI211_X1 g_129_26 (.ZN (n_129_26), .A (n_125_28), .B (n_122_28), .C1 (n_121_31), .C2 (n_126_27) );
AOI211_X1 g_131_25 (.ZN (n_131_25), .A (n_127_27), .B (n_121_30), .C1 (n_120_29), .C2 (n_124_28) );
AOI211_X1 g_130_27 (.ZN (n_130_27), .A (n_129_26), .B (n_123_29), .C1 (n_122_28), .C2 (n_122_29) );
AOI211_X1 g_132_26 (.ZN (n_132_26), .A (n_131_25), .B (n_125_28), .C1 (n_121_30), .C2 (n_121_31) );
AOI211_X1 g_131_24 (.ZN (n_131_24), .A (n_130_27), .B (n_127_27), .C1 (n_123_29), .C2 (n_120_29) );
AOI211_X1 g_133_23 (.ZN (n_133_23), .A (n_132_26), .B (n_129_26), .C1 (n_125_28), .C2 (n_122_28) );
AOI211_X1 g_135_22 (.ZN (n_135_22), .A (n_131_24), .B (n_131_25), .C1 (n_127_27), .C2 (n_121_30) );
AOI211_X1 g_137_21 (.ZN (n_137_21), .A (n_133_23), .B (n_130_27), .C1 (n_129_26), .C2 (n_123_29) );
AOI211_X1 g_139_20 (.ZN (n_139_20), .A (n_135_22), .B (n_132_26), .C1 (n_131_25), .C2 (n_125_28) );
AOI211_X1 g_138_22 (.ZN (n_138_22), .A (n_137_21), .B (n_131_24), .C1 (n_130_27), .C2 (n_127_27) );
AOI211_X1 g_140_21 (.ZN (n_140_21), .A (n_139_20), .B (n_133_23), .C1 (n_132_26), .C2 (n_129_26) );
AOI211_X1 g_142_20 (.ZN (n_142_20), .A (n_138_22), .B (n_135_22), .C1 (n_131_24), .C2 (n_131_25) );
AOI211_X1 g_144_19 (.ZN (n_144_19), .A (n_140_21), .B (n_137_21), .C1 (n_133_23), .C2 (n_130_27) );
AOI211_X1 g_146_18 (.ZN (n_146_18), .A (n_142_20), .B (n_139_20), .C1 (n_135_22), .C2 (n_132_26) );
AOI211_X1 g_147_20 (.ZN (n_147_20), .A (n_144_19), .B (n_138_22), .C1 (n_137_21), .C2 (n_131_24) );
AOI211_X1 g_149_21 (.ZN (n_149_21), .A (n_146_18), .B (n_140_21), .C1 (n_139_20), .C2 (n_133_23) );
AOI211_X1 g_148_19 (.ZN (n_148_19), .A (n_147_20), .B (n_142_20), .C1 (n_138_22), .C2 (n_135_22) );
AOI211_X1 g_146_20 (.ZN (n_146_20), .A (n_149_21), .B (n_144_19), .C1 (n_140_21), .C2 (n_137_21) );
AOI211_X1 g_147_22 (.ZN (n_147_22), .A (n_148_19), .B (n_146_18), .C1 (n_142_20), .C2 (n_139_20) );
AOI211_X1 g_145_21 (.ZN (n_145_21), .A (n_146_20), .B (n_147_20), .C1 (n_144_19), .C2 (n_138_22) );
AOI211_X1 g_146_19 (.ZN (n_146_19), .A (n_147_22), .B (n_149_21), .C1 (n_146_18), .C2 (n_140_21) );
AOI211_X1 g_144_18 (.ZN (n_144_18), .A (n_145_21), .B (n_148_19), .C1 (n_147_20), .C2 (n_142_20) );
AOI211_X1 g_143_20 (.ZN (n_143_20), .A (n_146_19), .B (n_146_20), .C1 (n_149_21), .C2 (n_144_19) );
AOI211_X1 g_141_21 (.ZN (n_141_21), .A (n_144_18), .B (n_147_22), .C1 (n_148_19), .C2 (n_146_18) );
AOI211_X1 g_142_19 (.ZN (n_142_19), .A (n_143_20), .B (n_145_21), .C1 (n_146_20), .C2 (n_147_20) );
AOI211_X1 g_144_20 (.ZN (n_144_20), .A (n_141_21), .B (n_146_19), .C1 (n_147_22), .C2 (n_149_21) );
AOI211_X1 g_143_22 (.ZN (n_143_22), .A (n_142_19), .B (n_144_18), .C1 (n_145_21), .C2 (n_148_19) );
AOI211_X1 g_145_23 (.ZN (n_145_23), .A (n_144_20), .B (n_143_20), .C1 (n_146_19), .C2 (n_146_20) );
AOI211_X1 g_144_21 (.ZN (n_144_21), .A (n_143_22), .B (n_141_21), .C1 (n_144_18), .C2 (n_147_22) );
AOI211_X1 g_142_22 (.ZN (n_142_22), .A (n_145_23), .B (n_142_19), .C1 (n_143_20), .C2 (n_145_21) );
AOI211_X1 g_140_23 (.ZN (n_140_23), .A (n_144_21), .B (n_144_20), .C1 (n_141_21), .C2 (n_146_19) );
AOI211_X1 g_138_24 (.ZN (n_138_24), .A (n_142_22), .B (n_143_22), .C1 (n_142_19), .C2 (n_144_18) );
AOI211_X1 g_136_23 (.ZN (n_136_23), .A (n_140_23), .B (n_145_23), .C1 (n_144_20), .C2 (n_143_20) );
AOI211_X1 g_134_24 (.ZN (n_134_24), .A (n_138_24), .B (n_144_21), .C1 (n_143_22), .C2 (n_141_21) );
AOI211_X1 g_132_25 (.ZN (n_132_25), .A (n_136_23), .B (n_142_22), .C1 (n_145_23), .C2 (n_142_19) );
AOI211_X1 g_130_26 (.ZN (n_130_26), .A (n_134_24), .B (n_140_23), .C1 (n_144_21), .C2 (n_144_20) );
AOI211_X1 g_128_27 (.ZN (n_128_27), .A (n_132_25), .B (n_138_24), .C1 (n_142_22), .C2 (n_143_22) );
AOI211_X1 g_129_25 (.ZN (n_129_25), .A (n_130_26), .B (n_136_23), .C1 (n_140_23), .C2 (n_145_23) );
AOI211_X1 g_127_26 (.ZN (n_127_26), .A (n_128_27), .B (n_134_24), .C1 (n_138_24), .C2 (n_144_21) );
AOI211_X1 g_125_27 (.ZN (n_125_27), .A (n_129_25), .B (n_132_25), .C1 (n_136_23), .C2 (n_142_22) );
AOI211_X1 g_123_28 (.ZN (n_123_28), .A (n_127_26), .B (n_130_26), .C1 (n_134_24), .C2 (n_140_23) );
AOI211_X1 g_121_29 (.ZN (n_121_29), .A (n_125_27), .B (n_128_27), .C1 (n_132_25), .C2 (n_138_24) );
AOI211_X1 g_119_30 (.ZN (n_119_30), .A (n_123_28), .B (n_129_25), .C1 (n_130_26), .C2 (n_136_23) );
AOI211_X1 g_117_31 (.ZN (n_117_31), .A (n_121_29), .B (n_127_26), .C1 (n_128_27), .C2 (n_134_24) );
AOI211_X1 g_119_32 (.ZN (n_119_32), .A (n_119_30), .B (n_125_27), .C1 (n_129_25), .C2 (n_132_25) );
AOI211_X1 g_118_30 (.ZN (n_118_30), .A (n_117_31), .B (n_123_28), .C1 (n_127_26), .C2 (n_130_26) );
AOI211_X1 g_116_31 (.ZN (n_116_31), .A (n_119_32), .B (n_121_29), .C1 (n_125_27), .C2 (n_128_27) );
AOI211_X1 g_114_32 (.ZN (n_114_32), .A (n_118_30), .B (n_119_30), .C1 (n_123_28), .C2 (n_129_25) );
AOI211_X1 g_112_33 (.ZN (n_112_33), .A (n_116_31), .B (n_117_31), .C1 (n_121_29), .C2 (n_127_26) );
AOI211_X1 g_113_31 (.ZN (n_113_31), .A (n_114_32), .B (n_119_32), .C1 (n_119_30), .C2 (n_125_27) );
AOI211_X1 g_111_32 (.ZN (n_111_32), .A (n_112_33), .B (n_118_30), .C1 (n_117_31), .C2 (n_123_28) );
AOI211_X1 g_109_33 (.ZN (n_109_33), .A (n_113_31), .B (n_116_31), .C1 (n_119_32), .C2 (n_121_29) );
AOI211_X1 g_107_34 (.ZN (n_107_34), .A (n_111_32), .B (n_114_32), .C1 (n_118_30), .C2 (n_119_30) );
AOI211_X1 g_105_33 (.ZN (n_105_33), .A (n_109_33), .B (n_112_33), .C1 (n_116_31), .C2 (n_117_31) );
AOI211_X1 g_103_34 (.ZN (n_103_34), .A (n_107_34), .B (n_113_31), .C1 (n_114_32), .C2 (n_119_32) );
AOI211_X1 g_101_35 (.ZN (n_101_35), .A (n_105_33), .B (n_111_32), .C1 (n_112_33), .C2 (n_118_30) );
AOI211_X1 g_99_36 (.ZN (n_99_36), .A (n_103_34), .B (n_109_33), .C1 (n_113_31), .C2 (n_116_31) );
AOI211_X1 g_97_37 (.ZN (n_97_37), .A (n_101_35), .B (n_107_34), .C1 (n_111_32), .C2 (n_114_32) );
AOI211_X1 g_95_38 (.ZN (n_95_38), .A (n_99_36), .B (n_105_33), .C1 (n_109_33), .C2 (n_112_33) );
AOI211_X1 g_93_39 (.ZN (n_93_39), .A (n_97_37), .B (n_103_34), .C1 (n_107_34), .C2 (n_113_31) );
AOI211_X1 g_91_40 (.ZN (n_91_40), .A (n_95_38), .B (n_101_35), .C1 (n_105_33), .C2 (n_111_32) );
AOI211_X1 g_89_41 (.ZN (n_89_41), .A (n_93_39), .B (n_99_36), .C1 (n_103_34), .C2 (n_109_33) );
AOI211_X1 g_87_42 (.ZN (n_87_42), .A (n_91_40), .B (n_97_37), .C1 (n_101_35), .C2 (n_107_34) );
AOI211_X1 g_85_43 (.ZN (n_85_43), .A (n_89_41), .B (n_95_38), .C1 (n_99_36), .C2 (n_105_33) );
AOI211_X1 g_83_44 (.ZN (n_83_44), .A (n_87_42), .B (n_93_39), .C1 (n_97_37), .C2 (n_103_34) );
AOI211_X1 g_81_45 (.ZN (n_81_45), .A (n_85_43), .B (n_91_40), .C1 (n_95_38), .C2 (n_101_35) );
AOI211_X1 g_79_46 (.ZN (n_79_46), .A (n_83_44), .B (n_89_41), .C1 (n_93_39), .C2 (n_99_36) );
AOI211_X1 g_77_47 (.ZN (n_77_47), .A (n_81_45), .B (n_87_42), .C1 (n_91_40), .C2 (n_97_37) );
AOI211_X1 g_75_48 (.ZN (n_75_48), .A (n_79_46), .B (n_85_43), .C1 (n_89_41), .C2 (n_95_38) );
AOI211_X1 g_73_49 (.ZN (n_73_49), .A (n_77_47), .B (n_83_44), .C1 (n_87_42), .C2 (n_93_39) );
AOI211_X1 g_72_51 (.ZN (n_72_51), .A (n_75_48), .B (n_81_45), .C1 (n_85_43), .C2 (n_91_40) );
AOI211_X1 g_74_50 (.ZN (n_74_50), .A (n_73_49), .B (n_79_46), .C1 (n_83_44), .C2 (n_89_41) );
AOI211_X1 g_76_49 (.ZN (n_76_49), .A (n_72_51), .B (n_77_47), .C1 (n_81_45), .C2 (n_87_42) );
AOI211_X1 g_78_48 (.ZN (n_78_48), .A (n_74_50), .B (n_75_48), .C1 (n_79_46), .C2 (n_85_43) );
AOI211_X1 g_80_47 (.ZN (n_80_47), .A (n_76_49), .B (n_73_49), .C1 (n_77_47), .C2 (n_83_44) );
AOI211_X1 g_82_46 (.ZN (n_82_46), .A (n_78_48), .B (n_72_51), .C1 (n_75_48), .C2 (n_81_45) );
AOI211_X1 g_84_45 (.ZN (n_84_45), .A (n_80_47), .B (n_74_50), .C1 (n_73_49), .C2 (n_79_46) );
AOI211_X1 g_86_44 (.ZN (n_86_44), .A (n_82_46), .B (n_76_49), .C1 (n_72_51), .C2 (n_77_47) );
AOI211_X1 g_88_43 (.ZN (n_88_43), .A (n_84_45), .B (n_78_48), .C1 (n_74_50), .C2 (n_75_48) );
AOI211_X1 g_90_42 (.ZN (n_90_42), .A (n_86_44), .B (n_80_47), .C1 (n_76_49), .C2 (n_73_49) );
AOI211_X1 g_92_41 (.ZN (n_92_41), .A (n_88_43), .B (n_82_46), .C1 (n_78_48), .C2 (n_72_51) );
AOI211_X1 g_94_40 (.ZN (n_94_40), .A (n_90_42), .B (n_84_45), .C1 (n_80_47), .C2 (n_74_50) );
AOI211_X1 g_96_39 (.ZN (n_96_39), .A (n_92_41), .B (n_86_44), .C1 (n_82_46), .C2 (n_76_49) );
AOI211_X1 g_98_38 (.ZN (n_98_38), .A (n_94_40), .B (n_88_43), .C1 (n_84_45), .C2 (n_78_48) );
AOI211_X1 g_100_37 (.ZN (n_100_37), .A (n_96_39), .B (n_90_42), .C1 (n_86_44), .C2 (n_80_47) );
AOI211_X1 g_102_36 (.ZN (n_102_36), .A (n_98_38), .B (n_92_41), .C1 (n_88_43), .C2 (n_82_46) );
AOI211_X1 g_104_35 (.ZN (n_104_35), .A (n_100_37), .B (n_94_40), .C1 (n_90_42), .C2 (n_84_45) );
AOI211_X1 g_106_34 (.ZN (n_106_34), .A (n_102_36), .B (n_96_39), .C1 (n_92_41), .C2 (n_86_44) );
AOI211_X1 g_108_33 (.ZN (n_108_33), .A (n_104_35), .B (n_98_38), .C1 (n_94_40), .C2 (n_88_43) );
AOI211_X1 g_110_34 (.ZN (n_110_34), .A (n_106_34), .B (n_100_37), .C1 (n_96_39), .C2 (n_90_42) );
AOI211_X1 g_108_35 (.ZN (n_108_35), .A (n_108_33), .B (n_102_36), .C1 (n_98_38), .C2 (n_92_41) );
AOI211_X1 g_106_36 (.ZN (n_106_36), .A (n_110_34), .B (n_104_35), .C1 (n_100_37), .C2 (n_94_40) );
AOI211_X1 g_104_37 (.ZN (n_104_37), .A (n_108_35), .B (n_106_34), .C1 (n_102_36), .C2 (n_96_39) );
AOI211_X1 g_105_35 (.ZN (n_105_35), .A (n_106_36), .B (n_108_33), .C1 (n_104_35), .C2 (n_98_38) );
AOI211_X1 g_103_36 (.ZN (n_103_36), .A (n_104_37), .B (n_110_34), .C1 (n_106_34), .C2 (n_100_37) );
AOI211_X1 g_101_37 (.ZN (n_101_37), .A (n_105_35), .B (n_108_35), .C1 (n_108_33), .C2 (n_102_36) );
AOI211_X1 g_99_38 (.ZN (n_99_38), .A (n_103_36), .B (n_106_36), .C1 (n_110_34), .C2 (n_104_35) );
AOI211_X1 g_97_39 (.ZN (n_97_39), .A (n_101_37), .B (n_104_37), .C1 (n_108_35), .C2 (n_106_34) );
AOI211_X1 g_95_40 (.ZN (n_95_40), .A (n_99_38), .B (n_105_35), .C1 (n_106_36), .C2 (n_108_33) );
AOI211_X1 g_93_41 (.ZN (n_93_41), .A (n_97_39), .B (n_103_36), .C1 (n_104_37), .C2 (n_110_34) );
AOI211_X1 g_91_42 (.ZN (n_91_42), .A (n_95_40), .B (n_101_37), .C1 (n_105_35), .C2 (n_108_35) );
AOI211_X1 g_89_43 (.ZN (n_89_43), .A (n_93_41), .B (n_99_38), .C1 (n_103_36), .C2 (n_106_36) );
AOI211_X1 g_87_44 (.ZN (n_87_44), .A (n_91_42), .B (n_97_39), .C1 (n_101_37), .C2 (n_104_37) );
AOI211_X1 g_85_45 (.ZN (n_85_45), .A (n_89_43), .B (n_95_40), .C1 (n_99_38), .C2 (n_105_35) );
AOI211_X1 g_83_46 (.ZN (n_83_46), .A (n_87_44), .B (n_93_41), .C1 (n_97_39), .C2 (n_103_36) );
AOI211_X1 g_81_47 (.ZN (n_81_47), .A (n_85_45), .B (n_91_42), .C1 (n_95_40), .C2 (n_101_37) );
AOI211_X1 g_79_48 (.ZN (n_79_48), .A (n_83_46), .B (n_89_43), .C1 (n_93_41), .C2 (n_99_38) );
AOI211_X1 g_77_49 (.ZN (n_77_49), .A (n_81_47), .B (n_87_44), .C1 (n_91_42), .C2 (n_97_39) );
AOI211_X1 g_75_50 (.ZN (n_75_50), .A (n_79_48), .B (n_85_45), .C1 (n_89_43), .C2 (n_95_40) );
AOI211_X1 g_73_51 (.ZN (n_73_51), .A (n_77_49), .B (n_83_46), .C1 (n_87_44), .C2 (n_93_41) );
AOI211_X1 g_71_52 (.ZN (n_71_52), .A (n_75_50), .B (n_81_47), .C1 (n_85_45), .C2 (n_91_42) );
AOI211_X1 g_69_53 (.ZN (n_69_53), .A (n_73_51), .B (n_79_48), .C1 (n_83_46), .C2 (n_89_43) );
AOI211_X1 g_67_54 (.ZN (n_67_54), .A (n_71_52), .B (n_77_49), .C1 (n_81_47), .C2 (n_87_44) );
AOI211_X1 g_65_55 (.ZN (n_65_55), .A (n_69_53), .B (n_75_50), .C1 (n_79_48), .C2 (n_85_45) );
AOI211_X1 g_63_56 (.ZN (n_63_56), .A (n_67_54), .B (n_73_51), .C1 (n_77_49), .C2 (n_83_46) );
AOI211_X1 g_61_57 (.ZN (n_61_57), .A (n_65_55), .B (n_71_52), .C1 (n_75_50), .C2 (n_81_47) );
AOI211_X1 g_59_58 (.ZN (n_59_58), .A (n_63_56), .B (n_69_53), .C1 (n_73_51), .C2 (n_79_48) );
AOI211_X1 g_57_59 (.ZN (n_57_59), .A (n_61_57), .B (n_67_54), .C1 (n_71_52), .C2 (n_77_49) );
AOI211_X1 g_55_60 (.ZN (n_55_60), .A (n_59_58), .B (n_65_55), .C1 (n_69_53), .C2 (n_75_50) );
AOI211_X1 g_53_61 (.ZN (n_53_61), .A (n_57_59), .B (n_63_56), .C1 (n_67_54), .C2 (n_73_51) );
AOI211_X1 g_51_62 (.ZN (n_51_62), .A (n_55_60), .B (n_61_57), .C1 (n_65_55), .C2 (n_71_52) );
AOI211_X1 g_49_63 (.ZN (n_49_63), .A (n_53_61), .B (n_59_58), .C1 (n_63_56), .C2 (n_69_53) );
AOI211_X1 g_47_64 (.ZN (n_47_64), .A (n_51_62), .B (n_57_59), .C1 (n_61_57), .C2 (n_67_54) );
AOI211_X1 g_45_65 (.ZN (n_45_65), .A (n_49_63), .B (n_55_60), .C1 (n_59_58), .C2 (n_65_55) );
AOI211_X1 g_43_66 (.ZN (n_43_66), .A (n_47_64), .B (n_53_61), .C1 (n_57_59), .C2 (n_63_56) );
AOI211_X1 g_41_67 (.ZN (n_41_67), .A (n_45_65), .B (n_51_62), .C1 (n_55_60), .C2 (n_61_57) );
AOI211_X1 g_39_68 (.ZN (n_39_68), .A (n_43_66), .B (n_49_63), .C1 (n_53_61), .C2 (n_59_58) );
AOI211_X1 g_37_69 (.ZN (n_37_69), .A (n_41_67), .B (n_47_64), .C1 (n_51_62), .C2 (n_57_59) );
AOI211_X1 g_35_70 (.ZN (n_35_70), .A (n_39_68), .B (n_45_65), .C1 (n_49_63), .C2 (n_55_60) );
AOI211_X1 g_33_71 (.ZN (n_33_71), .A (n_37_69), .B (n_43_66), .C1 (n_47_64), .C2 (n_53_61) );
AOI211_X1 g_31_72 (.ZN (n_31_72), .A (n_35_70), .B (n_41_67), .C1 (n_45_65), .C2 (n_51_62) );
AOI211_X1 g_29_73 (.ZN (n_29_73), .A (n_33_71), .B (n_39_68), .C1 (n_43_66), .C2 (n_49_63) );
AOI211_X1 g_27_72 (.ZN (n_27_72), .A (n_31_72), .B (n_37_69), .C1 (n_41_67), .C2 (n_47_64) );
AOI211_X1 g_25_73 (.ZN (n_25_73), .A (n_29_73), .B (n_35_70), .C1 (n_39_68), .C2 (n_45_65) );
AOI211_X1 g_23_74 (.ZN (n_23_74), .A (n_27_72), .B (n_33_71), .C1 (n_37_69), .C2 (n_43_66) );
AOI211_X1 g_21_75 (.ZN (n_21_75), .A (n_25_73), .B (n_31_72), .C1 (n_35_70), .C2 (n_41_67) );
AOI211_X1 g_19_76 (.ZN (n_19_76), .A (n_23_74), .B (n_29_73), .C1 (n_33_71), .C2 (n_39_68) );
AOI211_X1 g_17_77 (.ZN (n_17_77), .A (n_21_75), .B (n_27_72), .C1 (n_31_72), .C2 (n_37_69) );
AOI211_X1 g_15_78 (.ZN (n_15_78), .A (n_19_76), .B (n_25_73), .C1 (n_29_73), .C2 (n_35_70) );
AOI211_X1 g_13_79 (.ZN (n_13_79), .A (n_17_77), .B (n_23_74), .C1 (n_27_72), .C2 (n_33_71) );
AOI211_X1 g_11_80 (.ZN (n_11_80), .A (n_15_78), .B (n_21_75), .C1 (n_25_73), .C2 (n_31_72) );
AOI211_X1 g_9_81 (.ZN (n_9_81), .A (n_13_79), .B (n_19_76), .C1 (n_23_74), .C2 (n_29_73) );
AOI211_X1 g_8_83 (.ZN (n_8_83), .A (n_11_80), .B (n_17_77), .C1 (n_21_75), .C2 (n_27_72) );
AOI211_X1 g_10_82 (.ZN (n_10_82), .A (n_9_81), .B (n_15_78), .C1 (n_19_76), .C2 (n_25_73) );
AOI211_X1 g_12_81 (.ZN (n_12_81), .A (n_8_83), .B (n_13_79), .C1 (n_17_77), .C2 (n_23_74) );
AOI211_X1 g_14_80 (.ZN (n_14_80), .A (n_10_82), .B (n_11_80), .C1 (n_15_78), .C2 (n_21_75) );
AOI211_X1 g_16_79 (.ZN (n_16_79), .A (n_12_81), .B (n_9_81), .C1 (n_13_79), .C2 (n_19_76) );
AOI211_X1 g_18_78 (.ZN (n_18_78), .A (n_14_80), .B (n_8_83), .C1 (n_11_80), .C2 (n_17_77) );
AOI211_X1 g_20_77 (.ZN (n_20_77), .A (n_16_79), .B (n_10_82), .C1 (n_9_81), .C2 (n_15_78) );
AOI211_X1 g_22_76 (.ZN (n_22_76), .A (n_18_78), .B (n_12_81), .C1 (n_8_83), .C2 (n_13_79) );
AOI211_X1 g_24_75 (.ZN (n_24_75), .A (n_20_77), .B (n_14_80), .C1 (n_10_82), .C2 (n_11_80) );
AOI211_X1 g_26_74 (.ZN (n_26_74), .A (n_22_76), .B (n_16_79), .C1 (n_12_81), .C2 (n_9_81) );
AOI211_X1 g_28_73 (.ZN (n_28_73), .A (n_24_75), .B (n_18_78), .C1 (n_14_80), .C2 (n_8_83) );
AOI211_X1 g_30_72 (.ZN (n_30_72), .A (n_26_74), .B (n_20_77), .C1 (n_16_79), .C2 (n_10_82) );
AOI211_X1 g_32_71 (.ZN (n_32_71), .A (n_28_73), .B (n_22_76), .C1 (n_18_78), .C2 (n_12_81) );
AOI211_X1 g_34_70 (.ZN (n_34_70), .A (n_30_72), .B (n_24_75), .C1 (n_20_77), .C2 (n_14_80) );
AOI211_X1 g_36_69 (.ZN (n_36_69), .A (n_32_71), .B (n_26_74), .C1 (n_22_76), .C2 (n_16_79) );
AOI211_X1 g_38_68 (.ZN (n_38_68), .A (n_34_70), .B (n_28_73), .C1 (n_24_75), .C2 (n_18_78) );
AOI211_X1 g_40_67 (.ZN (n_40_67), .A (n_36_69), .B (n_30_72), .C1 (n_26_74), .C2 (n_20_77) );
AOI211_X1 g_42_66 (.ZN (n_42_66), .A (n_38_68), .B (n_32_71), .C1 (n_28_73), .C2 (n_22_76) );
AOI211_X1 g_41_68 (.ZN (n_41_68), .A (n_40_67), .B (n_34_70), .C1 (n_30_72), .C2 (n_24_75) );
AOI211_X1 g_43_67 (.ZN (n_43_67), .A (n_42_66), .B (n_36_69), .C1 (n_32_71), .C2 (n_26_74) );
AOI211_X1 g_45_66 (.ZN (n_45_66), .A (n_41_68), .B (n_38_68), .C1 (n_34_70), .C2 (n_28_73) );
AOI211_X1 g_47_65 (.ZN (n_47_65), .A (n_43_67), .B (n_40_67), .C1 (n_36_69), .C2 (n_30_72) );
AOI211_X1 g_49_64 (.ZN (n_49_64), .A (n_45_66), .B (n_42_66), .C1 (n_38_68), .C2 (n_32_71) );
AOI211_X1 g_51_63 (.ZN (n_51_63), .A (n_47_65), .B (n_41_68), .C1 (n_40_67), .C2 (n_34_70) );
AOI211_X1 g_53_62 (.ZN (n_53_62), .A (n_49_64), .B (n_43_67), .C1 (n_42_66), .C2 (n_36_69) );
AOI211_X1 g_55_61 (.ZN (n_55_61), .A (n_51_63), .B (n_45_66), .C1 (n_41_68), .C2 (n_38_68) );
AOI211_X1 g_56_59 (.ZN (n_56_59), .A (n_53_62), .B (n_47_65), .C1 (n_43_67), .C2 (n_40_67) );
AOI211_X1 g_58_58 (.ZN (n_58_58), .A (n_55_61), .B (n_49_64), .C1 (n_45_66), .C2 (n_42_66) );
AOI211_X1 g_60_57 (.ZN (n_60_57), .A (n_56_59), .B (n_51_63), .C1 (n_47_65), .C2 (n_41_68) );
AOI211_X1 g_62_56 (.ZN (n_62_56), .A (n_58_58), .B (n_53_62), .C1 (n_49_64), .C2 (n_43_67) );
AOI211_X1 g_64_55 (.ZN (n_64_55), .A (n_60_57), .B (n_55_61), .C1 (n_51_63), .C2 (n_45_66) );
AOI211_X1 g_66_54 (.ZN (n_66_54), .A (n_62_56), .B (n_56_59), .C1 (n_53_62), .C2 (n_47_65) );
AOI211_X1 g_68_53 (.ZN (n_68_53), .A (n_64_55), .B (n_58_58), .C1 (n_55_61), .C2 (n_49_64) );
AOI211_X1 g_70_52 (.ZN (n_70_52), .A (n_66_54), .B (n_60_57), .C1 (n_56_59), .C2 (n_51_63) );
AOI211_X1 g_69_54 (.ZN (n_69_54), .A (n_68_53), .B (n_62_56), .C1 (n_58_58), .C2 (n_53_62) );
AOI211_X1 g_71_53 (.ZN (n_71_53), .A (n_70_52), .B (n_64_55), .C1 (n_60_57), .C2 (n_55_61) );
AOI211_X1 g_73_52 (.ZN (n_73_52), .A (n_69_54), .B (n_66_54), .C1 (n_62_56), .C2 (n_56_59) );
AOI211_X1 g_75_51 (.ZN (n_75_51), .A (n_71_53), .B (n_68_53), .C1 (n_64_55), .C2 (n_58_58) );
AOI211_X1 g_77_50 (.ZN (n_77_50), .A (n_73_52), .B (n_70_52), .C1 (n_66_54), .C2 (n_60_57) );
AOI211_X1 g_79_49 (.ZN (n_79_49), .A (n_75_51), .B (n_69_54), .C1 (n_68_53), .C2 (n_62_56) );
AOI211_X1 g_81_48 (.ZN (n_81_48), .A (n_77_50), .B (n_71_53), .C1 (n_70_52), .C2 (n_64_55) );
AOI211_X1 g_83_47 (.ZN (n_83_47), .A (n_79_49), .B (n_73_52), .C1 (n_69_54), .C2 (n_66_54) );
AOI211_X1 g_85_46 (.ZN (n_85_46), .A (n_81_48), .B (n_75_51), .C1 (n_71_53), .C2 (n_68_53) );
AOI211_X1 g_87_45 (.ZN (n_87_45), .A (n_83_47), .B (n_77_50), .C1 (n_73_52), .C2 (n_70_52) );
AOI211_X1 g_89_44 (.ZN (n_89_44), .A (n_85_46), .B (n_79_49), .C1 (n_75_51), .C2 (n_69_54) );
AOI211_X1 g_91_43 (.ZN (n_91_43), .A (n_87_45), .B (n_81_48), .C1 (n_77_50), .C2 (n_71_53) );
AOI211_X1 g_93_42 (.ZN (n_93_42), .A (n_89_44), .B (n_83_47), .C1 (n_79_49), .C2 (n_73_52) );
AOI211_X1 g_95_41 (.ZN (n_95_41), .A (n_91_43), .B (n_85_46), .C1 (n_81_48), .C2 (n_75_51) );
AOI211_X1 g_97_40 (.ZN (n_97_40), .A (n_93_42), .B (n_87_45), .C1 (n_83_47), .C2 (n_77_50) );
AOI211_X1 g_99_39 (.ZN (n_99_39), .A (n_95_41), .B (n_89_44), .C1 (n_85_46), .C2 (n_79_49) );
AOI211_X1 g_101_38 (.ZN (n_101_38), .A (n_97_40), .B (n_91_43), .C1 (n_87_45), .C2 (n_81_48) );
AOI211_X1 g_103_37 (.ZN (n_103_37), .A (n_99_39), .B (n_93_42), .C1 (n_89_44), .C2 (n_83_47) );
AOI211_X1 g_105_36 (.ZN (n_105_36), .A (n_101_38), .B (n_95_41), .C1 (n_91_43), .C2 (n_85_46) );
AOI211_X1 g_107_35 (.ZN (n_107_35), .A (n_103_37), .B (n_97_40), .C1 (n_93_42), .C2 (n_87_45) );
AOI211_X1 g_109_34 (.ZN (n_109_34), .A (n_105_36), .B (n_99_39), .C1 (n_95_41), .C2 (n_89_44) );
AOI211_X1 g_108_36 (.ZN (n_108_36), .A (n_107_35), .B (n_101_38), .C1 (n_97_40), .C2 (n_91_43) );
AOI211_X1 g_106_35 (.ZN (n_106_35), .A (n_109_34), .B (n_103_37), .C1 (n_99_39), .C2 (n_93_42) );
AOI211_X1 g_108_34 (.ZN (n_108_34), .A (n_108_36), .B (n_105_36), .C1 (n_101_38), .C2 (n_95_41) );
AOI211_X1 g_110_33 (.ZN (n_110_33), .A (n_106_35), .B (n_107_35), .C1 (n_103_37), .C2 (n_97_40) );
AOI211_X1 g_112_32 (.ZN (n_112_32), .A (n_108_34), .B (n_109_34), .C1 (n_105_36), .C2 (n_99_39) );
AOI211_X1 g_114_31 (.ZN (n_114_31), .A (n_110_33), .B (n_108_36), .C1 (n_107_35), .C2 (n_101_38) );
AOI211_X1 g_116_30 (.ZN (n_116_30), .A (n_112_32), .B (n_106_35), .C1 (n_109_34), .C2 (n_103_37) );
AOI211_X1 g_115_32 (.ZN (n_115_32), .A (n_114_31), .B (n_108_34), .C1 (n_108_36), .C2 (n_105_36) );
AOI211_X1 g_113_33 (.ZN (n_113_33), .A (n_116_30), .B (n_110_33), .C1 (n_106_35), .C2 (n_107_35) );
AOI211_X1 g_111_34 (.ZN (n_111_34), .A (n_115_32), .B (n_112_32), .C1 (n_108_34), .C2 (n_109_34) );
AOI211_X1 g_109_35 (.ZN (n_109_35), .A (n_113_33), .B (n_114_31), .C1 (n_110_33), .C2 (n_108_36) );
AOI211_X1 g_107_36 (.ZN (n_107_36), .A (n_111_34), .B (n_116_30), .C1 (n_112_32), .C2 (n_106_35) );
AOI211_X1 g_105_37 (.ZN (n_105_37), .A (n_109_35), .B (n_115_32), .C1 (n_114_31), .C2 (n_108_34) );
AOI211_X1 g_103_38 (.ZN (n_103_38), .A (n_107_36), .B (n_113_33), .C1 (n_116_30), .C2 (n_110_33) );
AOI211_X1 g_104_36 (.ZN (n_104_36), .A (n_105_37), .B (n_111_34), .C1 (n_115_32), .C2 (n_112_32) );
AOI211_X1 g_102_37 (.ZN (n_102_37), .A (n_103_38), .B (n_109_35), .C1 (n_113_33), .C2 (n_114_31) );
AOI211_X1 g_100_38 (.ZN (n_100_38), .A (n_104_36), .B (n_107_36), .C1 (n_111_34), .C2 (n_116_30) );
AOI211_X1 g_98_39 (.ZN (n_98_39), .A (n_102_37), .B (n_105_37), .C1 (n_109_35), .C2 (n_115_32) );
AOI211_X1 g_96_40 (.ZN (n_96_40), .A (n_100_38), .B (n_103_38), .C1 (n_107_36), .C2 (n_113_33) );
AOI211_X1 g_94_41 (.ZN (n_94_41), .A (n_98_39), .B (n_104_36), .C1 (n_105_37), .C2 (n_111_34) );
AOI211_X1 g_92_42 (.ZN (n_92_42), .A (n_96_40), .B (n_102_37), .C1 (n_103_38), .C2 (n_109_35) );
AOI211_X1 g_90_43 (.ZN (n_90_43), .A (n_94_41), .B (n_100_38), .C1 (n_104_36), .C2 (n_107_36) );
AOI211_X1 g_88_44 (.ZN (n_88_44), .A (n_92_42), .B (n_98_39), .C1 (n_102_37), .C2 (n_105_37) );
AOI211_X1 g_86_45 (.ZN (n_86_45), .A (n_90_43), .B (n_96_40), .C1 (n_100_38), .C2 (n_103_38) );
AOI211_X1 g_84_46 (.ZN (n_84_46), .A (n_88_44), .B (n_94_41), .C1 (n_98_39), .C2 (n_104_36) );
AOI211_X1 g_82_47 (.ZN (n_82_47), .A (n_86_45), .B (n_92_42), .C1 (n_96_40), .C2 (n_102_37) );
AOI211_X1 g_80_48 (.ZN (n_80_48), .A (n_84_46), .B (n_90_43), .C1 (n_94_41), .C2 (n_100_38) );
AOI211_X1 g_78_49 (.ZN (n_78_49), .A (n_82_47), .B (n_88_44), .C1 (n_92_42), .C2 (n_98_39) );
AOI211_X1 g_76_50 (.ZN (n_76_50), .A (n_80_48), .B (n_86_45), .C1 (n_90_43), .C2 (n_96_40) );
AOI211_X1 g_74_51 (.ZN (n_74_51), .A (n_78_49), .B (n_84_46), .C1 (n_88_44), .C2 (n_94_41) );
AOI211_X1 g_72_52 (.ZN (n_72_52), .A (n_76_50), .B (n_82_47), .C1 (n_86_45), .C2 (n_92_42) );
AOI211_X1 g_70_53 (.ZN (n_70_53), .A (n_74_51), .B (n_80_48), .C1 (n_84_46), .C2 (n_90_43) );
AOI211_X1 g_68_54 (.ZN (n_68_54), .A (n_72_52), .B (n_78_49), .C1 (n_82_47), .C2 (n_88_44) );
AOI211_X1 g_66_55 (.ZN (n_66_55), .A (n_70_53), .B (n_76_50), .C1 (n_80_48), .C2 (n_86_45) );
AOI211_X1 g_64_56 (.ZN (n_64_56), .A (n_68_54), .B (n_74_51), .C1 (n_78_49), .C2 (n_84_46) );
AOI211_X1 g_62_57 (.ZN (n_62_57), .A (n_66_55), .B (n_72_52), .C1 (n_76_50), .C2 (n_82_47) );
AOI211_X1 g_60_58 (.ZN (n_60_58), .A (n_64_56), .B (n_70_53), .C1 (n_74_51), .C2 (n_80_48) );
AOI211_X1 g_58_59 (.ZN (n_58_59), .A (n_62_57), .B (n_68_54), .C1 (n_72_52), .C2 (n_78_49) );
AOI211_X1 g_56_60 (.ZN (n_56_60), .A (n_60_58), .B (n_66_55), .C1 (n_70_53), .C2 (n_76_50) );
AOI211_X1 g_54_61 (.ZN (n_54_61), .A (n_58_59), .B (n_64_56), .C1 (n_68_54), .C2 (n_74_51) );
AOI211_X1 g_52_62 (.ZN (n_52_62), .A (n_56_60), .B (n_62_57), .C1 (n_66_55), .C2 (n_72_52) );
AOI211_X1 g_50_63 (.ZN (n_50_63), .A (n_54_61), .B (n_60_58), .C1 (n_64_56), .C2 (n_70_53) );
AOI211_X1 g_48_64 (.ZN (n_48_64), .A (n_52_62), .B (n_58_59), .C1 (n_62_57), .C2 (n_68_54) );
AOI211_X1 g_46_65 (.ZN (n_46_65), .A (n_50_63), .B (n_56_60), .C1 (n_60_58), .C2 (n_66_55) );
AOI211_X1 g_44_66 (.ZN (n_44_66), .A (n_48_64), .B (n_54_61), .C1 (n_58_59), .C2 (n_64_56) );
AOI211_X1 g_42_67 (.ZN (n_42_67), .A (n_46_65), .B (n_52_62), .C1 (n_56_60), .C2 (n_62_57) );
AOI211_X1 g_40_68 (.ZN (n_40_68), .A (n_44_66), .B (n_50_63), .C1 (n_54_61), .C2 (n_60_58) );
AOI211_X1 g_38_69 (.ZN (n_38_69), .A (n_42_67), .B (n_48_64), .C1 (n_52_62), .C2 (n_58_59) );
AOI211_X1 g_36_70 (.ZN (n_36_70), .A (n_40_68), .B (n_46_65), .C1 (n_50_63), .C2 (n_56_60) );
AOI211_X1 g_34_71 (.ZN (n_34_71), .A (n_38_69), .B (n_44_66), .C1 (n_48_64), .C2 (n_54_61) );
AOI211_X1 g_32_72 (.ZN (n_32_72), .A (n_36_70), .B (n_42_67), .C1 (n_46_65), .C2 (n_52_62) );
AOI211_X1 g_30_73 (.ZN (n_30_73), .A (n_34_71), .B (n_40_68), .C1 (n_44_66), .C2 (n_50_63) );
AOI211_X1 g_28_74 (.ZN (n_28_74), .A (n_32_72), .B (n_38_69), .C1 (n_42_67), .C2 (n_48_64) );
AOI211_X1 g_26_75 (.ZN (n_26_75), .A (n_30_73), .B (n_36_70), .C1 (n_40_68), .C2 (n_46_65) );
AOI211_X1 g_24_76 (.ZN (n_24_76), .A (n_28_74), .B (n_34_71), .C1 (n_38_69), .C2 (n_44_66) );
AOI211_X1 g_22_77 (.ZN (n_22_77), .A (n_26_75), .B (n_32_72), .C1 (n_36_70), .C2 (n_42_67) );
AOI211_X1 g_21_79 (.ZN (n_21_79), .A (n_24_76), .B (n_30_73), .C1 (n_34_71), .C2 (n_40_68) );
AOI211_X1 g_19_78 (.ZN (n_19_78), .A (n_22_77), .B (n_28_74), .C1 (n_32_72), .C2 (n_38_69) );
AOI211_X1 g_21_77 (.ZN (n_21_77), .A (n_21_79), .B (n_26_75), .C1 (n_30_73), .C2 (n_36_70) );
AOI211_X1 g_23_76 (.ZN (n_23_76), .A (n_19_78), .B (n_24_76), .C1 (n_28_74), .C2 (n_34_71) );
AOI211_X1 g_25_75 (.ZN (n_25_75), .A (n_21_77), .B (n_22_77), .C1 (n_26_75), .C2 (n_32_72) );
AOI211_X1 g_27_74 (.ZN (n_27_74), .A (n_23_76), .B (n_21_79), .C1 (n_24_76), .C2 (n_30_73) );
AOI211_X1 g_26_76 (.ZN (n_26_76), .A (n_25_75), .B (n_19_78), .C1 (n_22_77), .C2 (n_28_74) );
AOI211_X1 g_28_75 (.ZN (n_28_75), .A (n_27_74), .B (n_21_77), .C1 (n_21_79), .C2 (n_26_75) );
AOI211_X1 g_30_74 (.ZN (n_30_74), .A (n_26_76), .B (n_23_76), .C1 (n_19_78), .C2 (n_24_76) );
AOI211_X1 g_32_73 (.ZN (n_32_73), .A (n_28_75), .B (n_25_75), .C1 (n_21_77), .C2 (n_22_77) );
AOI211_X1 g_34_72 (.ZN (n_34_72), .A (n_30_74), .B (n_27_74), .C1 (n_23_76), .C2 (n_21_79) );
AOI211_X1 g_36_71 (.ZN (n_36_71), .A (n_32_73), .B (n_26_76), .C1 (n_25_75), .C2 (n_19_78) );
AOI211_X1 g_38_70 (.ZN (n_38_70), .A (n_34_72), .B (n_28_75), .C1 (n_27_74), .C2 (n_21_77) );
AOI211_X1 g_40_69 (.ZN (n_40_69), .A (n_36_71), .B (n_30_74), .C1 (n_26_76), .C2 (n_23_76) );
AOI211_X1 g_42_68 (.ZN (n_42_68), .A (n_38_70), .B (n_32_73), .C1 (n_28_75), .C2 (n_25_75) );
AOI211_X1 g_44_67 (.ZN (n_44_67), .A (n_40_69), .B (n_34_72), .C1 (n_30_74), .C2 (n_27_74) );
AOI211_X1 g_46_66 (.ZN (n_46_66), .A (n_42_68), .B (n_36_71), .C1 (n_32_73), .C2 (n_26_76) );
AOI211_X1 g_48_65 (.ZN (n_48_65), .A (n_44_67), .B (n_38_70), .C1 (n_34_72), .C2 (n_28_75) );
AOI211_X1 g_50_64 (.ZN (n_50_64), .A (n_46_66), .B (n_40_69), .C1 (n_36_71), .C2 (n_30_74) );
AOI211_X1 g_52_63 (.ZN (n_52_63), .A (n_48_65), .B (n_42_68), .C1 (n_38_70), .C2 (n_32_73) );
AOI211_X1 g_54_62 (.ZN (n_54_62), .A (n_50_64), .B (n_44_67), .C1 (n_40_69), .C2 (n_34_72) );
AOI211_X1 g_56_61 (.ZN (n_56_61), .A (n_52_63), .B (n_46_66), .C1 (n_42_68), .C2 (n_36_71) );
AOI211_X1 g_58_60 (.ZN (n_58_60), .A (n_54_62), .B (n_48_65), .C1 (n_44_67), .C2 (n_38_70) );
AOI211_X1 g_60_59 (.ZN (n_60_59), .A (n_56_61), .B (n_50_64), .C1 (n_46_66), .C2 (n_40_69) );
AOI211_X1 g_62_58 (.ZN (n_62_58), .A (n_58_60), .B (n_52_63), .C1 (n_48_65), .C2 (n_42_68) );
AOI211_X1 g_64_57 (.ZN (n_64_57), .A (n_60_59), .B (n_54_62), .C1 (n_50_64), .C2 (n_44_67) );
AOI211_X1 g_66_56 (.ZN (n_66_56), .A (n_62_58), .B (n_56_61), .C1 (n_52_63), .C2 (n_46_66) );
AOI211_X1 g_68_55 (.ZN (n_68_55), .A (n_64_57), .B (n_58_60), .C1 (n_54_62), .C2 (n_48_65) );
AOI211_X1 g_70_54 (.ZN (n_70_54), .A (n_66_56), .B (n_60_59), .C1 (n_56_61), .C2 (n_50_64) );
AOI211_X1 g_72_53 (.ZN (n_72_53), .A (n_68_55), .B (n_62_58), .C1 (n_58_60), .C2 (n_52_63) );
AOI211_X1 g_74_52 (.ZN (n_74_52), .A (n_70_54), .B (n_64_57), .C1 (n_60_59), .C2 (n_54_62) );
AOI211_X1 g_76_51 (.ZN (n_76_51), .A (n_72_53), .B (n_66_56), .C1 (n_62_58), .C2 (n_56_61) );
AOI211_X1 g_78_50 (.ZN (n_78_50), .A (n_74_52), .B (n_68_55), .C1 (n_64_57), .C2 (n_58_60) );
AOI211_X1 g_80_49 (.ZN (n_80_49), .A (n_76_51), .B (n_70_54), .C1 (n_66_56), .C2 (n_60_59) );
AOI211_X1 g_82_48 (.ZN (n_82_48), .A (n_78_50), .B (n_72_53), .C1 (n_68_55), .C2 (n_62_58) );
AOI211_X1 g_84_47 (.ZN (n_84_47), .A (n_80_49), .B (n_74_52), .C1 (n_70_54), .C2 (n_64_57) );
AOI211_X1 g_86_46 (.ZN (n_86_46), .A (n_82_48), .B (n_76_51), .C1 (n_72_53), .C2 (n_66_56) );
AOI211_X1 g_88_45 (.ZN (n_88_45), .A (n_84_47), .B (n_78_50), .C1 (n_74_52), .C2 (n_68_55) );
AOI211_X1 g_90_44 (.ZN (n_90_44), .A (n_86_46), .B (n_80_49), .C1 (n_76_51), .C2 (n_70_54) );
AOI211_X1 g_92_43 (.ZN (n_92_43), .A (n_88_45), .B (n_82_48), .C1 (n_78_50), .C2 (n_72_53) );
AOI211_X1 g_94_42 (.ZN (n_94_42), .A (n_90_44), .B (n_84_47), .C1 (n_80_49), .C2 (n_74_52) );
AOI211_X1 g_96_41 (.ZN (n_96_41), .A (n_92_43), .B (n_86_46), .C1 (n_82_48), .C2 (n_76_51) );
AOI211_X1 g_98_40 (.ZN (n_98_40), .A (n_94_42), .B (n_88_45), .C1 (n_84_47), .C2 (n_78_50) );
AOI211_X1 g_100_39 (.ZN (n_100_39), .A (n_96_41), .B (n_90_44), .C1 (n_86_46), .C2 (n_80_49) );
AOI211_X1 g_102_38 (.ZN (n_102_38), .A (n_98_40), .B (n_92_43), .C1 (n_88_45), .C2 (n_82_48) );
AOI211_X1 g_101_40 (.ZN (n_101_40), .A (n_100_39), .B (n_94_42), .C1 (n_90_44), .C2 (n_84_47) );
AOI211_X1 g_103_39 (.ZN (n_103_39), .A (n_102_38), .B (n_96_41), .C1 (n_92_43), .C2 (n_86_46) );
AOI211_X1 g_105_38 (.ZN (n_105_38), .A (n_101_40), .B (n_98_40), .C1 (n_94_42), .C2 (n_88_45) );
AOI211_X1 g_107_37 (.ZN (n_107_37), .A (n_103_39), .B (n_100_39), .C1 (n_96_41), .C2 (n_90_44) );
AOI211_X1 g_109_36 (.ZN (n_109_36), .A (n_105_38), .B (n_102_38), .C1 (n_98_40), .C2 (n_92_43) );
AOI211_X1 g_111_35 (.ZN (n_111_35), .A (n_107_37), .B (n_101_40), .C1 (n_100_39), .C2 (n_94_42) );
AOI211_X1 g_113_34 (.ZN (n_113_34), .A (n_109_36), .B (n_103_39), .C1 (n_102_38), .C2 (n_96_41) );
AOI211_X1 g_115_33 (.ZN (n_115_33), .A (n_111_35), .B (n_105_38), .C1 (n_101_40), .C2 (n_98_40) );
AOI211_X1 g_117_32 (.ZN (n_117_32), .A (n_113_34), .B (n_107_37), .C1 (n_103_39), .C2 (n_100_39) );
AOI211_X1 g_119_31 (.ZN (n_119_31), .A (n_115_33), .B (n_109_36), .C1 (n_105_38), .C2 (n_102_38) );
AOI211_X1 g_118_33 (.ZN (n_118_33), .A (n_117_32), .B (n_111_35), .C1 (n_107_37), .C2 (n_101_40) );
AOI211_X1 g_116_32 (.ZN (n_116_32), .A (n_119_31), .B (n_113_34), .C1 (n_109_36), .C2 (n_103_39) );
AOI211_X1 g_118_31 (.ZN (n_118_31), .A (n_118_33), .B (n_115_33), .C1 (n_111_35), .C2 (n_105_38) );
AOI211_X1 g_117_33 (.ZN (n_117_33), .A (n_116_32), .B (n_117_32), .C1 (n_113_34), .C2 (n_107_37) );
AOI211_X1 g_115_34 (.ZN (n_115_34), .A (n_118_31), .B (n_119_31), .C1 (n_115_33), .C2 (n_109_36) );
AOI211_X1 g_113_35 (.ZN (n_113_35), .A (n_117_33), .B (n_118_33), .C1 (n_117_32), .C2 (n_111_35) );
AOI211_X1 g_114_33 (.ZN (n_114_33), .A (n_115_34), .B (n_116_32), .C1 (n_119_31), .C2 (n_113_34) );
AOI211_X1 g_112_34 (.ZN (n_112_34), .A (n_113_35), .B (n_118_31), .C1 (n_118_33), .C2 (n_115_33) );
AOI211_X1 g_110_35 (.ZN (n_110_35), .A (n_114_33), .B (n_117_33), .C1 (n_116_32), .C2 (n_117_32) );
AOI211_X1 g_109_37 (.ZN (n_109_37), .A (n_112_34), .B (n_115_34), .C1 (n_118_31), .C2 (n_119_31) );
AOI211_X1 g_111_36 (.ZN (n_111_36), .A (n_110_35), .B (n_113_35), .C1 (n_117_33), .C2 (n_118_33) );
AOI211_X1 g_110_38 (.ZN (n_110_38), .A (n_109_37), .B (n_114_33), .C1 (n_115_34), .C2 (n_116_32) );
AOI211_X1 g_108_37 (.ZN (n_108_37), .A (n_111_36), .B (n_112_34), .C1 (n_113_35), .C2 (n_118_31) );
AOI211_X1 g_110_36 (.ZN (n_110_36), .A (n_110_38), .B (n_110_35), .C1 (n_114_33), .C2 (n_117_33) );
AOI211_X1 g_112_35 (.ZN (n_112_35), .A (n_108_37), .B (n_109_37), .C1 (n_112_34), .C2 (n_115_34) );
AOI211_X1 g_114_34 (.ZN (n_114_34), .A (n_110_36), .B (n_111_36), .C1 (n_110_35), .C2 (n_113_35) );
AOI211_X1 g_116_33 (.ZN (n_116_33), .A (n_112_35), .B (n_110_38), .C1 (n_109_37), .C2 (n_114_33) );
AOI211_X1 g_118_32 (.ZN (n_118_32), .A (n_114_34), .B (n_108_37), .C1 (n_111_36), .C2 (n_112_34) );
AOI211_X1 g_120_31 (.ZN (n_120_31), .A (n_116_33), .B (n_110_36), .C1 (n_110_38), .C2 (n_110_35) );
AOI211_X1 g_122_30 (.ZN (n_122_30), .A (n_118_32), .B (n_112_35), .C1 (n_108_37), .C2 (n_109_37) );
AOI211_X1 g_124_29 (.ZN (n_124_29), .A (n_120_31), .B (n_114_34), .C1 (n_110_36), .C2 (n_111_36) );
AOI211_X1 g_126_28 (.ZN (n_126_28), .A (n_122_30), .B (n_116_33), .C1 (n_112_35), .C2 (n_110_38) );
AOI211_X1 g_125_30 (.ZN (n_125_30), .A (n_124_29), .B (n_118_32), .C1 (n_114_34), .C2 (n_108_37) );
AOI211_X1 g_127_29 (.ZN (n_127_29), .A (n_126_28), .B (n_120_31), .C1 (n_116_33), .C2 (n_110_36) );
AOI211_X1 g_129_28 (.ZN (n_129_28), .A (n_125_30), .B (n_122_30), .C1 (n_118_32), .C2 (n_112_35) );
AOI211_X1 g_131_27 (.ZN (n_131_27), .A (n_127_29), .B (n_124_29), .C1 (n_120_31), .C2 (n_114_34) );
AOI211_X1 g_133_26 (.ZN (n_133_26), .A (n_129_28), .B (n_126_28), .C1 (n_122_30), .C2 (n_116_33) );
AOI211_X1 g_135_25 (.ZN (n_135_25), .A (n_131_27), .B (n_125_30), .C1 (n_124_29), .C2 (n_118_32) );
AOI211_X1 g_137_24 (.ZN (n_137_24), .A (n_133_26), .B (n_127_29), .C1 (n_126_28), .C2 (n_120_31) );
AOI211_X1 g_136_22 (.ZN (n_136_22), .A (n_135_25), .B (n_129_28), .C1 (n_125_30), .C2 (n_122_30) );
AOI211_X1 g_138_21 (.ZN (n_138_21), .A (n_137_24), .B (n_131_27), .C1 (n_127_29), .C2 (n_124_29) );
AOI211_X1 g_140_20 (.ZN (n_140_20), .A (n_136_22), .B (n_133_26), .C1 (n_129_28), .C2 (n_126_28) );
AOI211_X1 g_139_22 (.ZN (n_139_22), .A (n_138_21), .B (n_135_25), .C1 (n_131_27), .C2 (n_125_30) );
AOI211_X1 g_137_23 (.ZN (n_137_23), .A (n_140_20), .B (n_137_24), .C1 (n_133_26), .C2 (n_127_29) );
AOI211_X1 g_135_24 (.ZN (n_135_24), .A (n_139_22), .B (n_136_22), .C1 (n_135_25), .C2 (n_129_28) );
AOI211_X1 g_133_25 (.ZN (n_133_25), .A (n_137_23), .B (n_138_21), .C1 (n_137_24), .C2 (n_131_27) );
AOI211_X1 g_131_26 (.ZN (n_131_26), .A (n_135_24), .B (n_140_20), .C1 (n_136_22), .C2 (n_133_26) );
AOI211_X1 g_129_27 (.ZN (n_129_27), .A (n_133_25), .B (n_139_22), .C1 (n_138_21), .C2 (n_135_25) );
AOI211_X1 g_127_28 (.ZN (n_127_28), .A (n_131_26), .B (n_137_23), .C1 (n_140_20), .C2 (n_137_24) );
AOI211_X1 g_125_29 (.ZN (n_125_29), .A (n_129_27), .B (n_135_24), .C1 (n_139_22), .C2 (n_136_22) );
AOI211_X1 g_123_30 (.ZN (n_123_30), .A (n_127_28), .B (n_133_25), .C1 (n_137_23), .C2 (n_138_21) );
AOI211_X1 g_122_32 (.ZN (n_122_32), .A (n_125_29), .B (n_131_26), .C1 (n_135_24), .C2 (n_140_20) );
AOI211_X1 g_124_31 (.ZN (n_124_31), .A (n_123_30), .B (n_129_27), .C1 (n_133_25), .C2 (n_139_22) );
AOI211_X1 g_126_30 (.ZN (n_126_30), .A (n_122_32), .B (n_127_28), .C1 (n_131_26), .C2 (n_137_23) );
AOI211_X1 g_128_29 (.ZN (n_128_29), .A (n_124_31), .B (n_125_29), .C1 (n_129_27), .C2 (n_135_24) );
AOI211_X1 g_130_28 (.ZN (n_130_28), .A (n_126_30), .B (n_123_30), .C1 (n_127_28), .C2 (n_133_25) );
AOI211_X1 g_132_27 (.ZN (n_132_27), .A (n_128_29), .B (n_122_32), .C1 (n_125_29), .C2 (n_131_26) );
AOI211_X1 g_134_26 (.ZN (n_134_26), .A (n_130_28), .B (n_124_31), .C1 (n_123_30), .C2 (n_129_27) );
AOI211_X1 g_136_25 (.ZN (n_136_25), .A (n_132_27), .B (n_126_30), .C1 (n_122_32), .C2 (n_127_28) );
AOI211_X1 g_135_27 (.ZN (n_135_27), .A (n_134_26), .B (n_128_29), .C1 (n_124_31), .C2 (n_125_29) );
AOI211_X1 g_133_28 (.ZN (n_133_28), .A (n_136_25), .B (n_130_28), .C1 (n_126_30), .C2 (n_123_30) );
AOI211_X1 g_131_29 (.ZN (n_131_29), .A (n_135_27), .B (n_132_27), .C1 (n_128_29), .C2 (n_122_32) );
AOI211_X1 g_129_30 (.ZN (n_129_30), .A (n_133_28), .B (n_134_26), .C1 (n_130_28), .C2 (n_124_31) );
AOI211_X1 g_128_28 (.ZN (n_128_28), .A (n_131_29), .B (n_136_25), .C1 (n_132_27), .C2 (n_126_30) );
AOI211_X1 g_126_29 (.ZN (n_126_29), .A (n_129_30), .B (n_135_27), .C1 (n_134_26), .C2 (n_128_29) );
AOI211_X1 g_124_30 (.ZN (n_124_30), .A (n_128_28), .B (n_133_28), .C1 (n_136_25), .C2 (n_130_28) );
AOI211_X1 g_122_31 (.ZN (n_122_31), .A (n_126_29), .B (n_131_29), .C1 (n_135_27), .C2 (n_132_27) );
AOI211_X1 g_120_32 (.ZN (n_120_32), .A (n_124_30), .B (n_129_30), .C1 (n_133_28), .C2 (n_134_26) );
AOI211_X1 g_119_34 (.ZN (n_119_34), .A (n_122_31), .B (n_128_28), .C1 (n_131_29), .C2 (n_136_25) );
AOI211_X1 g_121_33 (.ZN (n_121_33), .A (n_120_32), .B (n_126_29), .C1 (n_129_30), .C2 (n_135_27) );
AOI211_X1 g_123_32 (.ZN (n_123_32), .A (n_119_34), .B (n_124_30), .C1 (n_128_28), .C2 (n_133_28) );
AOI211_X1 g_125_31 (.ZN (n_125_31), .A (n_121_33), .B (n_122_31), .C1 (n_126_29), .C2 (n_131_29) );
AOI211_X1 g_127_30 (.ZN (n_127_30), .A (n_123_32), .B (n_120_32), .C1 (n_124_30), .C2 (n_129_30) );
AOI211_X1 g_129_29 (.ZN (n_129_29), .A (n_125_31), .B (n_119_34), .C1 (n_122_31), .C2 (n_128_28) );
AOI211_X1 g_131_28 (.ZN (n_131_28), .A (n_127_30), .B (n_121_33), .C1 (n_120_32), .C2 (n_126_29) );
AOI211_X1 g_133_27 (.ZN (n_133_27), .A (n_129_29), .B (n_123_32), .C1 (n_119_34), .C2 (n_124_30) );
AOI211_X1 g_135_26 (.ZN (n_135_26), .A (n_131_28), .B (n_125_31), .C1 (n_121_33), .C2 (n_122_31) );
AOI211_X1 g_136_24 (.ZN (n_136_24), .A (n_133_27), .B (n_127_30), .C1 (n_123_32), .C2 (n_120_32) );
AOI211_X1 g_138_23 (.ZN (n_138_23), .A (n_135_26), .B (n_129_29), .C1 (n_125_31), .C2 (n_119_34) );
AOI211_X1 g_140_22 (.ZN (n_140_22), .A (n_136_24), .B (n_131_28), .C1 (n_127_30), .C2 (n_121_33) );
AOI211_X1 g_142_21 (.ZN (n_142_21), .A (n_138_23), .B (n_133_27), .C1 (n_129_29), .C2 (n_123_32) );
AOI211_X1 g_141_23 (.ZN (n_141_23), .A (n_140_22), .B (n_135_26), .C1 (n_131_28), .C2 (n_125_31) );
AOI211_X1 g_139_24 (.ZN (n_139_24), .A (n_142_21), .B (n_136_24), .C1 (n_133_27), .C2 (n_127_30) );
AOI211_X1 g_137_25 (.ZN (n_137_25), .A (n_141_23), .B (n_138_23), .C1 (n_135_26), .C2 (n_129_29) );
AOI211_X1 g_136_27 (.ZN (n_136_27), .A (n_139_24), .B (n_140_22), .C1 (n_136_24), .C2 (n_131_28) );
AOI211_X1 g_138_26 (.ZN (n_138_26), .A (n_137_25), .B (n_142_21), .C1 (n_138_23), .C2 (n_133_27) );
AOI211_X1 g_140_25 (.ZN (n_140_25), .A (n_136_27), .B (n_141_23), .C1 (n_140_22), .C2 (n_135_26) );
AOI211_X1 g_139_23 (.ZN (n_139_23), .A (n_138_26), .B (n_139_24), .C1 (n_142_21), .C2 (n_136_24) );
AOI211_X1 g_141_22 (.ZN (n_141_22), .A (n_140_25), .B (n_137_25), .C1 (n_141_23), .C2 (n_138_23) );
AOI211_X1 g_143_21 (.ZN (n_143_21), .A (n_139_23), .B (n_136_27), .C1 (n_139_24), .C2 (n_140_22) );
AOI211_X1 g_145_20 (.ZN (n_145_20), .A (n_141_22), .B (n_138_26), .C1 (n_137_25), .C2 (n_142_21) );
AOI211_X1 g_147_21 (.ZN (n_147_21), .A (n_143_21), .B (n_140_25), .C1 (n_136_27), .C2 (n_141_23) );
AOI211_X1 g_145_22 (.ZN (n_145_22), .A (n_145_20), .B (n_139_23), .C1 (n_138_26), .C2 (n_139_24) );
AOI211_X1 g_143_23 (.ZN (n_143_23), .A (n_147_21), .B (n_141_22), .C1 (n_140_25), .C2 (n_137_25) );
AOI211_X1 g_141_24 (.ZN (n_141_24), .A (n_145_22), .B (n_143_21), .C1 (n_139_23), .C2 (n_136_27) );
AOI211_X1 g_139_25 (.ZN (n_139_25), .A (n_143_23), .B (n_145_20), .C1 (n_141_22), .C2 (n_138_26) );
AOI211_X1 g_137_26 (.ZN (n_137_26), .A (n_141_24), .B (n_147_21), .C1 (n_143_21), .C2 (n_140_25) );
AOI211_X1 g_136_28 (.ZN (n_136_28), .A (n_139_25), .B (n_145_22), .C1 (n_145_20), .C2 (n_139_23) );
AOI211_X1 g_134_27 (.ZN (n_134_27), .A (n_137_26), .B (n_143_23), .C1 (n_147_21), .C2 (n_141_22) );
AOI211_X1 g_136_26 (.ZN (n_136_26), .A (n_136_28), .B (n_141_24), .C1 (n_145_22), .C2 (n_143_21) );
AOI211_X1 g_138_25 (.ZN (n_138_25), .A (n_134_27), .B (n_139_25), .C1 (n_143_23), .C2 (n_145_20) );
AOI211_X1 g_140_24 (.ZN (n_140_24), .A (n_136_26), .B (n_137_26), .C1 (n_141_24), .C2 (n_147_21) );
AOI211_X1 g_142_23 (.ZN (n_142_23), .A (n_138_25), .B (n_136_28), .C1 (n_139_25), .C2 (n_145_22) );
AOI211_X1 g_144_22 (.ZN (n_144_22), .A (n_140_24), .B (n_134_27), .C1 (n_137_26), .C2 (n_143_23) );
AOI211_X1 g_146_23 (.ZN (n_146_23), .A (n_142_23), .B (n_136_26), .C1 (n_136_28), .C2 (n_141_24) );
AOI211_X1 g_144_24 (.ZN (n_144_24), .A (n_144_22), .B (n_138_25), .C1 (n_134_27), .C2 (n_139_25) );
AOI211_X1 g_142_25 (.ZN (n_142_25), .A (n_146_23), .B (n_140_24), .C1 (n_136_26), .C2 (n_137_26) );
AOI211_X1 g_140_26 (.ZN (n_140_26), .A (n_144_24), .B (n_142_23), .C1 (n_138_25), .C2 (n_136_28) );
AOI211_X1 g_138_27 (.ZN (n_138_27), .A (n_142_25), .B (n_144_22), .C1 (n_140_24), .C2 (n_134_27) );
AOI211_X1 g_137_29 (.ZN (n_137_29), .A (n_140_26), .B (n_146_23), .C1 (n_142_23), .C2 (n_136_26) );
AOI211_X1 g_135_28 (.ZN (n_135_28), .A (n_138_27), .B (n_144_24), .C1 (n_144_22), .C2 (n_138_25) );
AOI211_X1 g_137_27 (.ZN (n_137_27), .A (n_137_29), .B (n_142_25), .C1 (n_146_23), .C2 (n_140_24) );
AOI211_X1 g_139_26 (.ZN (n_139_26), .A (n_135_28), .B (n_140_26), .C1 (n_144_24), .C2 (n_142_23) );
AOI211_X1 g_141_25 (.ZN (n_141_25), .A (n_137_27), .B (n_138_27), .C1 (n_142_25), .C2 (n_144_22) );
AOI211_X1 g_143_24 (.ZN (n_143_24), .A (n_139_26), .B (n_137_29), .C1 (n_140_26), .C2 (n_146_23) );
AOI211_X1 g_142_26 (.ZN (n_142_26), .A (n_141_25), .B (n_135_28), .C1 (n_138_27), .C2 (n_144_24) );
AOI211_X1 g_140_27 (.ZN (n_140_27), .A (n_143_24), .B (n_137_27), .C1 (n_137_29), .C2 (n_142_25) );
AOI211_X1 g_138_28 (.ZN (n_138_28), .A (n_142_26), .B (n_139_26), .C1 (n_135_28), .C2 (n_140_26) );
AOI211_X1 g_136_29 (.ZN (n_136_29), .A (n_140_27), .B (n_141_25), .C1 (n_137_27), .C2 (n_138_27) );
AOI211_X1 g_134_28 (.ZN (n_134_28), .A (n_138_28), .B (n_143_24), .C1 (n_139_26), .C2 (n_137_29) );
AOI211_X1 g_132_29 (.ZN (n_132_29), .A (n_136_29), .B (n_142_26), .C1 (n_141_25), .C2 (n_135_28) );
AOI211_X1 g_130_30 (.ZN (n_130_30), .A (n_134_28), .B (n_140_27), .C1 (n_143_24), .C2 (n_137_27) );
AOI211_X1 g_128_31 (.ZN (n_128_31), .A (n_132_29), .B (n_138_28), .C1 (n_142_26), .C2 (n_139_26) );
AOI211_X1 g_126_32 (.ZN (n_126_32), .A (n_130_30), .B (n_136_29), .C1 (n_140_27), .C2 (n_141_25) );
AOI211_X1 g_124_33 (.ZN (n_124_33), .A (n_128_31), .B (n_134_28), .C1 (n_138_28), .C2 (n_143_24) );
AOI211_X1 g_123_31 (.ZN (n_123_31), .A (n_126_32), .B (n_132_29), .C1 (n_136_29), .C2 (n_142_26) );
AOI211_X1 g_121_32 (.ZN (n_121_32), .A (n_124_33), .B (n_130_30), .C1 (n_134_28), .C2 (n_140_27) );
AOI211_X1 g_119_33 (.ZN (n_119_33), .A (n_123_31), .B (n_128_31), .C1 (n_132_29), .C2 (n_138_28) );
AOI211_X1 g_117_34 (.ZN (n_117_34), .A (n_121_32), .B (n_126_32), .C1 (n_130_30), .C2 (n_136_29) );
AOI211_X1 g_115_35 (.ZN (n_115_35), .A (n_119_33), .B (n_124_33), .C1 (n_128_31), .C2 (n_134_28) );
AOI211_X1 g_113_36 (.ZN (n_113_36), .A (n_117_34), .B (n_123_31), .C1 (n_126_32), .C2 (n_132_29) );
AOI211_X1 g_111_37 (.ZN (n_111_37), .A (n_115_35), .B (n_121_32), .C1 (n_124_33), .C2 (n_130_30) );
AOI211_X1 g_109_38 (.ZN (n_109_38), .A (n_113_36), .B (n_119_33), .C1 (n_123_31), .C2 (n_128_31) );
AOI211_X1 g_107_39 (.ZN (n_107_39), .A (n_111_37), .B (n_117_34), .C1 (n_121_32), .C2 (n_126_32) );
AOI211_X1 g_106_37 (.ZN (n_106_37), .A (n_109_38), .B (n_115_35), .C1 (n_119_33), .C2 (n_124_33) );
AOI211_X1 g_104_38 (.ZN (n_104_38), .A (n_107_39), .B (n_113_36), .C1 (n_117_34), .C2 (n_123_31) );
AOI211_X1 g_102_39 (.ZN (n_102_39), .A (n_106_37), .B (n_111_37), .C1 (n_115_35), .C2 (n_121_32) );
AOI211_X1 g_100_40 (.ZN (n_100_40), .A (n_104_38), .B (n_109_38), .C1 (n_113_36), .C2 (n_119_33) );
AOI211_X1 g_98_41 (.ZN (n_98_41), .A (n_102_39), .B (n_107_39), .C1 (n_111_37), .C2 (n_117_34) );
AOI211_X1 g_96_42 (.ZN (n_96_42), .A (n_100_40), .B (n_106_37), .C1 (n_109_38), .C2 (n_115_35) );
AOI211_X1 g_94_43 (.ZN (n_94_43), .A (n_98_41), .B (n_104_38), .C1 (n_107_39), .C2 (n_113_36) );
AOI211_X1 g_92_44 (.ZN (n_92_44), .A (n_96_42), .B (n_102_39), .C1 (n_106_37), .C2 (n_111_37) );
AOI211_X1 g_90_45 (.ZN (n_90_45), .A (n_94_43), .B (n_100_40), .C1 (n_104_38), .C2 (n_109_38) );
AOI211_X1 g_88_46 (.ZN (n_88_46), .A (n_92_44), .B (n_98_41), .C1 (n_102_39), .C2 (n_107_39) );
AOI211_X1 g_86_47 (.ZN (n_86_47), .A (n_90_45), .B (n_96_42), .C1 (n_100_40), .C2 (n_106_37) );
AOI211_X1 g_84_48 (.ZN (n_84_48), .A (n_88_46), .B (n_94_43), .C1 (n_98_41), .C2 (n_104_38) );
AOI211_X1 g_82_49 (.ZN (n_82_49), .A (n_86_47), .B (n_92_44), .C1 (n_96_42), .C2 (n_102_39) );
AOI211_X1 g_80_50 (.ZN (n_80_50), .A (n_84_48), .B (n_90_45), .C1 (n_94_43), .C2 (n_100_40) );
AOI211_X1 g_78_51 (.ZN (n_78_51), .A (n_82_49), .B (n_88_46), .C1 (n_92_44), .C2 (n_98_41) );
AOI211_X1 g_76_52 (.ZN (n_76_52), .A (n_80_50), .B (n_86_47), .C1 (n_90_45), .C2 (n_96_42) );
AOI211_X1 g_74_53 (.ZN (n_74_53), .A (n_78_51), .B (n_84_48), .C1 (n_88_46), .C2 (n_94_43) );
AOI211_X1 g_72_54 (.ZN (n_72_54), .A (n_76_52), .B (n_82_49), .C1 (n_86_47), .C2 (n_92_44) );
AOI211_X1 g_70_55 (.ZN (n_70_55), .A (n_74_53), .B (n_80_50), .C1 (n_84_48), .C2 (n_90_45) );
AOI211_X1 g_68_56 (.ZN (n_68_56), .A (n_72_54), .B (n_78_51), .C1 (n_82_49), .C2 (n_88_46) );
AOI211_X1 g_66_57 (.ZN (n_66_57), .A (n_70_55), .B (n_76_52), .C1 (n_80_50), .C2 (n_86_47) );
AOI211_X1 g_67_55 (.ZN (n_67_55), .A (n_68_56), .B (n_74_53), .C1 (n_78_51), .C2 (n_84_48) );
AOI211_X1 g_65_56 (.ZN (n_65_56), .A (n_66_57), .B (n_72_54), .C1 (n_76_52), .C2 (n_82_49) );
AOI211_X1 g_63_57 (.ZN (n_63_57), .A (n_67_55), .B (n_70_55), .C1 (n_74_53), .C2 (n_80_50) );
AOI211_X1 g_61_58 (.ZN (n_61_58), .A (n_65_56), .B (n_68_56), .C1 (n_72_54), .C2 (n_78_51) );
AOI211_X1 g_59_59 (.ZN (n_59_59), .A (n_63_57), .B (n_66_57), .C1 (n_70_55), .C2 (n_76_52) );
AOI211_X1 g_57_60 (.ZN (n_57_60), .A (n_61_58), .B (n_67_55), .C1 (n_68_56), .C2 (n_74_53) );
AOI211_X1 g_56_62 (.ZN (n_56_62), .A (n_59_59), .B (n_65_56), .C1 (n_66_57), .C2 (n_72_54) );
AOI211_X1 g_58_61 (.ZN (n_58_61), .A (n_57_60), .B (n_63_57), .C1 (n_67_55), .C2 (n_70_55) );
AOI211_X1 g_60_60 (.ZN (n_60_60), .A (n_56_62), .B (n_61_58), .C1 (n_65_56), .C2 (n_68_56) );
AOI211_X1 g_62_59 (.ZN (n_62_59), .A (n_58_61), .B (n_59_59), .C1 (n_63_57), .C2 (n_66_57) );
AOI211_X1 g_64_58 (.ZN (n_64_58), .A (n_60_60), .B (n_57_60), .C1 (n_61_58), .C2 (n_67_55) );
AOI211_X1 g_63_60 (.ZN (n_63_60), .A (n_62_59), .B (n_56_62), .C1 (n_59_59), .C2 (n_65_56) );
AOI211_X1 g_61_59 (.ZN (n_61_59), .A (n_64_58), .B (n_58_61), .C1 (n_57_60), .C2 (n_63_57) );
AOI211_X1 g_63_58 (.ZN (n_63_58), .A (n_63_60), .B (n_60_60), .C1 (n_56_62), .C2 (n_61_58) );
AOI211_X1 g_65_57 (.ZN (n_65_57), .A (n_61_59), .B (n_62_59), .C1 (n_58_61), .C2 (n_59_59) );
AOI211_X1 g_67_56 (.ZN (n_67_56), .A (n_63_58), .B (n_64_58), .C1 (n_60_60), .C2 (n_57_60) );
AOI211_X1 g_69_55 (.ZN (n_69_55), .A (n_65_57), .B (n_63_60), .C1 (n_62_59), .C2 (n_56_62) );
AOI211_X1 g_71_54 (.ZN (n_71_54), .A (n_67_56), .B (n_61_59), .C1 (n_64_58), .C2 (n_58_61) );
AOI211_X1 g_73_53 (.ZN (n_73_53), .A (n_69_55), .B (n_63_58), .C1 (n_63_60), .C2 (n_60_60) );
AOI211_X1 g_75_52 (.ZN (n_75_52), .A (n_71_54), .B (n_65_57), .C1 (n_61_59), .C2 (n_62_59) );
AOI211_X1 g_77_51 (.ZN (n_77_51), .A (n_73_53), .B (n_67_56), .C1 (n_63_58), .C2 (n_64_58) );
AOI211_X1 g_79_50 (.ZN (n_79_50), .A (n_75_52), .B (n_69_55), .C1 (n_65_57), .C2 (n_63_60) );
AOI211_X1 g_81_49 (.ZN (n_81_49), .A (n_77_51), .B (n_71_54), .C1 (n_67_56), .C2 (n_61_59) );
AOI211_X1 g_83_48 (.ZN (n_83_48), .A (n_79_50), .B (n_73_53), .C1 (n_69_55), .C2 (n_63_58) );
AOI211_X1 g_85_47 (.ZN (n_85_47), .A (n_81_49), .B (n_75_52), .C1 (n_71_54), .C2 (n_65_57) );
AOI211_X1 g_87_46 (.ZN (n_87_46), .A (n_83_48), .B (n_77_51), .C1 (n_73_53), .C2 (n_67_56) );
AOI211_X1 g_89_45 (.ZN (n_89_45), .A (n_85_47), .B (n_79_50), .C1 (n_75_52), .C2 (n_69_55) );
AOI211_X1 g_91_44 (.ZN (n_91_44), .A (n_87_46), .B (n_81_49), .C1 (n_77_51), .C2 (n_71_54) );
AOI211_X1 g_93_43 (.ZN (n_93_43), .A (n_89_45), .B (n_83_48), .C1 (n_79_50), .C2 (n_73_53) );
AOI211_X1 g_95_42 (.ZN (n_95_42), .A (n_91_44), .B (n_85_47), .C1 (n_81_49), .C2 (n_75_52) );
AOI211_X1 g_97_41 (.ZN (n_97_41), .A (n_93_43), .B (n_87_46), .C1 (n_83_48), .C2 (n_77_51) );
AOI211_X1 g_99_40 (.ZN (n_99_40), .A (n_95_42), .B (n_89_45), .C1 (n_85_47), .C2 (n_79_50) );
AOI211_X1 g_101_39 (.ZN (n_101_39), .A (n_97_41), .B (n_91_44), .C1 (n_87_46), .C2 (n_81_49) );
AOI211_X1 g_100_41 (.ZN (n_100_41), .A (n_99_40), .B (n_93_43), .C1 (n_89_45), .C2 (n_83_48) );
AOI211_X1 g_102_40 (.ZN (n_102_40), .A (n_101_39), .B (n_95_42), .C1 (n_91_44), .C2 (n_85_47) );
AOI211_X1 g_104_39 (.ZN (n_104_39), .A (n_100_41), .B (n_97_41), .C1 (n_93_43), .C2 (n_87_46) );
AOI211_X1 g_106_38 (.ZN (n_106_38), .A (n_102_40), .B (n_99_40), .C1 (n_95_42), .C2 (n_89_45) );
AOI211_X1 g_105_40 (.ZN (n_105_40), .A (n_104_39), .B (n_101_39), .C1 (n_97_41), .C2 (n_91_44) );
AOI211_X1 g_103_41 (.ZN (n_103_41), .A (n_106_38), .B (n_100_41), .C1 (n_99_40), .C2 (n_93_43) );
AOI211_X1 g_101_42 (.ZN (n_101_42), .A (n_105_40), .B (n_102_40), .C1 (n_101_39), .C2 (n_95_42) );
AOI211_X1 g_99_41 (.ZN (n_99_41), .A (n_103_41), .B (n_104_39), .C1 (n_100_41), .C2 (n_97_41) );
AOI211_X1 g_97_42 (.ZN (n_97_42), .A (n_101_42), .B (n_106_38), .C1 (n_102_40), .C2 (n_99_40) );
AOI211_X1 g_95_43 (.ZN (n_95_43), .A (n_99_41), .B (n_105_40), .C1 (n_104_39), .C2 (n_101_39) );
AOI211_X1 g_93_44 (.ZN (n_93_44), .A (n_97_42), .B (n_103_41), .C1 (n_106_38), .C2 (n_100_41) );
AOI211_X1 g_91_45 (.ZN (n_91_45), .A (n_95_43), .B (n_101_42), .C1 (n_105_40), .C2 (n_102_40) );
AOI211_X1 g_89_46 (.ZN (n_89_46), .A (n_93_44), .B (n_99_41), .C1 (n_103_41), .C2 (n_104_39) );
AOI211_X1 g_87_47 (.ZN (n_87_47), .A (n_91_45), .B (n_97_42), .C1 (n_101_42), .C2 (n_106_38) );
AOI211_X1 g_85_48 (.ZN (n_85_48), .A (n_89_46), .B (n_95_43), .C1 (n_99_41), .C2 (n_105_40) );
AOI211_X1 g_83_49 (.ZN (n_83_49), .A (n_87_47), .B (n_93_44), .C1 (n_97_42), .C2 (n_103_41) );
AOI211_X1 g_81_50 (.ZN (n_81_50), .A (n_85_48), .B (n_91_45), .C1 (n_95_43), .C2 (n_101_42) );
AOI211_X1 g_79_51 (.ZN (n_79_51), .A (n_83_49), .B (n_89_46), .C1 (n_93_44), .C2 (n_99_41) );
AOI211_X1 g_77_52 (.ZN (n_77_52), .A (n_81_50), .B (n_87_47), .C1 (n_91_45), .C2 (n_97_42) );
AOI211_X1 g_75_53 (.ZN (n_75_53), .A (n_79_51), .B (n_85_48), .C1 (n_89_46), .C2 (n_95_43) );
AOI211_X1 g_73_54 (.ZN (n_73_54), .A (n_77_52), .B (n_83_49), .C1 (n_87_47), .C2 (n_93_44) );
AOI211_X1 g_71_55 (.ZN (n_71_55), .A (n_75_53), .B (n_81_50), .C1 (n_85_48), .C2 (n_91_45) );
AOI211_X1 g_69_56 (.ZN (n_69_56), .A (n_73_54), .B (n_79_51), .C1 (n_83_49), .C2 (n_89_46) );
AOI211_X1 g_67_57 (.ZN (n_67_57), .A (n_71_55), .B (n_77_52), .C1 (n_81_50), .C2 (n_87_47) );
AOI211_X1 g_65_58 (.ZN (n_65_58), .A (n_69_56), .B (n_75_53), .C1 (n_79_51), .C2 (n_85_48) );
AOI211_X1 g_63_59 (.ZN (n_63_59), .A (n_67_57), .B (n_73_54), .C1 (n_77_52), .C2 (n_83_49) );
AOI211_X1 g_61_60 (.ZN (n_61_60), .A (n_65_58), .B (n_71_55), .C1 (n_75_53), .C2 (n_81_50) );
AOI211_X1 g_59_61 (.ZN (n_59_61), .A (n_63_59), .B (n_69_56), .C1 (n_73_54), .C2 (n_79_51) );
AOI211_X1 g_57_62 (.ZN (n_57_62), .A (n_61_60), .B (n_67_57), .C1 (n_71_55), .C2 (n_77_52) );
AOI211_X1 g_55_63 (.ZN (n_55_63), .A (n_59_61), .B (n_65_58), .C1 (n_69_56), .C2 (n_75_53) );
AOI211_X1 g_53_64 (.ZN (n_53_64), .A (n_57_62), .B (n_63_59), .C1 (n_67_57), .C2 (n_73_54) );
AOI211_X1 g_51_65 (.ZN (n_51_65), .A (n_55_63), .B (n_61_60), .C1 (n_65_58), .C2 (n_71_55) );
AOI211_X1 g_49_66 (.ZN (n_49_66), .A (n_53_64), .B (n_59_61), .C1 (n_63_59), .C2 (n_69_56) );
AOI211_X1 g_47_67 (.ZN (n_47_67), .A (n_51_65), .B (n_57_62), .C1 (n_61_60), .C2 (n_67_57) );
AOI211_X1 g_45_68 (.ZN (n_45_68), .A (n_49_66), .B (n_55_63), .C1 (n_59_61), .C2 (n_65_58) );
AOI211_X1 g_43_69 (.ZN (n_43_69), .A (n_47_67), .B (n_53_64), .C1 (n_57_62), .C2 (n_63_59) );
AOI211_X1 g_41_70 (.ZN (n_41_70), .A (n_45_68), .B (n_51_65), .C1 (n_55_63), .C2 (n_61_60) );
AOI211_X1 g_39_69 (.ZN (n_39_69), .A (n_43_69), .B (n_49_66), .C1 (n_53_64), .C2 (n_59_61) );
AOI211_X1 g_37_70 (.ZN (n_37_70), .A (n_41_70), .B (n_47_67), .C1 (n_51_65), .C2 (n_57_62) );
AOI211_X1 g_35_71 (.ZN (n_35_71), .A (n_39_69), .B (n_45_68), .C1 (n_49_66), .C2 (n_55_63) );
AOI211_X1 g_33_72 (.ZN (n_33_72), .A (n_37_70), .B (n_43_69), .C1 (n_47_67), .C2 (n_53_64) );
AOI211_X1 g_31_73 (.ZN (n_31_73), .A (n_35_71), .B (n_41_70), .C1 (n_45_68), .C2 (n_51_65) );
AOI211_X1 g_29_74 (.ZN (n_29_74), .A (n_33_72), .B (n_39_69), .C1 (n_43_69), .C2 (n_49_66) );
AOI211_X1 g_27_75 (.ZN (n_27_75), .A (n_31_73), .B (n_37_70), .C1 (n_41_70), .C2 (n_47_67) );
AOI211_X1 g_25_76 (.ZN (n_25_76), .A (n_29_74), .B (n_35_71), .C1 (n_39_69), .C2 (n_45_68) );
AOI211_X1 g_23_77 (.ZN (n_23_77), .A (n_27_75), .B (n_33_72), .C1 (n_37_70), .C2 (n_43_69) );
AOI211_X1 g_21_78 (.ZN (n_21_78), .A (n_25_76), .B (n_31_73), .C1 (n_35_71), .C2 (n_41_70) );
AOI211_X1 g_19_79 (.ZN (n_19_79), .A (n_23_77), .B (n_29_74), .C1 (n_33_72), .C2 (n_39_69) );
AOI211_X1 g_17_80 (.ZN (n_17_80), .A (n_21_78), .B (n_27_75), .C1 (n_31_73), .C2 (n_37_70) );
AOI211_X1 g_15_81 (.ZN (n_15_81), .A (n_19_79), .B (n_25_76), .C1 (n_29_74), .C2 (n_35_71) );
AOI211_X1 g_13_82 (.ZN (n_13_82), .A (n_17_80), .B (n_23_77), .C1 (n_27_75), .C2 (n_33_72) );
AOI211_X1 g_11_83 (.ZN (n_11_83), .A (n_15_81), .B (n_21_78), .C1 (n_25_76), .C2 (n_31_73) );
AOI211_X1 g_9_84 (.ZN (n_9_84), .A (n_13_82), .B (n_19_79), .C1 (n_23_77), .C2 (n_29_74) );
AOI211_X1 g_8_86 (.ZN (n_8_86), .A (n_11_83), .B (n_17_80), .C1 (n_21_78), .C2 (n_27_75) );
AOI211_X1 g_7_84 (.ZN (n_7_84), .A (n_9_84), .B (n_15_81), .C1 (n_19_79), .C2 (n_25_76) );
AOI211_X1 g_5_85 (.ZN (n_5_85), .A (n_8_86), .B (n_13_82), .C1 (n_17_80), .C2 (n_23_77) );
AOI211_X1 g_4_87 (.ZN (n_4_87), .A (n_7_84), .B (n_11_83), .C1 (n_15_81), .C2 (n_21_78) );
AOI211_X1 g_3_89 (.ZN (n_3_89), .A (n_5_85), .B (n_9_84), .C1 (n_13_82), .C2 (n_19_79) );
AOI211_X1 g_5_90 (.ZN (n_5_90), .A (n_4_87), .B (n_8_86), .C1 (n_11_83), .C2 (n_17_80) );
AOI211_X1 g_3_91 (.ZN (n_3_91), .A (n_3_89), .B (n_7_84), .C1 (n_9_84), .C2 (n_15_81) );
AOI211_X1 g_1_92 (.ZN (n_1_92), .A (n_5_90), .B (n_5_85), .C1 (n_8_86), .C2 (n_13_82) );
AOI211_X1 g_2_90 (.ZN (n_2_90), .A (n_3_91), .B (n_4_87), .C1 (n_7_84), .C2 (n_11_83) );
AOI211_X1 g_4_89 (.ZN (n_4_89), .A (n_1_92), .B (n_3_89), .C1 (n_5_85), .C2 (n_9_84) );
AOI211_X1 g_6_88 (.ZN (n_6_88), .A (n_2_90), .B (n_5_90), .C1 (n_4_87), .C2 (n_8_86) );
AOI211_X1 g_7_86 (.ZN (n_7_86), .A (n_4_89), .B (n_3_91), .C1 (n_3_89), .C2 (n_7_84) );
AOI211_X1 g_8_84 (.ZN (n_8_84), .A (n_6_88), .B (n_1_92), .C1 (n_5_90), .C2 (n_5_85) );
AOI211_X1 g_6_85 (.ZN (n_6_85), .A (n_7_86), .B (n_2_90), .C1 (n_3_91), .C2 (n_4_87) );
AOI211_X1 g_4_86 (.ZN (n_4_86), .A (n_8_84), .B (n_4_89), .C1 (n_1_92), .C2 (n_3_89) );
AOI211_X1 g_3_88 (.ZN (n_3_88), .A (n_6_85), .B (n_6_88), .C1 (n_2_90), .C2 (n_5_90) );
AOI211_X1 g_5_87 (.ZN (n_5_87), .A (n_4_86), .B (n_7_86), .C1 (n_4_89), .C2 (n_3_91) );
AOI211_X1 g_6_89 (.ZN (n_6_89), .A (n_3_88), .B (n_8_84), .C1 (n_6_88), .C2 (n_1_92) );
AOI211_X1 g_4_90 (.ZN (n_4_90), .A (n_5_87), .B (n_6_85), .C1 (n_7_86), .C2 (n_2_90) );
AOI211_X1 g_5_88 (.ZN (n_5_88), .A (n_6_89), .B (n_4_86), .C1 (n_8_84), .C2 (n_4_89) );
AOI211_X1 g_6_86 (.ZN (n_6_86), .A (n_4_90), .B (n_3_88), .C1 (n_6_85), .C2 (n_6_88) );
AOI211_X1 g_8_85 (.ZN (n_8_85), .A (n_5_88), .B (n_5_87), .C1 (n_4_86), .C2 (n_7_86) );
AOI211_X1 g_9_83 (.ZN (n_9_83), .A (n_6_86), .B (n_6_89), .C1 (n_3_88), .C2 (n_8_84) );
AOI211_X1 g_11_82 (.ZN (n_11_82), .A (n_8_85), .B (n_4_90), .C1 (n_5_87), .C2 (n_6_85) );
AOI211_X1 g_13_81 (.ZN (n_13_81), .A (n_9_83), .B (n_5_88), .C1 (n_6_89), .C2 (n_4_86) );
AOI211_X1 g_15_80 (.ZN (n_15_80), .A (n_11_82), .B (n_6_86), .C1 (n_4_90), .C2 (n_3_88) );
AOI211_X1 g_17_79 (.ZN (n_17_79), .A (n_13_81), .B (n_8_85), .C1 (n_5_88), .C2 (n_5_87) );
AOI211_X1 g_19_80 (.ZN (n_19_80), .A (n_15_80), .B (n_9_83), .C1 (n_6_86), .C2 (n_6_89) );
AOI211_X1 g_17_81 (.ZN (n_17_81), .A (n_17_79), .B (n_11_82), .C1 (n_8_85), .C2 (n_4_90) );
AOI211_X1 g_18_79 (.ZN (n_18_79), .A (n_19_80), .B (n_13_81), .C1 (n_9_83), .C2 (n_5_88) );
AOI211_X1 g_16_80 (.ZN (n_16_80), .A (n_17_81), .B (n_15_80), .C1 (n_11_82), .C2 (n_6_86) );
AOI211_X1 g_14_81 (.ZN (n_14_81), .A (n_18_79), .B (n_17_79), .C1 (n_13_81), .C2 (n_8_85) );
AOI211_X1 g_12_82 (.ZN (n_12_82), .A (n_16_80), .B (n_19_80), .C1 (n_15_80), .C2 (n_9_83) );
AOI211_X1 g_10_83 (.ZN (n_10_83), .A (n_14_81), .B (n_17_81), .C1 (n_17_79), .C2 (n_11_82) );
AOI211_X1 g_9_85 (.ZN (n_9_85), .A (n_12_82), .B (n_18_79), .C1 (n_19_80), .C2 (n_13_81) );
AOI211_X1 g_11_84 (.ZN (n_11_84), .A (n_10_83), .B (n_16_80), .C1 (n_17_81), .C2 (n_15_80) );
AOI211_X1 g_13_83 (.ZN (n_13_83), .A (n_9_85), .B (n_14_81), .C1 (n_18_79), .C2 (n_17_79) );
AOI211_X1 g_15_82 (.ZN (n_15_82), .A (n_11_84), .B (n_12_82), .C1 (n_16_80), .C2 (n_19_80) );
AOI211_X1 g_14_84 (.ZN (n_14_84), .A (n_13_83), .B (n_10_83), .C1 (n_14_81), .C2 (n_17_81) );
AOI211_X1 g_12_83 (.ZN (n_12_83), .A (n_15_82), .B (n_9_85), .C1 (n_12_82), .C2 (n_18_79) );
AOI211_X1 g_10_84 (.ZN (n_10_84), .A (n_14_84), .B (n_11_84), .C1 (n_10_83), .C2 (n_16_80) );
AOI211_X1 g_12_85 (.ZN (n_12_85), .A (n_12_83), .B (n_13_83), .C1 (n_9_85), .C2 (n_14_81) );
AOI211_X1 g_10_86 (.ZN (n_10_86), .A (n_10_84), .B (n_15_82), .C1 (n_11_84), .C2 (n_12_82) );
AOI211_X1 g_8_87 (.ZN (n_8_87), .A (n_12_85), .B (n_14_84), .C1 (n_13_83), .C2 (n_10_83) );
AOI211_X1 g_7_89 (.ZN (n_7_89), .A (n_10_86), .B (n_12_83), .C1 (n_15_82), .C2 (n_9_85) );
AOI211_X1 g_6_87 (.ZN (n_6_87), .A (n_8_87), .B (n_10_84), .C1 (n_14_84), .C2 (n_11_84) );
AOI211_X1 g_5_89 (.ZN (n_5_89), .A (n_7_89), .B (n_12_85), .C1 (n_12_83), .C2 (n_13_83) );
AOI211_X1 g_7_88 (.ZN (n_7_88), .A (n_6_87), .B (n_10_86), .C1 (n_10_84), .C2 (n_15_82) );
AOI211_X1 g_9_87 (.ZN (n_9_87), .A (n_5_89), .B (n_8_87), .C1 (n_12_85), .C2 (n_14_84) );
AOI211_X1 g_10_85 (.ZN (n_10_85), .A (n_7_88), .B (n_7_89), .C1 (n_10_86), .C2 (n_12_83) );
AOI211_X1 g_12_84 (.ZN (n_12_84), .A (n_9_87), .B (n_6_87), .C1 (n_8_87), .C2 (n_10_84) );
AOI211_X1 g_14_83 (.ZN (n_14_83), .A (n_10_85), .B (n_5_89), .C1 (n_7_89), .C2 (n_12_85) );
AOI211_X1 g_16_82 (.ZN (n_16_82), .A (n_12_84), .B (n_7_88), .C1 (n_6_87), .C2 (n_10_86) );
AOI211_X1 g_18_81 (.ZN (n_18_81), .A (n_14_83), .B (n_9_87), .C1 (n_5_89), .C2 (n_8_87) );
AOI211_X1 g_20_80 (.ZN (n_20_80), .A (n_16_82), .B (n_10_85), .C1 (n_7_88), .C2 (n_7_89) );
AOI211_X1 g_22_79 (.ZN (n_22_79), .A (n_18_81), .B (n_12_84), .C1 (n_9_87), .C2 (n_6_87) );
AOI211_X1 g_24_78 (.ZN (n_24_78), .A (n_20_80), .B (n_14_83), .C1 (n_10_85), .C2 (n_5_89) );
AOI211_X1 g_26_77 (.ZN (n_26_77), .A (n_22_79), .B (n_16_82), .C1 (n_12_84), .C2 (n_7_88) );
AOI211_X1 g_28_76 (.ZN (n_28_76), .A (n_24_78), .B (n_18_81), .C1 (n_14_83), .C2 (n_9_87) );
AOI211_X1 g_30_75 (.ZN (n_30_75), .A (n_26_77), .B (n_20_80), .C1 (n_16_82), .C2 (n_10_85) );
AOI211_X1 g_32_74 (.ZN (n_32_74), .A (n_28_76), .B (n_22_79), .C1 (n_18_81), .C2 (n_12_84) );
AOI211_X1 g_34_73 (.ZN (n_34_73), .A (n_30_75), .B (n_24_78), .C1 (n_20_80), .C2 (n_14_83) );
AOI211_X1 g_36_72 (.ZN (n_36_72), .A (n_32_74), .B (n_26_77), .C1 (n_22_79), .C2 (n_16_82) );
AOI211_X1 g_38_71 (.ZN (n_38_71), .A (n_34_73), .B (n_28_76), .C1 (n_24_78), .C2 (n_18_81) );
AOI211_X1 g_40_70 (.ZN (n_40_70), .A (n_36_72), .B (n_30_75), .C1 (n_26_77), .C2 (n_20_80) );
AOI211_X1 g_42_69 (.ZN (n_42_69), .A (n_38_71), .B (n_32_74), .C1 (n_28_76), .C2 (n_22_79) );
AOI211_X1 g_44_68 (.ZN (n_44_68), .A (n_40_70), .B (n_34_73), .C1 (n_30_75), .C2 (n_24_78) );
AOI211_X1 g_46_67 (.ZN (n_46_67), .A (n_42_69), .B (n_36_72), .C1 (n_32_74), .C2 (n_26_77) );
AOI211_X1 g_48_66 (.ZN (n_48_66), .A (n_44_68), .B (n_38_71), .C1 (n_34_73), .C2 (n_28_76) );
AOI211_X1 g_50_65 (.ZN (n_50_65), .A (n_46_67), .B (n_40_70), .C1 (n_36_72), .C2 (n_30_75) );
AOI211_X1 g_52_64 (.ZN (n_52_64), .A (n_48_66), .B (n_42_69), .C1 (n_38_71), .C2 (n_32_74) );
AOI211_X1 g_54_63 (.ZN (n_54_63), .A (n_50_65), .B (n_44_68), .C1 (n_40_70), .C2 (n_34_73) );
AOI211_X1 g_53_65 (.ZN (n_53_65), .A (n_52_64), .B (n_46_67), .C1 (n_42_69), .C2 (n_36_72) );
AOI211_X1 g_51_64 (.ZN (n_51_64), .A (n_54_63), .B (n_48_66), .C1 (n_44_68), .C2 (n_38_71) );
AOI211_X1 g_53_63 (.ZN (n_53_63), .A (n_53_65), .B (n_50_65), .C1 (n_46_67), .C2 (n_40_70) );
AOI211_X1 g_55_62 (.ZN (n_55_62), .A (n_51_64), .B (n_52_64), .C1 (n_48_66), .C2 (n_42_69) );
AOI211_X1 g_57_61 (.ZN (n_57_61), .A (n_53_63), .B (n_54_63), .C1 (n_50_65), .C2 (n_44_68) );
AOI211_X1 g_59_60 (.ZN (n_59_60), .A (n_55_62), .B (n_53_65), .C1 (n_52_64), .C2 (n_46_67) );
AOI211_X1 g_61_61 (.ZN (n_61_61), .A (n_57_61), .B (n_51_64), .C1 (n_54_63), .C2 (n_48_66) );
AOI211_X1 g_59_62 (.ZN (n_59_62), .A (n_59_60), .B (n_53_63), .C1 (n_53_65), .C2 (n_50_65) );
AOI211_X1 g_57_63 (.ZN (n_57_63), .A (n_61_61), .B (n_55_62), .C1 (n_51_64), .C2 (n_52_64) );
AOI211_X1 g_55_64 (.ZN (n_55_64), .A (n_59_62), .B (n_57_61), .C1 (n_53_63), .C2 (n_54_63) );
AOI211_X1 g_54_66 (.ZN (n_54_66), .A (n_57_63), .B (n_59_60), .C1 (n_55_62), .C2 (n_53_65) );
AOI211_X1 g_52_65 (.ZN (n_52_65), .A (n_55_64), .B (n_61_61), .C1 (n_57_61), .C2 (n_51_64) );
AOI211_X1 g_54_64 (.ZN (n_54_64), .A (n_54_66), .B (n_59_62), .C1 (n_59_60), .C2 (n_53_63) );
AOI211_X1 g_56_63 (.ZN (n_56_63), .A (n_52_65), .B (n_57_63), .C1 (n_61_61), .C2 (n_55_62) );
AOI211_X1 g_58_62 (.ZN (n_58_62), .A (n_54_64), .B (n_55_64), .C1 (n_59_62), .C2 (n_57_61) );
AOI211_X1 g_60_61 (.ZN (n_60_61), .A (n_56_63), .B (n_54_66), .C1 (n_57_63), .C2 (n_59_60) );
AOI211_X1 g_62_60 (.ZN (n_62_60), .A (n_58_62), .B (n_52_65), .C1 (n_55_64), .C2 (n_61_61) );
AOI211_X1 g_64_59 (.ZN (n_64_59), .A (n_60_61), .B (n_54_64), .C1 (n_54_66), .C2 (n_59_62) );
AOI211_X1 g_66_58 (.ZN (n_66_58), .A (n_62_60), .B (n_56_63), .C1 (n_52_65), .C2 (n_57_63) );
AOI211_X1 g_68_57 (.ZN (n_68_57), .A (n_64_59), .B (n_58_62), .C1 (n_54_64), .C2 (n_55_64) );
AOI211_X1 g_70_56 (.ZN (n_70_56), .A (n_66_58), .B (n_60_61), .C1 (n_56_63), .C2 (n_54_66) );
AOI211_X1 g_72_55 (.ZN (n_72_55), .A (n_68_57), .B (n_62_60), .C1 (n_58_62), .C2 (n_52_65) );
AOI211_X1 g_74_54 (.ZN (n_74_54), .A (n_70_56), .B (n_64_59), .C1 (n_60_61), .C2 (n_54_64) );
AOI211_X1 g_76_53 (.ZN (n_76_53), .A (n_72_55), .B (n_66_58), .C1 (n_62_60), .C2 (n_56_63) );
AOI211_X1 g_78_52 (.ZN (n_78_52), .A (n_74_54), .B (n_68_57), .C1 (n_64_59), .C2 (n_58_62) );
AOI211_X1 g_80_51 (.ZN (n_80_51), .A (n_76_53), .B (n_70_56), .C1 (n_66_58), .C2 (n_60_61) );
AOI211_X1 g_82_50 (.ZN (n_82_50), .A (n_78_52), .B (n_72_55), .C1 (n_68_57), .C2 (n_62_60) );
AOI211_X1 g_84_49 (.ZN (n_84_49), .A (n_80_51), .B (n_74_54), .C1 (n_70_56), .C2 (n_64_59) );
AOI211_X1 g_86_48 (.ZN (n_86_48), .A (n_82_50), .B (n_76_53), .C1 (n_72_55), .C2 (n_66_58) );
AOI211_X1 g_88_47 (.ZN (n_88_47), .A (n_84_49), .B (n_78_52), .C1 (n_74_54), .C2 (n_68_57) );
AOI211_X1 g_90_46 (.ZN (n_90_46), .A (n_86_48), .B (n_80_51), .C1 (n_76_53), .C2 (n_70_56) );
AOI211_X1 g_92_45 (.ZN (n_92_45), .A (n_88_47), .B (n_82_50), .C1 (n_78_52), .C2 (n_72_55) );
AOI211_X1 g_94_44 (.ZN (n_94_44), .A (n_90_46), .B (n_84_49), .C1 (n_80_51), .C2 (n_74_54) );
AOI211_X1 g_96_43 (.ZN (n_96_43), .A (n_92_45), .B (n_86_48), .C1 (n_82_50), .C2 (n_76_53) );
AOI211_X1 g_98_42 (.ZN (n_98_42), .A (n_94_44), .B (n_88_47), .C1 (n_84_49), .C2 (n_78_52) );
AOI211_X1 g_97_44 (.ZN (n_97_44), .A (n_96_43), .B (n_90_46), .C1 (n_86_48), .C2 (n_80_51) );
AOI211_X1 g_99_43 (.ZN (n_99_43), .A (n_98_42), .B (n_92_45), .C1 (n_88_47), .C2 (n_82_50) );
AOI211_X1 g_98_45 (.ZN (n_98_45), .A (n_97_44), .B (n_94_44), .C1 (n_90_46), .C2 (n_84_49) );
AOI211_X1 g_97_43 (.ZN (n_97_43), .A (n_99_43), .B (n_96_43), .C1 (n_92_45), .C2 (n_86_48) );
AOI211_X1 g_99_42 (.ZN (n_99_42), .A (n_98_45), .B (n_98_42), .C1 (n_94_44), .C2 (n_88_47) );
AOI211_X1 g_101_41 (.ZN (n_101_41), .A (n_97_43), .B (n_97_44), .C1 (n_96_43), .C2 (n_90_46) );
AOI211_X1 g_103_40 (.ZN (n_103_40), .A (n_99_42), .B (n_99_43), .C1 (n_98_42), .C2 (n_92_45) );
AOI211_X1 g_105_39 (.ZN (n_105_39), .A (n_101_41), .B (n_98_45), .C1 (n_97_44), .C2 (n_94_44) );
AOI211_X1 g_107_38 (.ZN (n_107_38), .A (n_103_40), .B (n_97_43), .C1 (n_99_43), .C2 (n_96_43) );
AOI211_X1 g_106_40 (.ZN (n_106_40), .A (n_105_39), .B (n_99_42), .C1 (n_98_45), .C2 (n_98_42) );
AOI211_X1 g_108_39 (.ZN (n_108_39), .A (n_107_38), .B (n_101_41), .C1 (n_97_43), .C2 (n_97_44) );
AOI211_X1 g_107_41 (.ZN (n_107_41), .A (n_106_40), .B (n_103_40), .C1 (n_99_42), .C2 (n_99_43) );
AOI211_X1 g_106_39 (.ZN (n_106_39), .A (n_108_39), .B (n_105_39), .C1 (n_101_41), .C2 (n_98_45) );
AOI211_X1 g_108_38 (.ZN (n_108_38), .A (n_107_41), .B (n_107_38), .C1 (n_103_40), .C2 (n_97_43) );
AOI211_X1 g_110_37 (.ZN (n_110_37), .A (n_106_39), .B (n_106_40), .C1 (n_105_39), .C2 (n_99_42) );
AOI211_X1 g_112_36 (.ZN (n_112_36), .A (n_108_38), .B (n_108_39), .C1 (n_107_38), .C2 (n_101_41) );
AOI211_X1 g_114_35 (.ZN (n_114_35), .A (n_110_37), .B (n_107_41), .C1 (n_106_40), .C2 (n_103_40) );
AOI211_X1 g_116_34 (.ZN (n_116_34), .A (n_112_36), .B (n_106_39), .C1 (n_108_39), .C2 (n_105_39) );
AOI211_X1 g_115_36 (.ZN (n_115_36), .A (n_114_35), .B (n_108_38), .C1 (n_107_41), .C2 (n_107_38) );
AOI211_X1 g_117_35 (.ZN (n_117_35), .A (n_116_34), .B (n_110_37), .C1 (n_106_39), .C2 (n_106_40) );
AOI211_X1 g_116_37 (.ZN (n_116_37), .A (n_115_36), .B (n_112_36), .C1 (n_108_38), .C2 (n_108_39) );
AOI211_X1 g_114_36 (.ZN (n_114_36), .A (n_117_35), .B (n_114_35), .C1 (n_110_37), .C2 (n_107_41) );
AOI211_X1 g_112_37 (.ZN (n_112_37), .A (n_116_37), .B (n_116_34), .C1 (n_112_36), .C2 (n_106_39) );
AOI211_X1 g_114_38 (.ZN (n_114_38), .A (n_114_36), .B (n_115_36), .C1 (n_114_35), .C2 (n_108_38) );
AOI211_X1 g_112_39 (.ZN (n_112_39), .A (n_112_37), .B (n_117_35), .C1 (n_116_34), .C2 (n_110_37) );
AOI211_X1 g_113_37 (.ZN (n_113_37), .A (n_114_38), .B (n_116_37), .C1 (n_115_36), .C2 (n_112_36) );
AOI211_X1 g_111_38 (.ZN (n_111_38), .A (n_112_39), .B (n_114_36), .C1 (n_117_35), .C2 (n_114_35) );
AOI211_X1 g_109_39 (.ZN (n_109_39), .A (n_113_37), .B (n_112_37), .C1 (n_116_37), .C2 (n_116_34) );
AOI211_X1 g_107_40 (.ZN (n_107_40), .A (n_111_38), .B (n_114_38), .C1 (n_114_36), .C2 (n_115_36) );
AOI211_X1 g_105_41 (.ZN (n_105_41), .A (n_109_39), .B (n_112_39), .C1 (n_112_37), .C2 (n_117_35) );
AOI211_X1 g_103_42 (.ZN (n_103_42), .A (n_107_40), .B (n_113_37), .C1 (n_114_38), .C2 (n_116_37) );
AOI211_X1 g_104_40 (.ZN (n_104_40), .A (n_105_41), .B (n_111_38), .C1 (n_112_39), .C2 (n_114_36) );
AOI211_X1 g_102_41 (.ZN (n_102_41), .A (n_103_42), .B (n_109_39), .C1 (n_113_37), .C2 (n_112_37) );
AOI211_X1 g_100_42 (.ZN (n_100_42), .A (n_104_40), .B (n_107_40), .C1 (n_111_38), .C2 (n_114_38) );
AOI211_X1 g_98_43 (.ZN (n_98_43), .A (n_102_41), .B (n_105_41), .C1 (n_109_39), .C2 (n_112_39) );
AOI211_X1 g_96_44 (.ZN (n_96_44), .A (n_100_42), .B (n_103_42), .C1 (n_107_40), .C2 (n_113_37) );
AOI211_X1 g_94_45 (.ZN (n_94_45), .A (n_98_43), .B (n_104_40), .C1 (n_105_41), .C2 (n_111_38) );
AOI211_X1 g_92_46 (.ZN (n_92_46), .A (n_96_44), .B (n_102_41), .C1 (n_103_42), .C2 (n_109_39) );
AOI211_X1 g_90_47 (.ZN (n_90_47), .A (n_94_45), .B (n_100_42), .C1 (n_104_40), .C2 (n_107_40) );
AOI211_X1 g_88_48 (.ZN (n_88_48), .A (n_92_46), .B (n_98_43), .C1 (n_102_41), .C2 (n_105_41) );
AOI211_X1 g_86_49 (.ZN (n_86_49), .A (n_90_47), .B (n_96_44), .C1 (n_100_42), .C2 (n_103_42) );
AOI211_X1 g_84_50 (.ZN (n_84_50), .A (n_88_48), .B (n_94_45), .C1 (n_98_43), .C2 (n_104_40) );
AOI211_X1 g_82_51 (.ZN (n_82_51), .A (n_86_49), .B (n_92_46), .C1 (n_96_44), .C2 (n_102_41) );
AOI211_X1 g_80_52 (.ZN (n_80_52), .A (n_84_50), .B (n_90_47), .C1 (n_94_45), .C2 (n_100_42) );
AOI211_X1 g_78_53 (.ZN (n_78_53), .A (n_82_51), .B (n_88_48), .C1 (n_92_46), .C2 (n_98_43) );
AOI211_X1 g_76_54 (.ZN (n_76_54), .A (n_80_52), .B (n_86_49), .C1 (n_90_47), .C2 (n_96_44) );
AOI211_X1 g_74_55 (.ZN (n_74_55), .A (n_78_53), .B (n_84_50), .C1 (n_88_48), .C2 (n_94_45) );
AOI211_X1 g_72_56 (.ZN (n_72_56), .A (n_76_54), .B (n_82_51), .C1 (n_86_49), .C2 (n_92_46) );
AOI211_X1 g_70_57 (.ZN (n_70_57), .A (n_74_55), .B (n_80_52), .C1 (n_84_50), .C2 (n_90_47) );
AOI211_X1 g_68_58 (.ZN (n_68_58), .A (n_72_56), .B (n_78_53), .C1 (n_82_51), .C2 (n_88_48) );
AOI211_X1 g_66_59 (.ZN (n_66_59), .A (n_70_57), .B (n_76_54), .C1 (n_80_52), .C2 (n_86_49) );
AOI211_X1 g_64_60 (.ZN (n_64_60), .A (n_68_58), .B (n_74_55), .C1 (n_78_53), .C2 (n_84_50) );
AOI211_X1 g_62_61 (.ZN (n_62_61), .A (n_66_59), .B (n_72_56), .C1 (n_76_54), .C2 (n_82_51) );
AOI211_X1 g_60_62 (.ZN (n_60_62), .A (n_64_60), .B (n_70_57), .C1 (n_74_55), .C2 (n_80_52) );
AOI211_X1 g_58_63 (.ZN (n_58_63), .A (n_62_61), .B (n_68_58), .C1 (n_72_56), .C2 (n_78_53) );
AOI211_X1 g_56_64 (.ZN (n_56_64), .A (n_60_62), .B (n_66_59), .C1 (n_70_57), .C2 (n_76_54) );
AOI211_X1 g_54_65 (.ZN (n_54_65), .A (n_58_63), .B (n_64_60), .C1 (n_68_58), .C2 (n_74_55) );
AOI211_X1 g_52_66 (.ZN (n_52_66), .A (n_56_64), .B (n_62_61), .C1 (n_66_59), .C2 (n_72_56) );
AOI211_X1 g_50_67 (.ZN (n_50_67), .A (n_54_65), .B (n_60_62), .C1 (n_64_60), .C2 (n_70_57) );
AOI211_X1 g_49_65 (.ZN (n_49_65), .A (n_52_66), .B (n_58_63), .C1 (n_62_61), .C2 (n_68_58) );
AOI211_X1 g_47_66 (.ZN (n_47_66), .A (n_50_67), .B (n_56_64), .C1 (n_60_62), .C2 (n_66_59) );
AOI211_X1 g_45_67 (.ZN (n_45_67), .A (n_49_65), .B (n_54_65), .C1 (n_58_63), .C2 (n_64_60) );
AOI211_X1 g_43_68 (.ZN (n_43_68), .A (n_47_66), .B (n_52_66), .C1 (n_56_64), .C2 (n_62_61) );
AOI211_X1 g_41_69 (.ZN (n_41_69), .A (n_45_67), .B (n_50_67), .C1 (n_54_65), .C2 (n_60_62) );
AOI211_X1 g_39_70 (.ZN (n_39_70), .A (n_43_68), .B (n_49_65), .C1 (n_52_66), .C2 (n_58_63) );
AOI211_X1 g_37_71 (.ZN (n_37_71), .A (n_41_69), .B (n_47_66), .C1 (n_50_67), .C2 (n_56_64) );
AOI211_X1 g_35_72 (.ZN (n_35_72), .A (n_39_70), .B (n_45_67), .C1 (n_49_65), .C2 (n_54_65) );
AOI211_X1 g_33_73 (.ZN (n_33_73), .A (n_37_71), .B (n_43_68), .C1 (n_47_66), .C2 (n_52_66) );
AOI211_X1 g_31_74 (.ZN (n_31_74), .A (n_35_72), .B (n_41_69), .C1 (n_45_67), .C2 (n_50_67) );
AOI211_X1 g_29_75 (.ZN (n_29_75), .A (n_33_73), .B (n_39_70), .C1 (n_43_68), .C2 (n_49_65) );
AOI211_X1 g_27_76 (.ZN (n_27_76), .A (n_31_74), .B (n_37_71), .C1 (n_41_69), .C2 (n_47_66) );
AOI211_X1 g_25_77 (.ZN (n_25_77), .A (n_29_75), .B (n_35_72), .C1 (n_39_70), .C2 (n_45_67) );
AOI211_X1 g_23_78 (.ZN (n_23_78), .A (n_27_76), .B (n_33_73), .C1 (n_37_71), .C2 (n_43_68) );
AOI211_X1 g_22_80 (.ZN (n_22_80), .A (n_25_77), .B (n_31_74), .C1 (n_35_72), .C2 (n_41_69) );
AOI211_X1 g_20_79 (.ZN (n_20_79), .A (n_23_78), .B (n_29_75), .C1 (n_33_73), .C2 (n_39_70) );
AOI211_X1 g_22_78 (.ZN (n_22_78), .A (n_22_80), .B (n_27_76), .C1 (n_31_74), .C2 (n_37_71) );
AOI211_X1 g_24_77 (.ZN (n_24_77), .A (n_20_79), .B (n_25_77), .C1 (n_29_75), .C2 (n_35_72) );
AOI211_X1 g_23_79 (.ZN (n_23_79), .A (n_22_78), .B (n_23_78), .C1 (n_27_76), .C2 (n_33_73) );
AOI211_X1 g_25_78 (.ZN (n_25_78), .A (n_24_77), .B (n_22_80), .C1 (n_25_77), .C2 (n_31_74) );
AOI211_X1 g_27_77 (.ZN (n_27_77), .A (n_23_79), .B (n_20_79), .C1 (n_23_78), .C2 (n_29_75) );
AOI211_X1 g_29_76 (.ZN (n_29_76), .A (n_25_78), .B (n_22_78), .C1 (n_22_80), .C2 (n_27_76) );
AOI211_X1 g_31_75 (.ZN (n_31_75), .A (n_27_77), .B (n_24_77), .C1 (n_20_79), .C2 (n_25_77) );
AOI211_X1 g_33_74 (.ZN (n_33_74), .A (n_29_76), .B (n_23_79), .C1 (n_22_78), .C2 (n_23_78) );
AOI211_X1 g_35_73 (.ZN (n_35_73), .A (n_31_75), .B (n_25_78), .C1 (n_24_77), .C2 (n_22_80) );
AOI211_X1 g_37_72 (.ZN (n_37_72), .A (n_33_74), .B (n_27_77), .C1 (n_23_79), .C2 (n_20_79) );
AOI211_X1 g_39_71 (.ZN (n_39_71), .A (n_35_73), .B (n_29_76), .C1 (n_25_78), .C2 (n_22_78) );
AOI211_X1 g_38_73 (.ZN (n_38_73), .A (n_37_72), .B (n_31_75), .C1 (n_27_77), .C2 (n_24_77) );
AOI211_X1 g_40_72 (.ZN (n_40_72), .A (n_39_71), .B (n_33_74), .C1 (n_29_76), .C2 (n_23_79) );
AOI211_X1 g_42_71 (.ZN (n_42_71), .A (n_38_73), .B (n_35_73), .C1 (n_31_75), .C2 (n_25_78) );
AOI211_X1 g_44_70 (.ZN (n_44_70), .A (n_40_72), .B (n_37_72), .C1 (n_33_74), .C2 (n_27_77) );
AOI211_X1 g_46_69 (.ZN (n_46_69), .A (n_42_71), .B (n_39_71), .C1 (n_35_73), .C2 (n_29_76) );
AOI211_X1 g_48_68 (.ZN (n_48_68), .A (n_44_70), .B (n_38_73), .C1 (n_37_72), .C2 (n_31_75) );
AOI211_X1 g_47_70 (.ZN (n_47_70), .A (n_46_69), .B (n_40_72), .C1 (n_39_71), .C2 (n_33_74) );
AOI211_X1 g_46_68 (.ZN (n_46_68), .A (n_48_68), .B (n_42_71), .C1 (n_38_73), .C2 (n_35_73) );
AOI211_X1 g_48_67 (.ZN (n_48_67), .A (n_47_70), .B (n_44_70), .C1 (n_40_72), .C2 (n_37_72) );
AOI211_X1 g_50_66 (.ZN (n_50_66), .A (n_46_68), .B (n_46_69), .C1 (n_42_71), .C2 (n_39_71) );
AOI211_X1 g_52_67 (.ZN (n_52_67), .A (n_48_67), .B (n_48_68), .C1 (n_44_70), .C2 (n_38_73) );
AOI211_X1 g_50_68 (.ZN (n_50_68), .A (n_50_66), .B (n_47_70), .C1 (n_46_69), .C2 (n_40_72) );
AOI211_X1 g_51_66 (.ZN (n_51_66), .A (n_52_67), .B (n_46_68), .C1 (n_48_68), .C2 (n_42_71) );
AOI211_X1 g_49_67 (.ZN (n_49_67), .A (n_50_68), .B (n_48_67), .C1 (n_47_70), .C2 (n_44_70) );
AOI211_X1 g_47_68 (.ZN (n_47_68), .A (n_51_66), .B (n_50_66), .C1 (n_46_68), .C2 (n_46_69) );
AOI211_X1 g_45_69 (.ZN (n_45_69), .A (n_49_67), .B (n_52_67), .C1 (n_48_67), .C2 (n_48_68) );
AOI211_X1 g_43_70 (.ZN (n_43_70), .A (n_47_68), .B (n_50_68), .C1 (n_50_66), .C2 (n_47_70) );
AOI211_X1 g_41_71 (.ZN (n_41_71), .A (n_45_69), .B (n_51_66), .C1 (n_52_67), .C2 (n_46_68) );
AOI211_X1 g_39_72 (.ZN (n_39_72), .A (n_43_70), .B (n_49_67), .C1 (n_50_68), .C2 (n_48_67) );
AOI211_X1 g_37_73 (.ZN (n_37_73), .A (n_41_71), .B (n_47_68), .C1 (n_51_66), .C2 (n_50_66) );
AOI211_X1 g_35_74 (.ZN (n_35_74), .A (n_39_72), .B (n_45_69), .C1 (n_49_67), .C2 (n_52_67) );
AOI211_X1 g_33_75 (.ZN (n_33_75), .A (n_37_73), .B (n_43_70), .C1 (n_47_68), .C2 (n_50_68) );
AOI211_X1 g_31_76 (.ZN (n_31_76), .A (n_35_74), .B (n_41_71), .C1 (n_45_69), .C2 (n_51_66) );
AOI211_X1 g_29_77 (.ZN (n_29_77), .A (n_33_75), .B (n_39_72), .C1 (n_43_70), .C2 (n_49_67) );
AOI211_X1 g_27_78 (.ZN (n_27_78), .A (n_31_76), .B (n_37_73), .C1 (n_41_71), .C2 (n_47_68) );
AOI211_X1 g_25_79 (.ZN (n_25_79), .A (n_29_77), .B (n_35_74), .C1 (n_39_72), .C2 (n_45_69) );
AOI211_X1 g_23_80 (.ZN (n_23_80), .A (n_27_78), .B (n_33_75), .C1 (n_37_73), .C2 (n_43_70) );
AOI211_X1 g_21_81 (.ZN (n_21_81), .A (n_25_79), .B (n_31_76), .C1 (n_35_74), .C2 (n_41_71) );
AOI211_X1 g_19_82 (.ZN (n_19_82), .A (n_23_80), .B (n_29_77), .C1 (n_33_75), .C2 (n_39_72) );
AOI211_X1 g_18_80 (.ZN (n_18_80), .A (n_21_81), .B (n_27_78), .C1 (n_31_76), .C2 (n_37_73) );
AOI211_X1 g_16_81 (.ZN (n_16_81), .A (n_19_82), .B (n_25_79), .C1 (n_29_77), .C2 (n_35_74) );
AOI211_X1 g_14_82 (.ZN (n_14_82), .A (n_18_80), .B (n_23_80), .C1 (n_27_78), .C2 (n_33_75) );
AOI211_X1 g_16_83 (.ZN (n_16_83), .A (n_16_81), .B (n_21_81), .C1 (n_25_79), .C2 (n_31_76) );
AOI211_X1 g_18_82 (.ZN (n_18_82), .A (n_14_82), .B (n_19_82), .C1 (n_23_80), .C2 (n_29_77) );
AOI211_X1 g_20_81 (.ZN (n_20_81), .A (n_16_83), .B (n_18_80), .C1 (n_21_81), .C2 (n_27_78) );
AOI211_X1 g_19_83 (.ZN (n_19_83), .A (n_18_82), .B (n_16_81), .C1 (n_19_82), .C2 (n_25_79) );
AOI211_X1 g_17_82 (.ZN (n_17_82), .A (n_20_81), .B (n_14_82), .C1 (n_18_80), .C2 (n_23_80) );
AOI211_X1 g_19_81 (.ZN (n_19_81), .A (n_19_83), .B (n_16_83), .C1 (n_16_81), .C2 (n_21_81) );
AOI211_X1 g_21_80 (.ZN (n_21_80), .A (n_17_82), .B (n_18_82), .C1 (n_14_82), .C2 (n_19_82) );
AOI211_X1 g_20_82 (.ZN (n_20_82), .A (n_19_81), .B (n_20_81), .C1 (n_16_83), .C2 (n_18_80) );
AOI211_X1 g_22_81 (.ZN (n_22_81), .A (n_21_80), .B (n_19_83), .C1 (n_18_82), .C2 (n_16_81) );
AOI211_X1 g_24_80 (.ZN (n_24_80), .A (n_20_82), .B (n_17_82), .C1 (n_20_81), .C2 (n_14_82) );
AOI211_X1 g_26_79 (.ZN (n_26_79), .A (n_22_81), .B (n_19_81), .C1 (n_19_83), .C2 (n_16_83) );
AOI211_X1 g_28_78 (.ZN (n_28_78), .A (n_24_80), .B (n_21_80), .C1 (n_17_82), .C2 (n_18_82) );
AOI211_X1 g_30_77 (.ZN (n_30_77), .A (n_26_79), .B (n_20_82), .C1 (n_19_81), .C2 (n_20_81) );
AOI211_X1 g_32_76 (.ZN (n_32_76), .A (n_28_78), .B (n_22_81), .C1 (n_21_80), .C2 (n_19_83) );
AOI211_X1 g_34_75 (.ZN (n_34_75), .A (n_30_77), .B (n_24_80), .C1 (n_20_82), .C2 (n_17_82) );
AOI211_X1 g_36_74 (.ZN (n_36_74), .A (n_32_76), .B (n_26_79), .C1 (n_22_81), .C2 (n_19_81) );
AOI211_X1 g_35_76 (.ZN (n_35_76), .A (n_34_75), .B (n_28_78), .C1 (n_24_80), .C2 (n_21_80) );
AOI211_X1 g_34_74 (.ZN (n_34_74), .A (n_36_74), .B (n_30_77), .C1 (n_26_79), .C2 (n_20_82) );
AOI211_X1 g_36_73 (.ZN (n_36_73), .A (n_35_76), .B (n_32_76), .C1 (n_28_78), .C2 (n_22_81) );
AOI211_X1 g_38_72 (.ZN (n_38_72), .A (n_34_74), .B (n_34_75), .C1 (n_30_77), .C2 (n_24_80) );
AOI211_X1 g_40_71 (.ZN (n_40_71), .A (n_36_73), .B (n_36_74), .C1 (n_32_76), .C2 (n_26_79) );
AOI211_X1 g_42_70 (.ZN (n_42_70), .A (n_38_72), .B (n_35_76), .C1 (n_34_75), .C2 (n_28_78) );
AOI211_X1 g_44_69 (.ZN (n_44_69), .A (n_40_71), .B (n_34_74), .C1 (n_36_74), .C2 (n_30_77) );
AOI211_X1 g_45_71 (.ZN (n_45_71), .A (n_42_70), .B (n_36_73), .C1 (n_35_76), .C2 (n_32_76) );
AOI211_X1 g_43_72 (.ZN (n_43_72), .A (n_44_69), .B (n_38_72), .C1 (n_34_74), .C2 (n_34_75) );
AOI211_X1 g_41_73 (.ZN (n_41_73), .A (n_45_71), .B (n_40_71), .C1 (n_36_73), .C2 (n_36_74) );
AOI211_X1 g_39_74 (.ZN (n_39_74), .A (n_43_72), .B (n_42_70), .C1 (n_38_72), .C2 (n_35_76) );
AOI211_X1 g_37_75 (.ZN (n_37_75), .A (n_41_73), .B (n_44_69), .C1 (n_40_71), .C2 (n_34_74) );
AOI211_X1 g_36_77 (.ZN (n_36_77), .A (n_39_74), .B (n_45_71), .C1 (n_42_70), .C2 (n_36_73) );
AOI211_X1 g_35_75 (.ZN (n_35_75), .A (n_37_75), .B (n_43_72), .C1 (n_44_69), .C2 (n_38_72) );
AOI211_X1 g_37_74 (.ZN (n_37_74), .A (n_36_77), .B (n_41_73), .C1 (n_45_71), .C2 (n_40_71) );
AOI211_X1 g_39_73 (.ZN (n_39_73), .A (n_35_75), .B (n_39_74), .C1 (n_43_72), .C2 (n_42_70) );
AOI211_X1 g_41_72 (.ZN (n_41_72), .A (n_37_74), .B (n_37_75), .C1 (n_41_73), .C2 (n_44_69) );
AOI211_X1 g_43_71 (.ZN (n_43_71), .A (n_39_73), .B (n_36_77), .C1 (n_39_74), .C2 (n_45_71) );
AOI211_X1 g_45_70 (.ZN (n_45_70), .A (n_41_72), .B (n_35_75), .C1 (n_37_75), .C2 (n_43_72) );
AOI211_X1 g_47_69 (.ZN (n_47_69), .A (n_43_71), .B (n_37_74), .C1 (n_36_77), .C2 (n_41_73) );
AOI211_X1 g_49_68 (.ZN (n_49_68), .A (n_45_70), .B (n_39_73), .C1 (n_35_75), .C2 (n_39_74) );
AOI211_X1 g_51_67 (.ZN (n_51_67), .A (n_47_69), .B (n_41_72), .C1 (n_37_74), .C2 (n_37_75) );
AOI211_X1 g_53_66 (.ZN (n_53_66), .A (n_49_68), .B (n_43_71), .C1 (n_39_73), .C2 (n_36_77) );
AOI211_X1 g_55_65 (.ZN (n_55_65), .A (n_51_67), .B (n_45_70), .C1 (n_41_72), .C2 (n_35_75) );
AOI211_X1 g_57_64 (.ZN (n_57_64), .A (n_53_66), .B (n_47_69), .C1 (n_43_71), .C2 (n_37_74) );
AOI211_X1 g_59_63 (.ZN (n_59_63), .A (n_55_65), .B (n_49_68), .C1 (n_45_70), .C2 (n_39_73) );
AOI211_X1 g_61_62 (.ZN (n_61_62), .A (n_57_64), .B (n_51_67), .C1 (n_47_69), .C2 (n_41_72) );
AOI211_X1 g_63_61 (.ZN (n_63_61), .A (n_59_63), .B (n_53_66), .C1 (n_49_68), .C2 (n_43_71) );
AOI211_X1 g_65_60 (.ZN (n_65_60), .A (n_61_62), .B (n_55_65), .C1 (n_51_67), .C2 (n_45_70) );
AOI211_X1 g_67_59 (.ZN (n_67_59), .A (n_63_61), .B (n_57_64), .C1 (n_53_66), .C2 (n_47_69) );
AOI211_X1 g_69_58 (.ZN (n_69_58), .A (n_65_60), .B (n_59_63), .C1 (n_55_65), .C2 (n_49_68) );
AOI211_X1 g_71_57 (.ZN (n_71_57), .A (n_67_59), .B (n_61_62), .C1 (n_57_64), .C2 (n_51_67) );
AOI211_X1 g_73_56 (.ZN (n_73_56), .A (n_69_58), .B (n_63_61), .C1 (n_59_63), .C2 (n_53_66) );
AOI211_X1 g_75_55 (.ZN (n_75_55), .A (n_71_57), .B (n_65_60), .C1 (n_61_62), .C2 (n_55_65) );
AOI211_X1 g_77_54 (.ZN (n_77_54), .A (n_73_56), .B (n_67_59), .C1 (n_63_61), .C2 (n_57_64) );
AOI211_X1 g_79_53 (.ZN (n_79_53), .A (n_75_55), .B (n_69_58), .C1 (n_65_60), .C2 (n_59_63) );
AOI211_X1 g_81_52 (.ZN (n_81_52), .A (n_77_54), .B (n_71_57), .C1 (n_67_59), .C2 (n_61_62) );
AOI211_X1 g_83_51 (.ZN (n_83_51), .A (n_79_53), .B (n_73_56), .C1 (n_69_58), .C2 (n_63_61) );
AOI211_X1 g_85_50 (.ZN (n_85_50), .A (n_81_52), .B (n_75_55), .C1 (n_71_57), .C2 (n_65_60) );
AOI211_X1 g_87_49 (.ZN (n_87_49), .A (n_83_51), .B (n_77_54), .C1 (n_73_56), .C2 (n_67_59) );
AOI211_X1 g_89_48 (.ZN (n_89_48), .A (n_85_50), .B (n_79_53), .C1 (n_75_55), .C2 (n_69_58) );
AOI211_X1 g_91_47 (.ZN (n_91_47), .A (n_87_49), .B (n_81_52), .C1 (n_77_54), .C2 (n_71_57) );
AOI211_X1 g_93_46 (.ZN (n_93_46), .A (n_89_48), .B (n_83_51), .C1 (n_79_53), .C2 (n_73_56) );
AOI211_X1 g_95_45 (.ZN (n_95_45), .A (n_91_47), .B (n_85_50), .C1 (n_81_52), .C2 (n_75_55) );
AOI211_X1 g_94_47 (.ZN (n_94_47), .A (n_93_46), .B (n_87_49), .C1 (n_83_51), .C2 (n_77_54) );
AOI211_X1 g_96_46 (.ZN (n_96_46), .A (n_95_45), .B (n_89_48), .C1 (n_85_50), .C2 (n_79_53) );
AOI211_X1 g_95_44 (.ZN (n_95_44), .A (n_94_47), .B (n_91_47), .C1 (n_87_49), .C2 (n_81_52) );
AOI211_X1 g_93_45 (.ZN (n_93_45), .A (n_96_46), .B (n_93_46), .C1 (n_89_48), .C2 (n_83_51) );
AOI211_X1 g_91_46 (.ZN (n_91_46), .A (n_95_44), .B (n_95_45), .C1 (n_91_47), .C2 (n_85_50) );
AOI211_X1 g_89_47 (.ZN (n_89_47), .A (n_93_45), .B (n_94_47), .C1 (n_93_46), .C2 (n_87_49) );
AOI211_X1 g_87_48 (.ZN (n_87_48), .A (n_91_46), .B (n_96_46), .C1 (n_95_45), .C2 (n_89_48) );
AOI211_X1 g_85_49 (.ZN (n_85_49), .A (n_89_47), .B (n_95_44), .C1 (n_94_47), .C2 (n_91_47) );
AOI211_X1 g_83_50 (.ZN (n_83_50), .A (n_87_48), .B (n_93_45), .C1 (n_96_46), .C2 (n_93_46) );
AOI211_X1 g_81_51 (.ZN (n_81_51), .A (n_85_49), .B (n_91_46), .C1 (n_95_44), .C2 (n_95_45) );
AOI211_X1 g_79_52 (.ZN (n_79_52), .A (n_83_50), .B (n_89_47), .C1 (n_93_45), .C2 (n_94_47) );
AOI211_X1 g_77_53 (.ZN (n_77_53), .A (n_81_51), .B (n_87_48), .C1 (n_91_46), .C2 (n_96_46) );
AOI211_X1 g_75_54 (.ZN (n_75_54), .A (n_79_52), .B (n_85_49), .C1 (n_89_47), .C2 (n_95_44) );
AOI211_X1 g_73_55 (.ZN (n_73_55), .A (n_77_53), .B (n_83_50), .C1 (n_87_48), .C2 (n_93_45) );
AOI211_X1 g_71_56 (.ZN (n_71_56), .A (n_75_54), .B (n_81_51), .C1 (n_85_49), .C2 (n_91_46) );
AOI211_X1 g_69_57 (.ZN (n_69_57), .A (n_73_55), .B (n_79_52), .C1 (n_83_50), .C2 (n_89_47) );
AOI211_X1 g_67_58 (.ZN (n_67_58), .A (n_71_56), .B (n_77_53), .C1 (n_81_51), .C2 (n_87_48) );
AOI211_X1 g_65_59 (.ZN (n_65_59), .A (n_69_57), .B (n_75_54), .C1 (n_79_52), .C2 (n_85_49) );
AOI211_X1 g_64_61 (.ZN (n_64_61), .A (n_67_58), .B (n_73_55), .C1 (n_77_53), .C2 (n_83_50) );
AOI211_X1 g_66_60 (.ZN (n_66_60), .A (n_65_59), .B (n_71_56), .C1 (n_75_54), .C2 (n_81_51) );
AOI211_X1 g_68_59 (.ZN (n_68_59), .A (n_64_61), .B (n_69_57), .C1 (n_73_55), .C2 (n_79_52) );
AOI211_X1 g_70_58 (.ZN (n_70_58), .A (n_66_60), .B (n_67_58), .C1 (n_71_56), .C2 (n_77_53) );
AOI211_X1 g_72_57 (.ZN (n_72_57), .A (n_68_59), .B (n_65_59), .C1 (n_69_57), .C2 (n_75_54) );
AOI211_X1 g_74_56 (.ZN (n_74_56), .A (n_70_58), .B (n_64_61), .C1 (n_67_58), .C2 (n_73_55) );
AOI211_X1 g_76_55 (.ZN (n_76_55), .A (n_72_57), .B (n_66_60), .C1 (n_65_59), .C2 (n_71_56) );
AOI211_X1 g_78_54 (.ZN (n_78_54), .A (n_74_56), .B (n_68_59), .C1 (n_64_61), .C2 (n_69_57) );
AOI211_X1 g_80_53 (.ZN (n_80_53), .A (n_76_55), .B (n_70_58), .C1 (n_66_60), .C2 (n_67_58) );
AOI211_X1 g_82_52 (.ZN (n_82_52), .A (n_78_54), .B (n_72_57), .C1 (n_68_59), .C2 (n_65_59) );
AOI211_X1 g_84_51 (.ZN (n_84_51), .A (n_80_53), .B (n_74_56), .C1 (n_70_58), .C2 (n_64_61) );
AOI211_X1 g_86_50 (.ZN (n_86_50), .A (n_82_52), .B (n_76_55), .C1 (n_72_57), .C2 (n_66_60) );
AOI211_X1 g_88_49 (.ZN (n_88_49), .A (n_84_51), .B (n_78_54), .C1 (n_74_56), .C2 (n_68_59) );
AOI211_X1 g_90_48 (.ZN (n_90_48), .A (n_86_50), .B (n_80_53), .C1 (n_76_55), .C2 (n_70_58) );
AOI211_X1 g_92_47 (.ZN (n_92_47), .A (n_88_49), .B (n_82_52), .C1 (n_78_54), .C2 (n_72_57) );
AOI211_X1 g_94_46 (.ZN (n_94_46), .A (n_90_48), .B (n_84_51), .C1 (n_80_53), .C2 (n_74_56) );
AOI211_X1 g_96_45 (.ZN (n_96_45), .A (n_92_47), .B (n_86_50), .C1 (n_82_52), .C2 (n_76_55) );
AOI211_X1 g_98_44 (.ZN (n_98_44), .A (n_94_46), .B (n_88_49), .C1 (n_84_51), .C2 (n_78_54) );
AOI211_X1 g_100_43 (.ZN (n_100_43), .A (n_96_45), .B (n_90_48), .C1 (n_86_50), .C2 (n_80_53) );
AOI211_X1 g_102_42 (.ZN (n_102_42), .A (n_98_44), .B (n_92_47), .C1 (n_88_49), .C2 (n_82_52) );
AOI211_X1 g_104_41 (.ZN (n_104_41), .A (n_100_43), .B (n_94_46), .C1 (n_90_48), .C2 (n_84_51) );
AOI211_X1 g_103_43 (.ZN (n_103_43), .A (n_102_42), .B (n_96_45), .C1 (n_92_47), .C2 (n_86_50) );
AOI211_X1 g_105_42 (.ZN (n_105_42), .A (n_104_41), .B (n_98_44), .C1 (n_94_46), .C2 (n_88_49) );
AOI211_X1 g_104_44 (.ZN (n_104_44), .A (n_103_43), .B (n_100_43), .C1 (n_96_45), .C2 (n_90_48) );
AOI211_X1 g_102_43 (.ZN (n_102_43), .A (n_105_42), .B (n_102_42), .C1 (n_98_44), .C2 (n_92_47) );
AOI211_X1 g_100_44 (.ZN (n_100_44), .A (n_104_44), .B (n_104_41), .C1 (n_100_43), .C2 (n_94_46) );
AOI211_X1 g_102_45 (.ZN (n_102_45), .A (n_102_43), .B (n_103_43), .C1 (n_102_42), .C2 (n_96_45) );
AOI211_X1 g_101_43 (.ZN (n_101_43), .A (n_100_44), .B (n_105_42), .C1 (n_104_41), .C2 (n_98_44) );
AOI211_X1 g_99_44 (.ZN (n_99_44), .A (n_102_45), .B (n_104_44), .C1 (n_103_43), .C2 (n_100_43) );
AOI211_X1 g_97_45 (.ZN (n_97_45), .A (n_101_43), .B (n_102_43), .C1 (n_105_42), .C2 (n_102_42) );
AOI211_X1 g_95_46 (.ZN (n_95_46), .A (n_99_44), .B (n_100_44), .C1 (n_104_44), .C2 (n_104_41) );
AOI211_X1 g_93_47 (.ZN (n_93_47), .A (n_97_45), .B (n_102_45), .C1 (n_102_43), .C2 (n_103_43) );
AOI211_X1 g_91_48 (.ZN (n_91_48), .A (n_95_46), .B (n_101_43), .C1 (n_100_44), .C2 (n_105_42) );
AOI211_X1 g_89_49 (.ZN (n_89_49), .A (n_93_47), .B (n_99_44), .C1 (n_102_45), .C2 (n_104_44) );
AOI211_X1 g_87_50 (.ZN (n_87_50), .A (n_91_48), .B (n_97_45), .C1 (n_101_43), .C2 (n_102_43) );
AOI211_X1 g_85_51 (.ZN (n_85_51), .A (n_89_49), .B (n_95_46), .C1 (n_99_44), .C2 (n_100_44) );
AOI211_X1 g_83_52 (.ZN (n_83_52), .A (n_87_50), .B (n_93_47), .C1 (n_97_45), .C2 (n_102_45) );
AOI211_X1 g_81_53 (.ZN (n_81_53), .A (n_85_51), .B (n_91_48), .C1 (n_95_46), .C2 (n_101_43) );
AOI211_X1 g_79_54 (.ZN (n_79_54), .A (n_83_52), .B (n_89_49), .C1 (n_93_47), .C2 (n_99_44) );
AOI211_X1 g_77_55 (.ZN (n_77_55), .A (n_81_53), .B (n_87_50), .C1 (n_91_48), .C2 (n_97_45) );
AOI211_X1 g_75_56 (.ZN (n_75_56), .A (n_79_54), .B (n_85_51), .C1 (n_89_49), .C2 (n_95_46) );
AOI211_X1 g_73_57 (.ZN (n_73_57), .A (n_77_55), .B (n_83_52), .C1 (n_87_50), .C2 (n_93_47) );
AOI211_X1 g_71_58 (.ZN (n_71_58), .A (n_75_56), .B (n_81_53), .C1 (n_85_51), .C2 (n_91_48) );
AOI211_X1 g_69_59 (.ZN (n_69_59), .A (n_73_57), .B (n_79_54), .C1 (n_83_52), .C2 (n_89_49) );
AOI211_X1 g_67_60 (.ZN (n_67_60), .A (n_71_58), .B (n_77_55), .C1 (n_81_53), .C2 (n_87_50) );
AOI211_X1 g_65_61 (.ZN (n_65_61), .A (n_69_59), .B (n_75_56), .C1 (n_79_54), .C2 (n_85_51) );
AOI211_X1 g_63_62 (.ZN (n_63_62), .A (n_67_60), .B (n_73_57), .C1 (n_77_55), .C2 (n_83_52) );
AOI211_X1 g_61_63 (.ZN (n_61_63), .A (n_65_61), .B (n_71_58), .C1 (n_75_56), .C2 (n_81_53) );
AOI211_X1 g_59_64 (.ZN (n_59_64), .A (n_63_62), .B (n_69_59), .C1 (n_73_57), .C2 (n_79_54) );
AOI211_X1 g_57_65 (.ZN (n_57_65), .A (n_61_63), .B (n_67_60), .C1 (n_71_58), .C2 (n_77_55) );
AOI211_X1 g_55_66 (.ZN (n_55_66), .A (n_59_64), .B (n_65_61), .C1 (n_69_59), .C2 (n_75_56) );
AOI211_X1 g_53_67 (.ZN (n_53_67), .A (n_57_65), .B (n_63_62), .C1 (n_67_60), .C2 (n_73_57) );
AOI211_X1 g_51_68 (.ZN (n_51_68), .A (n_55_66), .B (n_61_63), .C1 (n_65_61), .C2 (n_71_58) );
AOI211_X1 g_49_69 (.ZN (n_49_69), .A (n_53_67), .B (n_59_64), .C1 (n_63_62), .C2 (n_69_59) );
AOI211_X1 g_48_71 (.ZN (n_48_71), .A (n_51_68), .B (n_57_65), .C1 (n_61_63), .C2 (n_67_60) );
AOI211_X1 g_46_70 (.ZN (n_46_70), .A (n_49_69), .B (n_55_66), .C1 (n_59_64), .C2 (n_65_61) );
AOI211_X1 g_48_69 (.ZN (n_48_69), .A (n_48_71), .B (n_53_67), .C1 (n_57_65), .C2 (n_63_62) );
AOI211_X1 g_50_70 (.ZN (n_50_70), .A (n_46_70), .B (n_51_68), .C1 (n_55_66), .C2 (n_61_63) );
AOI211_X1 g_52_69 (.ZN (n_52_69), .A (n_48_69), .B (n_49_69), .C1 (n_53_67), .C2 (n_59_64) );
AOI211_X1 g_54_68 (.ZN (n_54_68), .A (n_50_70), .B (n_48_71), .C1 (n_51_68), .C2 (n_57_65) );
AOI211_X1 g_56_67 (.ZN (n_56_67), .A (n_52_69), .B (n_46_70), .C1 (n_49_69), .C2 (n_55_66) );
AOI211_X1 g_58_66 (.ZN (n_58_66), .A (n_54_68), .B (n_48_69), .C1 (n_48_71), .C2 (n_53_67) );
AOI211_X1 g_56_65 (.ZN (n_56_65), .A (n_56_67), .B (n_50_70), .C1 (n_46_70), .C2 (n_51_68) );
AOI211_X1 g_58_64 (.ZN (n_58_64), .A (n_58_66), .B (n_52_69), .C1 (n_48_69), .C2 (n_49_69) );
AOI211_X1 g_60_63 (.ZN (n_60_63), .A (n_56_65), .B (n_54_68), .C1 (n_50_70), .C2 (n_48_71) );
AOI211_X1 g_62_62 (.ZN (n_62_62), .A (n_58_64), .B (n_56_67), .C1 (n_52_69), .C2 (n_46_70) );
AOI211_X1 g_61_64 (.ZN (n_61_64), .A (n_60_63), .B (n_58_66), .C1 (n_54_68), .C2 (n_48_69) );
AOI211_X1 g_63_63 (.ZN (n_63_63), .A (n_62_62), .B (n_56_65), .C1 (n_56_67), .C2 (n_50_70) );
AOI211_X1 g_65_62 (.ZN (n_65_62), .A (n_61_64), .B (n_58_64), .C1 (n_58_66), .C2 (n_52_69) );
AOI211_X1 g_67_61 (.ZN (n_67_61), .A (n_63_63), .B (n_60_63), .C1 (n_56_65), .C2 (n_54_68) );
AOI211_X1 g_69_60 (.ZN (n_69_60), .A (n_65_62), .B (n_62_62), .C1 (n_58_64), .C2 (n_56_67) );
AOI211_X1 g_71_59 (.ZN (n_71_59), .A (n_67_61), .B (n_61_64), .C1 (n_60_63), .C2 (n_58_66) );
AOI211_X1 g_73_58 (.ZN (n_73_58), .A (n_69_60), .B (n_63_63), .C1 (n_62_62), .C2 (n_56_65) );
AOI211_X1 g_75_57 (.ZN (n_75_57), .A (n_71_59), .B (n_65_62), .C1 (n_61_64), .C2 (n_58_64) );
AOI211_X1 g_77_56 (.ZN (n_77_56), .A (n_73_58), .B (n_67_61), .C1 (n_63_63), .C2 (n_60_63) );
AOI211_X1 g_79_55 (.ZN (n_79_55), .A (n_75_57), .B (n_69_60), .C1 (n_65_62), .C2 (n_62_62) );
AOI211_X1 g_81_54 (.ZN (n_81_54), .A (n_77_56), .B (n_71_59), .C1 (n_67_61), .C2 (n_61_64) );
AOI211_X1 g_83_53 (.ZN (n_83_53), .A (n_79_55), .B (n_73_58), .C1 (n_69_60), .C2 (n_63_63) );
AOI211_X1 g_85_52 (.ZN (n_85_52), .A (n_81_54), .B (n_75_57), .C1 (n_71_59), .C2 (n_65_62) );
AOI211_X1 g_87_51 (.ZN (n_87_51), .A (n_83_53), .B (n_77_56), .C1 (n_73_58), .C2 (n_67_61) );
AOI211_X1 g_89_50 (.ZN (n_89_50), .A (n_85_52), .B (n_79_55), .C1 (n_75_57), .C2 (n_69_60) );
AOI211_X1 g_91_49 (.ZN (n_91_49), .A (n_87_51), .B (n_81_54), .C1 (n_77_56), .C2 (n_71_59) );
AOI211_X1 g_93_48 (.ZN (n_93_48), .A (n_89_50), .B (n_83_53), .C1 (n_79_55), .C2 (n_73_58) );
AOI211_X1 g_95_47 (.ZN (n_95_47), .A (n_91_49), .B (n_85_52), .C1 (n_81_54), .C2 (n_75_57) );
AOI211_X1 g_97_46 (.ZN (n_97_46), .A (n_93_48), .B (n_87_51), .C1 (n_83_53), .C2 (n_77_56) );
AOI211_X1 g_99_45 (.ZN (n_99_45), .A (n_95_47), .B (n_89_50), .C1 (n_85_52), .C2 (n_79_55) );
AOI211_X1 g_101_44 (.ZN (n_101_44), .A (n_97_46), .B (n_91_49), .C1 (n_87_51), .C2 (n_81_54) );
AOI211_X1 g_100_46 (.ZN (n_100_46), .A (n_99_45), .B (n_93_48), .C1 (n_89_50), .C2 (n_83_53) );
AOI211_X1 g_98_47 (.ZN (n_98_47), .A (n_101_44), .B (n_95_47), .C1 (n_91_49), .C2 (n_85_52) );
AOI211_X1 g_96_48 (.ZN (n_96_48), .A (n_100_46), .B (n_97_46), .C1 (n_93_48), .C2 (n_87_51) );
AOI211_X1 g_94_49 (.ZN (n_94_49), .A (n_98_47), .B (n_99_45), .C1 (n_95_47), .C2 (n_89_50) );
AOI211_X1 g_92_48 (.ZN (n_92_48), .A (n_96_48), .B (n_101_44), .C1 (n_97_46), .C2 (n_91_49) );
AOI211_X1 g_90_49 (.ZN (n_90_49), .A (n_94_49), .B (n_100_46), .C1 (n_99_45), .C2 (n_93_48) );
AOI211_X1 g_88_50 (.ZN (n_88_50), .A (n_92_48), .B (n_98_47), .C1 (n_101_44), .C2 (n_95_47) );
AOI211_X1 g_86_51 (.ZN (n_86_51), .A (n_90_49), .B (n_96_48), .C1 (n_100_46), .C2 (n_97_46) );
AOI211_X1 g_84_52 (.ZN (n_84_52), .A (n_88_50), .B (n_94_49), .C1 (n_98_47), .C2 (n_99_45) );
AOI211_X1 g_82_53 (.ZN (n_82_53), .A (n_86_51), .B (n_92_48), .C1 (n_96_48), .C2 (n_101_44) );
AOI211_X1 g_80_54 (.ZN (n_80_54), .A (n_84_52), .B (n_90_49), .C1 (n_94_49), .C2 (n_100_46) );
AOI211_X1 g_78_55 (.ZN (n_78_55), .A (n_82_53), .B (n_88_50), .C1 (n_92_48), .C2 (n_98_47) );
AOI211_X1 g_76_56 (.ZN (n_76_56), .A (n_80_54), .B (n_86_51), .C1 (n_90_49), .C2 (n_96_48) );
AOI211_X1 g_74_57 (.ZN (n_74_57), .A (n_78_55), .B (n_84_52), .C1 (n_88_50), .C2 (n_94_49) );
AOI211_X1 g_72_58 (.ZN (n_72_58), .A (n_76_56), .B (n_82_53), .C1 (n_86_51), .C2 (n_92_48) );
AOI211_X1 g_70_59 (.ZN (n_70_59), .A (n_74_57), .B (n_80_54), .C1 (n_84_52), .C2 (n_90_49) );
AOI211_X1 g_68_60 (.ZN (n_68_60), .A (n_72_58), .B (n_78_55), .C1 (n_82_53), .C2 (n_88_50) );
AOI211_X1 g_66_61 (.ZN (n_66_61), .A (n_70_59), .B (n_76_56), .C1 (n_80_54), .C2 (n_86_51) );
AOI211_X1 g_64_62 (.ZN (n_64_62), .A (n_68_60), .B (n_74_57), .C1 (n_78_55), .C2 (n_84_52) );
AOI211_X1 g_62_63 (.ZN (n_62_63), .A (n_66_61), .B (n_72_58), .C1 (n_76_56), .C2 (n_82_53) );
AOI211_X1 g_60_64 (.ZN (n_60_64), .A (n_64_62), .B (n_70_59), .C1 (n_74_57), .C2 (n_80_54) );
AOI211_X1 g_58_65 (.ZN (n_58_65), .A (n_62_63), .B (n_68_60), .C1 (n_72_58), .C2 (n_78_55) );
AOI211_X1 g_56_66 (.ZN (n_56_66), .A (n_60_64), .B (n_66_61), .C1 (n_70_59), .C2 (n_76_56) );
AOI211_X1 g_54_67 (.ZN (n_54_67), .A (n_58_65), .B (n_64_62), .C1 (n_68_60), .C2 (n_74_57) );
AOI211_X1 g_52_68 (.ZN (n_52_68), .A (n_56_66), .B (n_62_63), .C1 (n_66_61), .C2 (n_72_58) );
AOI211_X1 g_50_69 (.ZN (n_50_69), .A (n_54_67), .B (n_60_64), .C1 (n_64_62), .C2 (n_70_59) );
AOI211_X1 g_48_70 (.ZN (n_48_70), .A (n_52_68), .B (n_58_65), .C1 (n_62_63), .C2 (n_68_60) );
AOI211_X1 g_46_71 (.ZN (n_46_71), .A (n_50_69), .B (n_56_66), .C1 (n_60_64), .C2 (n_66_61) );
AOI211_X1 g_44_72 (.ZN (n_44_72), .A (n_48_70), .B (n_54_67), .C1 (n_58_65), .C2 (n_64_62) );
AOI211_X1 g_42_73 (.ZN (n_42_73), .A (n_46_71), .B (n_52_68), .C1 (n_56_66), .C2 (n_62_63) );
AOI211_X1 g_40_74 (.ZN (n_40_74), .A (n_44_72), .B (n_50_69), .C1 (n_54_67), .C2 (n_60_64) );
AOI211_X1 g_38_75 (.ZN (n_38_75), .A (n_42_73), .B (n_48_70), .C1 (n_52_68), .C2 (n_58_65) );
AOI211_X1 g_36_76 (.ZN (n_36_76), .A (n_40_74), .B (n_46_71), .C1 (n_50_69), .C2 (n_56_66) );
AOI211_X1 g_34_77 (.ZN (n_34_77), .A (n_38_75), .B (n_44_72), .C1 (n_48_70), .C2 (n_54_67) );
AOI211_X1 g_32_78 (.ZN (n_32_78), .A (n_36_76), .B (n_42_73), .C1 (n_46_71), .C2 (n_52_68) );
AOI211_X1 g_33_76 (.ZN (n_33_76), .A (n_34_77), .B (n_40_74), .C1 (n_44_72), .C2 (n_50_69) );
AOI211_X1 g_31_77 (.ZN (n_31_77), .A (n_32_78), .B (n_38_75), .C1 (n_42_73), .C2 (n_48_70) );
AOI211_X1 g_32_75 (.ZN (n_32_75), .A (n_33_76), .B (n_36_76), .C1 (n_40_74), .C2 (n_46_71) );
AOI211_X1 g_30_76 (.ZN (n_30_76), .A (n_31_77), .B (n_34_77), .C1 (n_38_75), .C2 (n_44_72) );
AOI211_X1 g_28_77 (.ZN (n_28_77), .A (n_32_75), .B (n_32_78), .C1 (n_36_76), .C2 (n_42_73) );
AOI211_X1 g_26_78 (.ZN (n_26_78), .A (n_30_76), .B (n_33_76), .C1 (n_34_77), .C2 (n_40_74) );
AOI211_X1 g_24_79 (.ZN (n_24_79), .A (n_28_77), .B (n_31_77), .C1 (n_32_78), .C2 (n_38_75) );
AOI211_X1 g_23_81 (.ZN (n_23_81), .A (n_26_78), .B (n_32_75), .C1 (n_33_76), .C2 (n_36_76) );
AOI211_X1 g_21_82 (.ZN (n_21_82), .A (n_24_79), .B (n_30_76), .C1 (n_31_77), .C2 (n_34_77) );
AOI211_X1 g_20_84 (.ZN (n_20_84), .A (n_23_81), .B (n_28_77), .C1 (n_32_75), .C2 (n_32_78) );
AOI211_X1 g_18_83 (.ZN (n_18_83), .A (n_21_82), .B (n_26_78), .C1 (n_30_76), .C2 (n_33_76) );
AOI211_X1 g_16_84 (.ZN (n_16_84), .A (n_20_84), .B (n_24_79), .C1 (n_28_77), .C2 (n_31_77) );
AOI211_X1 g_14_85 (.ZN (n_14_85), .A (n_18_83), .B (n_23_81), .C1 (n_26_78), .C2 (n_32_75) );
AOI211_X1 g_15_83 (.ZN (n_15_83), .A (n_16_84), .B (n_21_82), .C1 (n_24_79), .C2 (n_30_76) );
AOI211_X1 g_13_84 (.ZN (n_13_84), .A (n_14_85), .B (n_20_84), .C1 (n_23_81), .C2 (n_28_77) );
AOI211_X1 g_11_85 (.ZN (n_11_85), .A (n_15_83), .B (n_18_83), .C1 (n_21_82), .C2 (n_26_78) );
AOI211_X1 g_9_86 (.ZN (n_9_86), .A (n_13_84), .B (n_16_84), .C1 (n_20_84), .C2 (n_24_79) );
AOI211_X1 g_7_87 (.ZN (n_7_87), .A (n_11_85), .B (n_14_85), .C1 (n_18_83), .C2 (n_23_81) );
AOI211_X1 g_9_88 (.ZN (n_9_88), .A (n_9_86), .B (n_15_83), .C1 (n_16_84), .C2 (n_21_82) );
AOI211_X1 g_11_87 (.ZN (n_11_87), .A (n_7_87), .B (n_13_84), .C1 (n_14_85), .C2 (n_20_84) );
AOI211_X1 g_13_86 (.ZN (n_13_86), .A (n_9_88), .B (n_11_85), .C1 (n_15_83), .C2 (n_18_83) );
AOI211_X1 g_15_85 (.ZN (n_15_85), .A (n_11_87), .B (n_9_86), .C1 (n_13_84), .C2 (n_16_84) );
AOI211_X1 g_17_84 (.ZN (n_17_84), .A (n_13_86), .B (n_7_87), .C1 (n_11_85), .C2 (n_14_85) );
AOI211_X1 g_16_86 (.ZN (n_16_86), .A (n_15_85), .B (n_9_88), .C1 (n_9_86), .C2 (n_15_83) );
AOI211_X1 g_18_85 (.ZN (n_18_85), .A (n_17_84), .B (n_11_87), .C1 (n_7_87), .C2 (n_13_84) );
AOI211_X1 g_17_83 (.ZN (n_17_83), .A (n_16_86), .B (n_13_86), .C1 (n_9_88), .C2 (n_11_85) );
AOI211_X1 g_15_84 (.ZN (n_15_84), .A (n_18_85), .B (n_15_85), .C1 (n_11_87), .C2 (n_9_86) );
AOI211_X1 g_13_85 (.ZN (n_13_85), .A (n_17_83), .B (n_17_84), .C1 (n_13_86), .C2 (n_7_87) );
AOI211_X1 g_11_86 (.ZN (n_11_86), .A (n_15_84), .B (n_16_86), .C1 (n_15_85), .C2 (n_9_88) );
AOI211_X1 g_10_88 (.ZN (n_10_88), .A (n_13_85), .B (n_18_85), .C1 (n_17_84), .C2 (n_11_87) );
AOI211_X1 g_12_87 (.ZN (n_12_87), .A (n_11_86), .B (n_17_83), .C1 (n_16_86), .C2 (n_13_86) );
AOI211_X1 g_14_86 (.ZN (n_14_86), .A (n_10_88), .B (n_15_84), .C1 (n_18_85), .C2 (n_15_85) );
AOI211_X1 g_16_85 (.ZN (n_16_85), .A (n_12_87), .B (n_13_85), .C1 (n_17_83), .C2 (n_17_84) );
AOI211_X1 g_18_84 (.ZN (n_18_84), .A (n_14_86), .B (n_11_86), .C1 (n_15_84), .C2 (n_16_86) );
AOI211_X1 g_20_83 (.ZN (n_20_83), .A (n_16_85), .B (n_10_88), .C1 (n_13_85), .C2 (n_18_85) );
AOI211_X1 g_22_82 (.ZN (n_22_82), .A (n_18_84), .B (n_12_87), .C1 (n_11_86), .C2 (n_17_83) );
AOI211_X1 g_24_81 (.ZN (n_24_81), .A (n_20_83), .B (n_14_86), .C1 (n_10_88), .C2 (n_15_84) );
AOI211_X1 g_26_80 (.ZN (n_26_80), .A (n_22_82), .B (n_16_85), .C1 (n_12_87), .C2 (n_13_85) );
AOI211_X1 g_28_79 (.ZN (n_28_79), .A (n_24_81), .B (n_18_84), .C1 (n_14_86), .C2 (n_11_86) );
AOI211_X1 g_30_78 (.ZN (n_30_78), .A (n_26_80), .B (n_20_83), .C1 (n_16_85), .C2 (n_10_88) );
AOI211_X1 g_32_77 (.ZN (n_32_77), .A (n_28_79), .B (n_22_82), .C1 (n_18_84), .C2 (n_12_87) );
AOI211_X1 g_34_76 (.ZN (n_34_76), .A (n_30_78), .B (n_24_81), .C1 (n_20_83), .C2 (n_14_86) );
AOI211_X1 g_36_75 (.ZN (n_36_75), .A (n_32_77), .B (n_26_80), .C1 (n_22_82), .C2 (n_16_85) );
AOI211_X1 g_38_74 (.ZN (n_38_74), .A (n_34_76), .B (n_28_79), .C1 (n_24_81), .C2 (n_18_84) );
AOI211_X1 g_40_73 (.ZN (n_40_73), .A (n_36_75), .B (n_30_78), .C1 (n_26_80), .C2 (n_20_83) );
AOI211_X1 g_42_72 (.ZN (n_42_72), .A (n_38_74), .B (n_32_77), .C1 (n_28_79), .C2 (n_22_82) );
AOI211_X1 g_44_71 (.ZN (n_44_71), .A (n_40_73), .B (n_34_76), .C1 (n_30_78), .C2 (n_24_81) );
AOI211_X1 g_46_72 (.ZN (n_46_72), .A (n_42_72), .B (n_36_75), .C1 (n_32_77), .C2 (n_26_80) );
AOI211_X1 g_44_73 (.ZN (n_44_73), .A (n_44_71), .B (n_38_74), .C1 (n_34_76), .C2 (n_28_79) );
AOI211_X1 g_42_74 (.ZN (n_42_74), .A (n_46_72), .B (n_40_73), .C1 (n_36_75), .C2 (n_30_78) );
AOI211_X1 g_40_75 (.ZN (n_40_75), .A (n_44_73), .B (n_42_72), .C1 (n_38_74), .C2 (n_32_77) );
AOI211_X1 g_38_76 (.ZN (n_38_76), .A (n_42_74), .B (n_44_71), .C1 (n_40_73), .C2 (n_34_76) );
AOI211_X1 g_37_78 (.ZN (n_37_78), .A (n_40_75), .B (n_46_72), .C1 (n_42_72), .C2 (n_36_75) );
AOI211_X1 g_35_77 (.ZN (n_35_77), .A (n_38_76), .B (n_44_73), .C1 (n_44_71), .C2 (n_38_74) );
AOI211_X1 g_37_76 (.ZN (n_37_76), .A (n_37_78), .B (n_42_74), .C1 (n_46_72), .C2 (n_40_73) );
AOI211_X1 g_39_75 (.ZN (n_39_75), .A (n_35_77), .B (n_40_75), .C1 (n_44_73), .C2 (n_42_72) );
AOI211_X1 g_41_74 (.ZN (n_41_74), .A (n_37_76), .B (n_38_76), .C1 (n_42_74), .C2 (n_44_71) );
AOI211_X1 g_43_73 (.ZN (n_43_73), .A (n_39_75), .B (n_37_78), .C1 (n_40_75), .C2 (n_46_72) );
AOI211_X1 g_45_72 (.ZN (n_45_72), .A (n_41_74), .B (n_35_77), .C1 (n_38_76), .C2 (n_44_73) );
AOI211_X1 g_47_71 (.ZN (n_47_71), .A (n_43_73), .B (n_37_76), .C1 (n_37_78), .C2 (n_42_74) );
AOI211_X1 g_49_70 (.ZN (n_49_70), .A (n_45_72), .B (n_39_75), .C1 (n_35_77), .C2 (n_40_75) );
AOI211_X1 g_51_69 (.ZN (n_51_69), .A (n_47_71), .B (n_41_74), .C1 (n_37_76), .C2 (n_38_76) );
AOI211_X1 g_53_68 (.ZN (n_53_68), .A (n_49_70), .B (n_43_73), .C1 (n_39_75), .C2 (n_37_78) );
AOI211_X1 g_55_67 (.ZN (n_55_67), .A (n_51_69), .B (n_45_72), .C1 (n_41_74), .C2 (n_35_77) );
AOI211_X1 g_57_66 (.ZN (n_57_66), .A (n_53_68), .B (n_47_71), .C1 (n_43_73), .C2 (n_37_76) );
AOI211_X1 g_59_65 (.ZN (n_59_65), .A (n_55_67), .B (n_49_70), .C1 (n_45_72), .C2 (n_39_75) );
AOI211_X1 g_58_67 (.ZN (n_58_67), .A (n_57_66), .B (n_51_69), .C1 (n_47_71), .C2 (n_41_74) );
AOI211_X1 g_60_66 (.ZN (n_60_66), .A (n_59_65), .B (n_53_68), .C1 (n_49_70), .C2 (n_43_73) );
AOI211_X1 g_62_65 (.ZN (n_62_65), .A (n_58_67), .B (n_55_67), .C1 (n_51_69), .C2 (n_45_72) );
AOI211_X1 g_64_64 (.ZN (n_64_64), .A (n_60_66), .B (n_57_66), .C1 (n_53_68), .C2 (n_47_71) );
AOI211_X1 g_66_63 (.ZN (n_66_63), .A (n_62_65), .B (n_59_65), .C1 (n_55_67), .C2 (n_49_70) );
AOI211_X1 g_68_62 (.ZN (n_68_62), .A (n_64_64), .B (n_58_67), .C1 (n_57_66), .C2 (n_51_69) );
AOI211_X1 g_70_61 (.ZN (n_70_61), .A (n_66_63), .B (n_60_66), .C1 (n_59_65), .C2 (n_53_68) );
AOI211_X1 g_72_60 (.ZN (n_72_60), .A (n_68_62), .B (n_62_65), .C1 (n_58_67), .C2 (n_55_67) );
AOI211_X1 g_74_59 (.ZN (n_74_59), .A (n_70_61), .B (n_64_64), .C1 (n_60_66), .C2 (n_57_66) );
AOI211_X1 g_76_58 (.ZN (n_76_58), .A (n_72_60), .B (n_66_63), .C1 (n_62_65), .C2 (n_59_65) );
AOI211_X1 g_78_57 (.ZN (n_78_57), .A (n_74_59), .B (n_68_62), .C1 (n_64_64), .C2 (n_58_67) );
AOI211_X1 g_80_56 (.ZN (n_80_56), .A (n_76_58), .B (n_70_61), .C1 (n_66_63), .C2 (n_60_66) );
AOI211_X1 g_82_55 (.ZN (n_82_55), .A (n_78_57), .B (n_72_60), .C1 (n_68_62), .C2 (n_62_65) );
AOI211_X1 g_84_54 (.ZN (n_84_54), .A (n_80_56), .B (n_74_59), .C1 (n_70_61), .C2 (n_64_64) );
AOI211_X1 g_86_53 (.ZN (n_86_53), .A (n_82_55), .B (n_76_58), .C1 (n_72_60), .C2 (n_66_63) );
AOI211_X1 g_88_52 (.ZN (n_88_52), .A (n_84_54), .B (n_78_57), .C1 (n_74_59), .C2 (n_68_62) );
AOI211_X1 g_90_51 (.ZN (n_90_51), .A (n_86_53), .B (n_80_56), .C1 (n_76_58), .C2 (n_70_61) );
AOI211_X1 g_92_50 (.ZN (n_92_50), .A (n_88_52), .B (n_82_55), .C1 (n_78_57), .C2 (n_72_60) );
AOI211_X1 g_91_52 (.ZN (n_91_52), .A (n_90_51), .B (n_84_54), .C1 (n_80_56), .C2 (n_74_59) );
AOI211_X1 g_90_50 (.ZN (n_90_50), .A (n_92_50), .B (n_86_53), .C1 (n_82_55), .C2 (n_76_58) );
AOI211_X1 g_92_49 (.ZN (n_92_49), .A (n_91_52), .B (n_88_52), .C1 (n_84_54), .C2 (n_78_57) );
AOI211_X1 g_94_48 (.ZN (n_94_48), .A (n_90_50), .B (n_90_51), .C1 (n_86_53), .C2 (n_80_56) );
AOI211_X1 g_96_47 (.ZN (n_96_47), .A (n_92_49), .B (n_92_50), .C1 (n_88_52), .C2 (n_82_55) );
AOI211_X1 g_98_46 (.ZN (n_98_46), .A (n_94_48), .B (n_91_52), .C1 (n_90_51), .C2 (n_84_54) );
AOI211_X1 g_100_45 (.ZN (n_100_45), .A (n_96_47), .B (n_90_50), .C1 (n_92_50), .C2 (n_86_53) );
AOI211_X1 g_102_44 (.ZN (n_102_44), .A (n_98_46), .B (n_92_49), .C1 (n_91_52), .C2 (n_88_52) );
AOI211_X1 g_104_43 (.ZN (n_104_43), .A (n_100_45), .B (n_94_48), .C1 (n_90_50), .C2 (n_90_51) );
AOI211_X1 g_106_42 (.ZN (n_106_42), .A (n_102_44), .B (n_96_47), .C1 (n_92_49), .C2 (n_92_50) );
AOI211_X1 g_108_41 (.ZN (n_108_41), .A (n_104_43), .B (n_98_46), .C1 (n_94_48), .C2 (n_91_52) );
AOI211_X1 g_110_40 (.ZN (n_110_40), .A (n_106_42), .B (n_100_45), .C1 (n_96_47), .C2 (n_90_50) );
AOI211_X1 g_109_42 (.ZN (n_109_42), .A (n_108_41), .B (n_102_44), .C1 (n_98_46), .C2 (n_92_49) );
AOI211_X1 g_108_40 (.ZN (n_108_40), .A (n_110_40), .B (n_104_43), .C1 (n_100_45), .C2 (n_94_48) );
AOI211_X1 g_110_39 (.ZN (n_110_39), .A (n_109_42), .B (n_106_42), .C1 (n_102_44), .C2 (n_96_47) );
AOI211_X1 g_112_38 (.ZN (n_112_38), .A (n_108_40), .B (n_108_41), .C1 (n_104_43), .C2 (n_98_46) );
AOI211_X1 g_114_37 (.ZN (n_114_37), .A (n_110_39), .B (n_110_40), .C1 (n_106_42), .C2 (n_100_45) );
AOI211_X1 g_116_36 (.ZN (n_116_36), .A (n_112_38), .B (n_109_42), .C1 (n_108_41), .C2 (n_102_44) );
AOI211_X1 g_118_35 (.ZN (n_118_35), .A (n_114_37), .B (n_108_40), .C1 (n_110_40), .C2 (n_104_43) );
AOI211_X1 g_120_34 (.ZN (n_120_34), .A (n_116_36), .B (n_110_39), .C1 (n_109_42), .C2 (n_106_42) );
AOI211_X1 g_122_33 (.ZN (n_122_33), .A (n_118_35), .B (n_112_38), .C1 (n_108_40), .C2 (n_108_41) );
AOI211_X1 g_124_32 (.ZN (n_124_32), .A (n_120_34), .B (n_114_37), .C1 (n_110_39), .C2 (n_110_40) );
AOI211_X1 g_126_31 (.ZN (n_126_31), .A (n_122_33), .B (n_116_36), .C1 (n_112_38), .C2 (n_109_42) );
AOI211_X1 g_128_30 (.ZN (n_128_30), .A (n_124_32), .B (n_118_35), .C1 (n_114_37), .C2 (n_108_40) );
AOI211_X1 g_130_29 (.ZN (n_130_29), .A (n_126_31), .B (n_120_34), .C1 (n_116_36), .C2 (n_110_39) );
AOI211_X1 g_132_28 (.ZN (n_132_28), .A (n_128_30), .B (n_122_33), .C1 (n_118_35), .C2 (n_112_38) );
AOI211_X1 g_134_29 (.ZN (n_134_29), .A (n_130_29), .B (n_124_32), .C1 (n_120_34), .C2 (n_114_37) );
AOI211_X1 g_132_30 (.ZN (n_132_30), .A (n_132_28), .B (n_126_31), .C1 (n_122_33), .C2 (n_116_36) );
AOI211_X1 g_130_31 (.ZN (n_130_31), .A (n_134_29), .B (n_128_30), .C1 (n_124_32), .C2 (n_118_35) );
AOI211_X1 g_128_32 (.ZN (n_128_32), .A (n_132_30), .B (n_130_29), .C1 (n_126_31), .C2 (n_120_34) );
AOI211_X1 g_126_33 (.ZN (n_126_33), .A (n_130_31), .B (n_132_28), .C1 (n_128_30), .C2 (n_122_33) );
AOI211_X1 g_127_31 (.ZN (n_127_31), .A (n_128_32), .B (n_134_29), .C1 (n_130_29), .C2 (n_124_32) );
AOI211_X1 g_125_32 (.ZN (n_125_32), .A (n_126_33), .B (n_132_30), .C1 (n_132_28), .C2 (n_126_31) );
AOI211_X1 g_123_33 (.ZN (n_123_33), .A (n_127_31), .B (n_130_31), .C1 (n_134_29), .C2 (n_128_30) );
AOI211_X1 g_121_34 (.ZN (n_121_34), .A (n_125_32), .B (n_128_32), .C1 (n_132_30), .C2 (n_130_29) );
AOI211_X1 g_119_35 (.ZN (n_119_35), .A (n_123_33), .B (n_126_33), .C1 (n_130_31), .C2 (n_132_28) );
AOI211_X1 g_120_33 (.ZN (n_120_33), .A (n_121_34), .B (n_127_31), .C1 (n_128_32), .C2 (n_134_29) );
AOI211_X1 g_118_34 (.ZN (n_118_34), .A (n_119_35), .B (n_125_32), .C1 (n_126_33), .C2 (n_132_30) );
AOI211_X1 g_116_35 (.ZN (n_116_35), .A (n_120_33), .B (n_123_33), .C1 (n_127_31), .C2 (n_130_31) );
AOI211_X1 g_118_36 (.ZN (n_118_36), .A (n_118_34), .B (n_121_34), .C1 (n_125_32), .C2 (n_128_32) );
AOI211_X1 g_120_35 (.ZN (n_120_35), .A (n_116_35), .B (n_119_35), .C1 (n_123_33), .C2 (n_126_33) );
AOI211_X1 g_122_34 (.ZN (n_122_34), .A (n_118_36), .B (n_120_33), .C1 (n_121_34), .C2 (n_127_31) );
AOI211_X1 g_121_36 (.ZN (n_121_36), .A (n_120_35), .B (n_118_34), .C1 (n_119_35), .C2 (n_125_32) );
AOI211_X1 g_123_35 (.ZN (n_123_35), .A (n_122_34), .B (n_116_35), .C1 (n_120_33), .C2 (n_123_33) );
AOI211_X1 g_125_34 (.ZN (n_125_34), .A (n_121_36), .B (n_118_36), .C1 (n_118_34), .C2 (n_121_34) );
AOI211_X1 g_127_33 (.ZN (n_127_33), .A (n_123_35), .B (n_120_35), .C1 (n_116_35), .C2 (n_119_35) );
AOI211_X1 g_129_32 (.ZN (n_129_32), .A (n_125_34), .B (n_122_34), .C1 (n_118_36), .C2 (n_120_33) );
AOI211_X1 g_131_31 (.ZN (n_131_31), .A (n_127_33), .B (n_121_36), .C1 (n_120_35), .C2 (n_118_34) );
AOI211_X1 g_133_30 (.ZN (n_133_30), .A (n_129_32), .B (n_123_35), .C1 (n_122_34), .C2 (n_116_35) );
AOI211_X1 g_135_29 (.ZN (n_135_29), .A (n_131_31), .B (n_125_34), .C1 (n_121_36), .C2 (n_118_36) );
AOI211_X1 g_137_28 (.ZN (n_137_28), .A (n_133_30), .B (n_127_33), .C1 (n_123_35), .C2 (n_120_35) );
AOI211_X1 g_139_27 (.ZN (n_139_27), .A (n_135_29), .B (n_129_32), .C1 (n_125_34), .C2 (n_122_34) );
AOI211_X1 g_141_26 (.ZN (n_141_26), .A (n_137_28), .B (n_131_31), .C1 (n_127_33), .C2 (n_121_36) );
AOI211_X1 g_142_24 (.ZN (n_142_24), .A (n_139_27), .B (n_133_30), .C1 (n_129_32), .C2 (n_123_35) );
AOI211_X1 g_144_23 (.ZN (n_144_23), .A (n_141_26), .B (n_135_29), .C1 (n_131_31), .C2 (n_125_34) );
AOI211_X1 g_146_22 (.ZN (n_146_22), .A (n_142_24), .B (n_137_28), .C1 (n_133_30), .C2 (n_127_33) );
AOI211_X1 g_147_24 (.ZN (n_147_24), .A (n_144_23), .B (n_139_27), .C1 (n_135_29), .C2 (n_129_32) );
AOI211_X1 g_149_25 (.ZN (n_149_25), .A (n_146_22), .B (n_141_26), .C1 (n_137_28), .C2 (n_131_31) );
AOI211_X1 g_148_23 (.ZN (n_148_23), .A (n_147_24), .B (n_142_24), .C1 (n_139_27), .C2 (n_133_30) );
AOI211_X1 g_146_24 (.ZN (n_146_24), .A (n_149_25), .B (n_144_23), .C1 (n_141_26), .C2 (n_135_29) );
AOI211_X1 g_144_25 (.ZN (n_144_25), .A (n_148_23), .B (n_146_22), .C1 (n_142_24), .C2 (n_137_28) );
AOI211_X1 g_143_27 (.ZN (n_143_27), .A (n_146_24), .B (n_147_24), .C1 (n_144_23), .C2 (n_139_27) );
AOI211_X1 g_145_26 (.ZN (n_145_26), .A (n_144_25), .B (n_149_25), .C1 (n_146_22), .C2 (n_141_26) );
AOI211_X1 g_147_25 (.ZN (n_147_25), .A (n_143_27), .B (n_148_23), .C1 (n_147_24), .C2 (n_142_24) );
AOI211_X1 g_145_24 (.ZN (n_145_24), .A (n_145_26), .B (n_146_24), .C1 (n_149_25), .C2 (n_144_23) );
AOI211_X1 g_143_25 (.ZN (n_143_25), .A (n_147_25), .B (n_144_25), .C1 (n_148_23), .C2 (n_146_22) );
AOI211_X1 g_142_27 (.ZN (n_142_27), .A (n_145_24), .B (n_143_27), .C1 (n_146_24), .C2 (n_147_24) );
AOI211_X1 g_144_26 (.ZN (n_144_26), .A (n_143_25), .B (n_145_26), .C1 (n_144_25), .C2 (n_149_25) );
AOI211_X1 g_146_27 (.ZN (n_146_27), .A (n_142_27), .B (n_147_25), .C1 (n_143_27), .C2 (n_148_23) );
AOI211_X1 g_145_25 (.ZN (n_145_25), .A (n_144_26), .B (n_145_24), .C1 (n_145_26), .C2 (n_146_24) );
AOI211_X1 g_147_26 (.ZN (n_147_26), .A (n_146_27), .B (n_143_25), .C1 (n_147_25), .C2 (n_144_25) );
AOI211_X1 g_145_27 (.ZN (n_145_27), .A (n_145_25), .B (n_142_27), .C1 (n_145_24), .C2 (n_143_27) );
AOI211_X1 g_143_26 (.ZN (n_143_26), .A (n_147_26), .B (n_144_26), .C1 (n_143_25), .C2 (n_145_26) );
AOI211_X1 g_144_28 (.ZN (n_144_28), .A (n_145_27), .B (n_146_27), .C1 (n_142_27), .C2 (n_147_25) );
AOI211_X1 g_142_29 (.ZN (n_142_29), .A (n_143_26), .B (n_145_25), .C1 (n_144_26), .C2 (n_145_24) );
AOI211_X1 g_141_27 (.ZN (n_141_27), .A (n_144_28), .B (n_147_26), .C1 (n_146_27), .C2 (n_143_25) );
AOI211_X1 g_139_28 (.ZN (n_139_28), .A (n_142_29), .B (n_145_27), .C1 (n_145_25), .C2 (n_142_27) );
AOI211_X1 g_138_30 (.ZN (n_138_30), .A (n_141_27), .B (n_143_26), .C1 (n_147_26), .C2 (n_144_26) );
AOI211_X1 g_140_29 (.ZN (n_140_29), .A (n_139_28), .B (n_144_28), .C1 (n_145_27), .C2 (n_146_27) );
AOI211_X1 g_142_28 (.ZN (n_142_28), .A (n_138_30), .B (n_142_29), .C1 (n_143_26), .C2 (n_145_25) );
AOI211_X1 g_144_27 (.ZN (n_144_27), .A (n_140_29), .B (n_141_27), .C1 (n_144_28), .C2 (n_147_26) );
AOI211_X1 g_146_26 (.ZN (n_146_26), .A (n_142_28), .B (n_139_28), .C1 (n_142_29), .C2 (n_145_27) );
AOI211_X1 g_147_28 (.ZN (n_147_28), .A (n_144_27), .B (n_138_30), .C1 (n_141_27), .C2 (n_143_26) );
AOI211_X1 g_149_29 (.ZN (n_149_29), .A (n_146_26), .B (n_140_29), .C1 (n_139_28), .C2 (n_144_28) );
AOI211_X1 g_148_27 (.ZN (n_148_27), .A (n_147_28), .B (n_142_28), .C1 (n_138_30), .C2 (n_142_29) );
AOI211_X1 g_146_28 (.ZN (n_146_28), .A (n_149_29), .B (n_144_27), .C1 (n_140_29), .C2 (n_141_27) );
AOI211_X1 g_147_30 (.ZN (n_147_30), .A (n_148_27), .B (n_146_26), .C1 (n_142_28), .C2 (n_139_28) );
AOI211_X1 g_145_29 (.ZN (n_145_29), .A (n_146_28), .B (n_147_28), .C1 (n_144_27), .C2 (n_138_30) );
AOI211_X1 g_143_28 (.ZN (n_143_28), .A (n_147_30), .B (n_149_29), .C1 (n_146_26), .C2 (n_140_29) );
AOI211_X1 g_141_29 (.ZN (n_141_29), .A (n_145_29), .B (n_148_27), .C1 (n_147_28), .C2 (n_142_28) );
AOI211_X1 g_143_30 (.ZN (n_143_30), .A (n_143_28), .B (n_146_28), .C1 (n_149_29), .C2 (n_144_27) );
AOI211_X1 g_145_31 (.ZN (n_145_31), .A (n_141_29), .B (n_147_30), .C1 (n_148_27), .C2 (n_146_26) );
AOI211_X1 g_144_29 (.ZN (n_144_29), .A (n_143_30), .B (n_145_29), .C1 (n_146_28), .C2 (n_147_28) );
AOI211_X1 g_142_30 (.ZN (n_142_30), .A (n_145_31), .B (n_143_28), .C1 (n_147_30), .C2 (n_149_29) );
AOI211_X1 g_141_28 (.ZN (n_141_28), .A (n_144_29), .B (n_141_29), .C1 (n_145_29), .C2 (n_148_27) );
AOI211_X1 g_139_29 (.ZN (n_139_29), .A (n_142_30), .B (n_143_30), .C1 (n_143_28), .C2 (n_146_28) );
AOI211_X1 g_137_30 (.ZN (n_137_30), .A (n_141_28), .B (n_145_31), .C1 (n_141_29), .C2 (n_147_30) );
AOI211_X1 g_135_31 (.ZN (n_135_31), .A (n_139_29), .B (n_144_29), .C1 (n_143_30), .C2 (n_145_29) );
AOI211_X1 g_133_32 (.ZN (n_133_32), .A (n_137_30), .B (n_142_30), .C1 (n_145_31), .C2 (n_143_28) );
AOI211_X1 g_134_30 (.ZN (n_134_30), .A (n_135_31), .B (n_141_28), .C1 (n_144_29), .C2 (n_141_29) );
AOI211_X1 g_136_31 (.ZN (n_136_31), .A (n_133_32), .B (n_139_29), .C1 (n_142_30), .C2 (n_143_30) );
AOI211_X1 g_134_32 (.ZN (n_134_32), .A (n_134_30), .B (n_137_30), .C1 (n_141_28), .C2 (n_145_31) );
AOI211_X1 g_135_30 (.ZN (n_135_30), .A (n_136_31), .B (n_135_31), .C1 (n_139_29), .C2 (n_144_29) );
AOI211_X1 g_133_29 (.ZN (n_133_29), .A (n_134_32), .B (n_133_32), .C1 (n_137_30), .C2 (n_142_30) );
AOI211_X1 g_132_31 (.ZN (n_132_31), .A (n_135_30), .B (n_134_30), .C1 (n_135_31), .C2 (n_141_28) );
AOI211_X1 g_131_33 (.ZN (n_131_33), .A (n_133_29), .B (n_136_31), .C1 (n_133_32), .C2 (n_139_29) );
AOI211_X1 g_129_34 (.ZN (n_129_34), .A (n_132_31), .B (n_134_32), .C1 (n_134_30), .C2 (n_137_30) );
AOI211_X1 g_130_32 (.ZN (n_130_32), .A (n_131_33), .B (n_135_30), .C1 (n_136_31), .C2 (n_135_31) );
AOI211_X1 g_131_30 (.ZN (n_131_30), .A (n_129_34), .B (n_133_29), .C1 (n_134_32), .C2 (n_133_32) );
AOI211_X1 g_129_31 (.ZN (n_129_31), .A (n_130_32), .B (n_132_31), .C1 (n_135_30), .C2 (n_134_30) );
AOI211_X1 g_127_32 (.ZN (n_127_32), .A (n_131_30), .B (n_131_33), .C1 (n_133_29), .C2 (n_136_31) );
AOI211_X1 g_125_33 (.ZN (n_125_33), .A (n_129_31), .B (n_129_34), .C1 (n_132_31), .C2 (n_134_32) );
AOI211_X1 g_123_34 (.ZN (n_123_34), .A (n_127_32), .B (n_130_32), .C1 (n_131_33), .C2 (n_135_30) );
AOI211_X1 g_121_35 (.ZN (n_121_35), .A (n_125_33), .B (n_131_30), .C1 (n_129_34), .C2 (n_133_29) );
AOI211_X1 g_119_36 (.ZN (n_119_36), .A (n_123_34), .B (n_129_31), .C1 (n_130_32), .C2 (n_132_31) );
AOI211_X1 g_117_37 (.ZN (n_117_37), .A (n_121_35), .B (n_127_32), .C1 (n_131_30), .C2 (n_131_33) );
AOI211_X1 g_115_38 (.ZN (n_115_38), .A (n_119_36), .B (n_125_33), .C1 (n_129_31), .C2 (n_129_34) );
AOI211_X1 g_113_39 (.ZN (n_113_39), .A (n_117_37), .B (n_123_34), .C1 (n_127_32), .C2 (n_130_32) );
AOI211_X1 g_111_40 (.ZN (n_111_40), .A (n_115_38), .B (n_121_35), .C1 (n_125_33), .C2 (n_131_30) );
AOI211_X1 g_109_41 (.ZN (n_109_41), .A (n_113_39), .B (n_119_36), .C1 (n_123_34), .C2 (n_129_31) );
AOI211_X1 g_107_42 (.ZN (n_107_42), .A (n_111_40), .B (n_117_37), .C1 (n_121_35), .C2 (n_127_32) );
AOI211_X1 g_105_43 (.ZN (n_105_43), .A (n_109_41), .B (n_115_38), .C1 (n_119_36), .C2 (n_125_33) );
AOI211_X1 g_106_41 (.ZN (n_106_41), .A (n_107_42), .B (n_113_39), .C1 (n_117_37), .C2 (n_123_34) );
AOI211_X1 g_104_42 (.ZN (n_104_42), .A (n_105_43), .B (n_111_40), .C1 (n_115_38), .C2 (n_121_35) );
AOI211_X1 g_103_44 (.ZN (n_103_44), .A (n_106_41), .B (n_109_41), .C1 (n_113_39), .C2 (n_119_36) );
AOI211_X1 g_101_45 (.ZN (n_101_45), .A (n_104_42), .B (n_107_42), .C1 (n_111_40), .C2 (n_117_37) );
AOI211_X1 g_99_46 (.ZN (n_99_46), .A (n_103_44), .B (n_105_43), .C1 (n_109_41), .C2 (n_115_38) );
AOI211_X1 g_97_47 (.ZN (n_97_47), .A (n_101_45), .B (n_106_41), .C1 (n_107_42), .C2 (n_113_39) );
AOI211_X1 g_95_48 (.ZN (n_95_48), .A (n_99_46), .B (n_104_42), .C1 (n_105_43), .C2 (n_111_40) );
AOI211_X1 g_93_49 (.ZN (n_93_49), .A (n_97_47), .B (n_103_44), .C1 (n_106_41), .C2 (n_109_41) );
AOI211_X1 g_91_50 (.ZN (n_91_50), .A (n_95_48), .B (n_101_45), .C1 (n_104_42), .C2 (n_107_42) );
AOI211_X1 g_89_51 (.ZN (n_89_51), .A (n_93_49), .B (n_99_46), .C1 (n_103_44), .C2 (n_105_43) );
AOI211_X1 g_87_52 (.ZN (n_87_52), .A (n_91_50), .B (n_97_47), .C1 (n_101_45), .C2 (n_106_41) );
AOI211_X1 g_85_53 (.ZN (n_85_53), .A (n_89_51), .B (n_95_48), .C1 (n_99_46), .C2 (n_104_42) );
AOI211_X1 g_83_54 (.ZN (n_83_54), .A (n_87_52), .B (n_93_49), .C1 (n_97_47), .C2 (n_103_44) );
AOI211_X1 g_81_55 (.ZN (n_81_55), .A (n_85_53), .B (n_91_50), .C1 (n_95_48), .C2 (n_101_45) );
AOI211_X1 g_79_56 (.ZN (n_79_56), .A (n_83_54), .B (n_89_51), .C1 (n_93_49), .C2 (n_99_46) );
AOI211_X1 g_77_57 (.ZN (n_77_57), .A (n_81_55), .B (n_87_52), .C1 (n_91_50), .C2 (n_97_47) );
AOI211_X1 g_75_58 (.ZN (n_75_58), .A (n_79_56), .B (n_85_53), .C1 (n_89_51), .C2 (n_95_48) );
AOI211_X1 g_73_59 (.ZN (n_73_59), .A (n_77_57), .B (n_83_54), .C1 (n_87_52), .C2 (n_93_49) );
AOI211_X1 g_71_60 (.ZN (n_71_60), .A (n_75_58), .B (n_81_55), .C1 (n_85_53), .C2 (n_91_50) );
AOI211_X1 g_69_61 (.ZN (n_69_61), .A (n_73_59), .B (n_79_56), .C1 (n_83_54), .C2 (n_89_51) );
AOI211_X1 g_67_62 (.ZN (n_67_62), .A (n_71_60), .B (n_77_57), .C1 (n_81_55), .C2 (n_87_52) );
AOI211_X1 g_65_63 (.ZN (n_65_63), .A (n_69_61), .B (n_75_58), .C1 (n_79_56), .C2 (n_85_53) );
AOI211_X1 g_63_64 (.ZN (n_63_64), .A (n_67_62), .B (n_73_59), .C1 (n_77_57), .C2 (n_83_54) );
AOI211_X1 g_61_65 (.ZN (n_61_65), .A (n_65_63), .B (n_71_60), .C1 (n_75_58), .C2 (n_81_55) );
AOI211_X1 g_59_66 (.ZN (n_59_66), .A (n_63_64), .B (n_69_61), .C1 (n_73_59), .C2 (n_79_56) );
AOI211_X1 g_57_67 (.ZN (n_57_67), .A (n_61_65), .B (n_67_62), .C1 (n_71_60), .C2 (n_77_57) );
AOI211_X1 g_55_68 (.ZN (n_55_68), .A (n_59_66), .B (n_65_63), .C1 (n_69_61), .C2 (n_75_58) );
AOI211_X1 g_53_69 (.ZN (n_53_69), .A (n_57_67), .B (n_63_64), .C1 (n_67_62), .C2 (n_73_59) );
AOI211_X1 g_51_70 (.ZN (n_51_70), .A (n_55_68), .B (n_61_65), .C1 (n_65_63), .C2 (n_71_60) );
AOI211_X1 g_49_71 (.ZN (n_49_71), .A (n_53_69), .B (n_59_66), .C1 (n_63_64), .C2 (n_69_61) );
AOI211_X1 g_47_72 (.ZN (n_47_72), .A (n_51_70), .B (n_57_67), .C1 (n_61_65), .C2 (n_67_62) );
AOI211_X1 g_45_73 (.ZN (n_45_73), .A (n_49_71), .B (n_55_68), .C1 (n_59_66), .C2 (n_65_63) );
AOI211_X1 g_43_74 (.ZN (n_43_74), .A (n_47_72), .B (n_53_69), .C1 (n_57_67), .C2 (n_63_64) );
AOI211_X1 g_41_75 (.ZN (n_41_75), .A (n_45_73), .B (n_51_70), .C1 (n_55_68), .C2 (n_61_65) );
AOI211_X1 g_39_76 (.ZN (n_39_76), .A (n_43_74), .B (n_49_71), .C1 (n_53_69), .C2 (n_59_66) );
AOI211_X1 g_37_77 (.ZN (n_37_77), .A (n_41_75), .B (n_47_72), .C1 (n_51_70), .C2 (n_57_67) );
AOI211_X1 g_35_78 (.ZN (n_35_78), .A (n_39_76), .B (n_45_73), .C1 (n_49_71), .C2 (n_55_68) );
AOI211_X1 g_33_77 (.ZN (n_33_77), .A (n_37_77), .B (n_43_74), .C1 (n_47_72), .C2 (n_53_69) );
AOI211_X1 g_31_78 (.ZN (n_31_78), .A (n_35_78), .B (n_41_75), .C1 (n_45_73), .C2 (n_51_70) );
AOI211_X1 g_29_79 (.ZN (n_29_79), .A (n_33_77), .B (n_39_76), .C1 (n_43_74), .C2 (n_49_71) );
AOI211_X1 g_27_80 (.ZN (n_27_80), .A (n_31_78), .B (n_37_77), .C1 (n_41_75), .C2 (n_47_72) );
AOI211_X1 g_25_81 (.ZN (n_25_81), .A (n_29_79), .B (n_35_78), .C1 (n_39_76), .C2 (n_45_73) );
AOI211_X1 g_23_82 (.ZN (n_23_82), .A (n_27_80), .B (n_33_77), .C1 (n_37_77), .C2 (n_43_74) );
AOI211_X1 g_21_83 (.ZN (n_21_83), .A (n_25_81), .B (n_31_78), .C1 (n_35_78), .C2 (n_41_75) );
AOI211_X1 g_19_84 (.ZN (n_19_84), .A (n_23_82), .B (n_29_79), .C1 (n_33_77), .C2 (n_39_76) );
AOI211_X1 g_17_85 (.ZN (n_17_85), .A (n_21_83), .B (n_27_80), .C1 (n_31_78), .C2 (n_37_77) );
AOI211_X1 g_15_86 (.ZN (n_15_86), .A (n_19_84), .B (n_25_81), .C1 (n_29_79), .C2 (n_35_78) );
AOI211_X1 g_13_87 (.ZN (n_13_87), .A (n_17_85), .B (n_23_82), .C1 (n_27_80), .C2 (n_33_77) );
AOI211_X1 g_11_88 (.ZN (n_11_88), .A (n_15_86), .B (n_21_83), .C1 (n_25_81), .C2 (n_31_78) );
AOI211_X1 g_12_86 (.ZN (n_12_86), .A (n_13_87), .B (n_19_84), .C1 (n_23_82), .C2 (n_29_79) );
AOI211_X1 g_10_87 (.ZN (n_10_87), .A (n_11_88), .B (n_17_85), .C1 (n_21_83), .C2 (n_27_80) );
AOI211_X1 g_8_88 (.ZN (n_8_88), .A (n_12_86), .B (n_15_86), .C1 (n_19_84), .C2 (n_25_81) );
AOI211_X1 g_7_90 (.ZN (n_7_90), .A (n_10_87), .B (n_13_87), .C1 (n_17_85), .C2 (n_23_82) );
AOI211_X1 g_9_89 (.ZN (n_9_89), .A (n_8_88), .B (n_11_88), .C1 (n_15_86), .C2 (n_21_83) );
AOI211_X1 g_8_91 (.ZN (n_8_91), .A (n_7_90), .B (n_12_86), .C1 (n_13_87), .C2 (n_19_84) );
AOI211_X1 g_6_90 (.ZN (n_6_90), .A (n_9_89), .B (n_10_87), .C1 (n_11_88), .C2 (n_17_85) );
AOI211_X1 g_8_89 (.ZN (n_8_89), .A (n_8_91), .B (n_8_88), .C1 (n_12_86), .C2 (n_15_86) );
AOI211_X1 g_10_90 (.ZN (n_10_90), .A (n_6_90), .B (n_7_90), .C1 (n_10_87), .C2 (n_13_87) );
AOI211_X1 g_12_89 (.ZN (n_12_89), .A (n_8_89), .B (n_9_89), .C1 (n_8_88), .C2 (n_11_88) );
AOI211_X1 g_14_88 (.ZN (n_14_88), .A (n_10_90), .B (n_8_91), .C1 (n_7_90), .C2 (n_12_86) );
AOI211_X1 g_16_87 (.ZN (n_16_87), .A (n_12_89), .B (n_6_90), .C1 (n_9_89), .C2 (n_10_87) );
AOI211_X1 g_18_86 (.ZN (n_18_86), .A (n_14_88), .B (n_8_89), .C1 (n_8_91), .C2 (n_8_88) );
AOI211_X1 g_20_85 (.ZN (n_20_85), .A (n_16_87), .B (n_10_90), .C1 (n_6_90), .C2 (n_7_90) );
AOI211_X1 g_22_84 (.ZN (n_22_84), .A (n_18_86), .B (n_12_89), .C1 (n_8_89), .C2 (n_9_89) );
AOI211_X1 g_24_83 (.ZN (n_24_83), .A (n_20_85), .B (n_14_88), .C1 (n_10_90), .C2 (n_8_91) );
AOI211_X1 g_26_82 (.ZN (n_26_82), .A (n_22_84), .B (n_16_87), .C1 (n_12_89), .C2 (n_6_90) );
AOI211_X1 g_25_80 (.ZN (n_25_80), .A (n_24_83), .B (n_18_86), .C1 (n_14_88), .C2 (n_8_89) );
AOI211_X1 g_27_79 (.ZN (n_27_79), .A (n_26_82), .B (n_20_85), .C1 (n_16_87), .C2 (n_10_90) );
AOI211_X1 g_29_78 (.ZN (n_29_78), .A (n_25_80), .B (n_22_84), .C1 (n_18_86), .C2 (n_12_89) );
AOI211_X1 g_28_80 (.ZN (n_28_80), .A (n_27_79), .B (n_24_83), .C1 (n_20_85), .C2 (n_14_88) );
AOI211_X1 g_30_79 (.ZN (n_30_79), .A (n_29_78), .B (n_26_82), .C1 (n_22_84), .C2 (n_16_87) );
AOI211_X1 g_29_81 (.ZN (n_29_81), .A (n_28_80), .B (n_25_80), .C1 (n_24_83), .C2 (n_18_86) );
AOI211_X1 g_31_80 (.ZN (n_31_80), .A (n_30_79), .B (n_27_79), .C1 (n_26_82), .C2 (n_20_85) );
AOI211_X1 g_33_79 (.ZN (n_33_79), .A (n_29_81), .B (n_29_78), .C1 (n_25_80), .C2 (n_22_84) );
AOI211_X1 g_32_81 (.ZN (n_32_81), .A (n_31_80), .B (n_28_80), .C1 (n_27_79), .C2 (n_24_83) );
AOI211_X1 g_31_79 (.ZN (n_31_79), .A (n_33_79), .B (n_30_79), .C1 (n_29_78), .C2 (n_26_82) );
AOI211_X1 g_33_78 (.ZN (n_33_78), .A (n_32_81), .B (n_29_81), .C1 (n_28_80), .C2 (n_25_80) );
AOI211_X1 g_35_79 (.ZN (n_35_79), .A (n_31_79), .B (n_31_80), .C1 (n_30_79), .C2 (n_27_79) );
AOI211_X1 g_33_80 (.ZN (n_33_80), .A (n_33_78), .B (n_33_79), .C1 (n_29_81), .C2 (n_29_78) );
AOI211_X1 g_34_78 (.ZN (n_34_78), .A (n_35_79), .B (n_32_81), .C1 (n_31_80), .C2 (n_28_80) );
AOI211_X1 g_32_79 (.ZN (n_32_79), .A (n_33_80), .B (n_31_79), .C1 (n_33_79), .C2 (n_30_79) );
AOI211_X1 g_30_80 (.ZN (n_30_80), .A (n_34_78), .B (n_33_78), .C1 (n_32_81), .C2 (n_29_81) );
AOI211_X1 g_28_81 (.ZN (n_28_81), .A (n_32_79), .B (n_35_79), .C1 (n_31_79), .C2 (n_31_80) );
AOI211_X1 g_30_82 (.ZN (n_30_82), .A (n_30_80), .B (n_33_80), .C1 (n_33_78), .C2 (n_33_79) );
AOI211_X1 g_29_80 (.ZN (n_29_80), .A (n_28_81), .B (n_34_78), .C1 (n_35_79), .C2 (n_32_81) );
AOI211_X1 g_27_81 (.ZN (n_27_81), .A (n_30_82), .B (n_32_79), .C1 (n_33_80), .C2 (n_31_79) );
AOI211_X1 g_25_82 (.ZN (n_25_82), .A (n_29_80), .B (n_30_80), .C1 (n_34_78), .C2 (n_33_78) );
AOI211_X1 g_23_83 (.ZN (n_23_83), .A (n_27_81), .B (n_28_81), .C1 (n_32_79), .C2 (n_35_79) );
AOI211_X1 g_21_84 (.ZN (n_21_84), .A (n_25_82), .B (n_30_82), .C1 (n_30_80), .C2 (n_33_80) );
AOI211_X1 g_19_85 (.ZN (n_19_85), .A (n_23_83), .B (n_29_80), .C1 (n_28_81), .C2 (n_34_78) );
AOI211_X1 g_17_86 (.ZN (n_17_86), .A (n_21_84), .B (n_27_81), .C1 (n_30_82), .C2 (n_32_79) );
AOI211_X1 g_15_87 (.ZN (n_15_87), .A (n_19_85), .B (n_25_82), .C1 (n_29_80), .C2 (n_30_80) );
AOI211_X1 g_13_88 (.ZN (n_13_88), .A (n_17_86), .B (n_23_83), .C1 (n_27_81), .C2 (n_28_81) );
AOI211_X1 g_11_89 (.ZN (n_11_89), .A (n_15_87), .B (n_21_84), .C1 (n_25_82), .C2 (n_30_82) );
AOI211_X1 g_9_90 (.ZN (n_9_90), .A (n_13_88), .B (n_19_85), .C1 (n_23_83), .C2 (n_29_80) );
AOI211_X1 g_7_91 (.ZN (n_7_91), .A (n_11_89), .B (n_17_86), .C1 (n_21_84), .C2 (n_27_81) );
AOI211_X1 g_5_92 (.ZN (n_5_92), .A (n_9_90), .B (n_15_87), .C1 (n_19_85), .C2 (n_25_82) );
AOI211_X1 g_3_93 (.ZN (n_3_93), .A (n_7_91), .B (n_13_88), .C1 (n_17_86), .C2 (n_23_83) );
AOI211_X1 g_4_91 (.ZN (n_4_91), .A (n_5_92), .B (n_11_89), .C1 (n_15_87), .C2 (n_21_84) );
AOI211_X1 g_6_92 (.ZN (n_6_92), .A (n_3_93), .B (n_9_90), .C1 (n_13_88), .C2 (n_19_85) );
AOI211_X1 g_5_94 (.ZN (n_5_94), .A (n_4_91), .B (n_7_91), .C1 (n_11_89), .C2 (n_17_86) );
AOI211_X1 g_3_95 (.ZN (n_3_95), .A (n_6_92), .B (n_5_92), .C1 (n_9_90), .C2 (n_15_87) );
AOI211_X1 g_1_96 (.ZN (n_1_96), .A (n_5_94), .B (n_3_93), .C1 (n_7_91), .C2 (n_13_88) );
AOI211_X1 g_2_94 (.ZN (n_2_94), .A (n_3_95), .B (n_4_91), .C1 (n_5_92), .C2 (n_11_89) );
AOI211_X1 g_4_93 (.ZN (n_4_93), .A (n_1_96), .B (n_6_92), .C1 (n_3_93), .C2 (n_9_90) );
AOI211_X1 g_5_91 (.ZN (n_5_91), .A (n_2_94), .B (n_5_94), .C1 (n_4_91), .C2 (n_7_91) );
AOI211_X1 g_3_92 (.ZN (n_3_92), .A (n_4_93), .B (n_3_95), .C1 (n_6_92), .C2 (n_5_92) );
AOI211_X1 g_4_94 (.ZN (n_4_94), .A (n_5_91), .B (n_1_96), .C1 (n_5_94), .C2 (n_3_93) );
AOI211_X1 g_6_93 (.ZN (n_6_93), .A (n_3_92), .B (n_2_94), .C1 (n_3_95), .C2 (n_4_91) );
AOI211_X1 g_8_92 (.ZN (n_8_92), .A (n_4_94), .B (n_4_93), .C1 (n_1_96), .C2 (n_6_92) );
AOI211_X1 g_6_91 (.ZN (n_6_91), .A (n_6_93), .B (n_5_91), .C1 (n_2_94), .C2 (n_5_94) );
AOI211_X1 g_8_90 (.ZN (n_8_90), .A (n_8_92), .B (n_3_92), .C1 (n_4_93), .C2 (n_3_95) );
AOI211_X1 g_10_89 (.ZN (n_10_89), .A (n_6_91), .B (n_4_94), .C1 (n_5_91), .C2 (n_1_96) );
AOI211_X1 g_12_88 (.ZN (n_12_88), .A (n_8_90), .B (n_6_93), .C1 (n_3_92), .C2 (n_2_94) );
AOI211_X1 g_14_87 (.ZN (n_14_87), .A (n_10_89), .B (n_8_92), .C1 (n_4_94), .C2 (n_4_93) );
AOI211_X1 g_13_89 (.ZN (n_13_89), .A (n_12_88), .B (n_6_91), .C1 (n_6_93), .C2 (n_5_91) );
AOI211_X1 g_15_88 (.ZN (n_15_88), .A (n_14_87), .B (n_8_90), .C1 (n_8_92), .C2 (n_3_92) );
AOI211_X1 g_17_87 (.ZN (n_17_87), .A (n_13_89), .B (n_10_89), .C1 (n_6_91), .C2 (n_4_94) );
AOI211_X1 g_19_86 (.ZN (n_19_86), .A (n_15_88), .B (n_12_88), .C1 (n_8_90), .C2 (n_6_93) );
AOI211_X1 g_21_85 (.ZN (n_21_85), .A (n_17_87), .B (n_14_87), .C1 (n_10_89), .C2 (n_8_92) );
AOI211_X1 g_22_83 (.ZN (n_22_83), .A (n_19_86), .B (n_13_89), .C1 (n_12_88), .C2 (n_6_91) );
AOI211_X1 g_24_82 (.ZN (n_24_82), .A (n_21_85), .B (n_15_88), .C1 (n_14_87), .C2 (n_8_90) );
AOI211_X1 g_26_81 (.ZN (n_26_81), .A (n_22_83), .B (n_17_87), .C1 (n_13_89), .C2 (n_10_89) );
AOI211_X1 g_25_83 (.ZN (n_25_83), .A (n_24_82), .B (n_19_86), .C1 (n_15_88), .C2 (n_12_88) );
AOI211_X1 g_27_82 (.ZN (n_27_82), .A (n_26_81), .B (n_21_85), .C1 (n_17_87), .C2 (n_14_87) );
AOI211_X1 g_26_84 (.ZN (n_26_84), .A (n_25_83), .B (n_22_83), .C1 (n_19_86), .C2 (n_13_89) );
AOI211_X1 g_28_83 (.ZN (n_28_83), .A (n_27_82), .B (n_24_82), .C1 (n_21_85), .C2 (n_15_88) );
AOI211_X1 g_27_85 (.ZN (n_27_85), .A (n_26_84), .B (n_26_81), .C1 (n_22_83), .C2 (n_17_87) );
AOI211_X1 g_26_83 (.ZN (n_26_83), .A (n_28_83), .B (n_25_83), .C1 (n_24_82), .C2 (n_19_86) );
AOI211_X1 g_28_82 (.ZN (n_28_82), .A (n_27_85), .B (n_27_82), .C1 (n_26_81), .C2 (n_21_85) );
AOI211_X1 g_30_81 (.ZN (n_30_81), .A (n_26_83), .B (n_26_84), .C1 (n_25_83), .C2 (n_22_83) );
AOI211_X1 g_32_80 (.ZN (n_32_80), .A (n_28_82), .B (n_28_83), .C1 (n_27_82), .C2 (n_24_82) );
AOI211_X1 g_34_79 (.ZN (n_34_79), .A (n_30_81), .B (n_27_85), .C1 (n_26_84), .C2 (n_26_81) );
AOI211_X1 g_36_78 (.ZN (n_36_78), .A (n_32_80), .B (n_26_83), .C1 (n_28_83), .C2 (n_25_83) );
AOI211_X1 g_38_77 (.ZN (n_38_77), .A (n_34_79), .B (n_28_82), .C1 (n_27_85), .C2 (n_27_82) );
AOI211_X1 g_40_76 (.ZN (n_40_76), .A (n_36_78), .B (n_30_81), .C1 (n_26_83), .C2 (n_26_84) );
AOI211_X1 g_42_75 (.ZN (n_42_75), .A (n_38_77), .B (n_32_80), .C1 (n_28_82), .C2 (n_28_83) );
AOI211_X1 g_44_74 (.ZN (n_44_74), .A (n_40_76), .B (n_34_79), .C1 (n_30_81), .C2 (n_27_85) );
AOI211_X1 g_46_73 (.ZN (n_46_73), .A (n_42_75), .B (n_36_78), .C1 (n_32_80), .C2 (n_26_83) );
AOI211_X1 g_48_72 (.ZN (n_48_72), .A (n_44_74), .B (n_38_77), .C1 (n_34_79), .C2 (n_28_82) );
AOI211_X1 g_50_71 (.ZN (n_50_71), .A (n_46_73), .B (n_40_76), .C1 (n_36_78), .C2 (n_30_81) );
AOI211_X1 g_52_70 (.ZN (n_52_70), .A (n_48_72), .B (n_42_75), .C1 (n_38_77), .C2 (n_32_80) );
AOI211_X1 g_54_69 (.ZN (n_54_69), .A (n_50_71), .B (n_44_74), .C1 (n_40_76), .C2 (n_34_79) );
AOI211_X1 g_56_68 (.ZN (n_56_68), .A (n_52_70), .B (n_46_73), .C1 (n_42_75), .C2 (n_36_78) );
AOI211_X1 g_55_70 (.ZN (n_55_70), .A (n_54_69), .B (n_48_72), .C1 (n_44_74), .C2 (n_38_77) );
AOI211_X1 g_57_69 (.ZN (n_57_69), .A (n_56_68), .B (n_50_71), .C1 (n_46_73), .C2 (n_40_76) );
AOI211_X1 g_59_68 (.ZN (n_59_68), .A (n_55_70), .B (n_52_70), .C1 (n_48_72), .C2 (n_42_75) );
AOI211_X1 g_61_67 (.ZN (n_61_67), .A (n_57_69), .B (n_54_69), .C1 (n_50_71), .C2 (n_44_74) );
AOI211_X1 g_60_65 (.ZN (n_60_65), .A (n_59_68), .B (n_56_68), .C1 (n_52_70), .C2 (n_46_73) );
AOI211_X1 g_62_64 (.ZN (n_62_64), .A (n_61_67), .B (n_55_70), .C1 (n_54_69), .C2 (n_48_72) );
AOI211_X1 g_64_63 (.ZN (n_64_63), .A (n_60_65), .B (n_57_69), .C1 (n_56_68), .C2 (n_50_71) );
AOI211_X1 g_66_62 (.ZN (n_66_62), .A (n_62_64), .B (n_59_68), .C1 (n_55_70), .C2 (n_52_70) );
AOI211_X1 g_68_61 (.ZN (n_68_61), .A (n_64_63), .B (n_61_67), .C1 (n_57_69), .C2 (n_54_69) );
AOI211_X1 g_70_60 (.ZN (n_70_60), .A (n_66_62), .B (n_60_65), .C1 (n_59_68), .C2 (n_56_68) );
AOI211_X1 g_72_59 (.ZN (n_72_59), .A (n_68_61), .B (n_62_64), .C1 (n_61_67), .C2 (n_55_70) );
AOI211_X1 g_74_58 (.ZN (n_74_58), .A (n_70_60), .B (n_64_63), .C1 (n_60_65), .C2 (n_57_69) );
AOI211_X1 g_76_57 (.ZN (n_76_57), .A (n_72_59), .B (n_66_62), .C1 (n_62_64), .C2 (n_59_68) );
AOI211_X1 g_78_56 (.ZN (n_78_56), .A (n_74_58), .B (n_68_61), .C1 (n_64_63), .C2 (n_61_67) );
AOI211_X1 g_80_55 (.ZN (n_80_55), .A (n_76_57), .B (n_70_60), .C1 (n_66_62), .C2 (n_60_65) );
AOI211_X1 g_82_54 (.ZN (n_82_54), .A (n_78_56), .B (n_72_59), .C1 (n_68_61), .C2 (n_62_64) );
AOI211_X1 g_84_53 (.ZN (n_84_53), .A (n_80_55), .B (n_74_58), .C1 (n_70_60), .C2 (n_64_63) );
AOI211_X1 g_86_52 (.ZN (n_86_52), .A (n_82_54), .B (n_76_57), .C1 (n_72_59), .C2 (n_66_62) );
AOI211_X1 g_88_51 (.ZN (n_88_51), .A (n_84_53), .B (n_78_56), .C1 (n_74_58), .C2 (n_68_61) );
AOI211_X1 g_89_53 (.ZN (n_89_53), .A (n_86_52), .B (n_80_55), .C1 (n_76_57), .C2 (n_70_60) );
AOI211_X1 g_87_54 (.ZN (n_87_54), .A (n_88_51), .B (n_82_54), .C1 (n_78_56), .C2 (n_72_59) );
AOI211_X1 g_85_55 (.ZN (n_85_55), .A (n_89_53), .B (n_84_53), .C1 (n_80_55), .C2 (n_74_58) );
AOI211_X1 g_83_56 (.ZN (n_83_56), .A (n_87_54), .B (n_86_52), .C1 (n_82_54), .C2 (n_76_57) );
AOI211_X1 g_81_57 (.ZN (n_81_57), .A (n_85_55), .B (n_88_51), .C1 (n_84_53), .C2 (n_78_56) );
AOI211_X1 g_79_58 (.ZN (n_79_58), .A (n_83_56), .B (n_89_53), .C1 (n_86_52), .C2 (n_80_55) );
AOI211_X1 g_77_59 (.ZN (n_77_59), .A (n_81_57), .B (n_87_54), .C1 (n_88_51), .C2 (n_82_54) );
AOI211_X1 g_75_60 (.ZN (n_75_60), .A (n_79_58), .B (n_85_55), .C1 (n_89_53), .C2 (n_84_53) );
AOI211_X1 g_73_61 (.ZN (n_73_61), .A (n_77_59), .B (n_83_56), .C1 (n_87_54), .C2 (n_86_52) );
AOI211_X1 g_71_62 (.ZN (n_71_62), .A (n_75_60), .B (n_81_57), .C1 (n_85_55), .C2 (n_88_51) );
AOI211_X1 g_69_63 (.ZN (n_69_63), .A (n_73_61), .B (n_79_58), .C1 (n_83_56), .C2 (n_89_53) );
AOI211_X1 g_67_64 (.ZN (n_67_64), .A (n_71_62), .B (n_77_59), .C1 (n_81_57), .C2 (n_87_54) );
AOI211_X1 g_65_65 (.ZN (n_65_65), .A (n_69_63), .B (n_75_60), .C1 (n_79_58), .C2 (n_85_55) );
AOI211_X1 g_63_66 (.ZN (n_63_66), .A (n_67_64), .B (n_73_61), .C1 (n_77_59), .C2 (n_83_56) );
AOI211_X1 g_62_68 (.ZN (n_62_68), .A (n_65_65), .B (n_71_62), .C1 (n_75_60), .C2 (n_81_57) );
AOI211_X1 g_61_66 (.ZN (n_61_66), .A (n_63_66), .B (n_69_63), .C1 (n_73_61), .C2 (n_79_58) );
AOI211_X1 g_63_65 (.ZN (n_63_65), .A (n_62_68), .B (n_67_64), .C1 (n_71_62), .C2 (n_77_59) );
AOI211_X1 g_65_64 (.ZN (n_65_64), .A (n_61_66), .B (n_65_65), .C1 (n_69_63), .C2 (n_75_60) );
AOI211_X1 g_67_63 (.ZN (n_67_63), .A (n_63_65), .B (n_63_66), .C1 (n_67_64), .C2 (n_73_61) );
AOI211_X1 g_69_62 (.ZN (n_69_62), .A (n_65_64), .B (n_62_68), .C1 (n_65_65), .C2 (n_71_62) );
AOI211_X1 g_71_61 (.ZN (n_71_61), .A (n_67_63), .B (n_61_66), .C1 (n_63_66), .C2 (n_69_63) );
AOI211_X1 g_73_60 (.ZN (n_73_60), .A (n_69_62), .B (n_63_65), .C1 (n_62_68), .C2 (n_67_64) );
AOI211_X1 g_75_59 (.ZN (n_75_59), .A (n_71_61), .B (n_65_64), .C1 (n_61_66), .C2 (n_65_65) );
AOI211_X1 g_77_58 (.ZN (n_77_58), .A (n_73_60), .B (n_67_63), .C1 (n_63_65), .C2 (n_63_66) );
AOI211_X1 g_79_57 (.ZN (n_79_57), .A (n_75_59), .B (n_69_62), .C1 (n_65_64), .C2 (n_62_68) );
AOI211_X1 g_81_56 (.ZN (n_81_56), .A (n_77_58), .B (n_71_61), .C1 (n_67_63), .C2 (n_61_66) );
AOI211_X1 g_83_55 (.ZN (n_83_55), .A (n_79_57), .B (n_73_60), .C1 (n_69_62), .C2 (n_63_65) );
AOI211_X1 g_85_54 (.ZN (n_85_54), .A (n_81_56), .B (n_75_59), .C1 (n_71_61), .C2 (n_65_64) );
AOI211_X1 g_87_53 (.ZN (n_87_53), .A (n_83_55), .B (n_77_58), .C1 (n_73_60), .C2 (n_67_63) );
AOI211_X1 g_89_52 (.ZN (n_89_52), .A (n_85_54), .B (n_79_57), .C1 (n_75_59), .C2 (n_69_62) );
AOI211_X1 g_91_51 (.ZN (n_91_51), .A (n_87_53), .B (n_81_56), .C1 (n_77_58), .C2 (n_71_61) );
AOI211_X1 g_93_50 (.ZN (n_93_50), .A (n_89_52), .B (n_83_55), .C1 (n_79_57), .C2 (n_73_60) );
AOI211_X1 g_95_49 (.ZN (n_95_49), .A (n_91_51), .B (n_85_54), .C1 (n_81_56), .C2 (n_75_59) );
AOI211_X1 g_97_48 (.ZN (n_97_48), .A (n_93_50), .B (n_87_53), .C1 (n_83_55), .C2 (n_77_58) );
AOI211_X1 g_99_47 (.ZN (n_99_47), .A (n_95_49), .B (n_89_52), .C1 (n_85_54), .C2 (n_79_57) );
AOI211_X1 g_101_46 (.ZN (n_101_46), .A (n_97_48), .B (n_91_51), .C1 (n_87_53), .C2 (n_81_56) );
AOI211_X1 g_103_45 (.ZN (n_103_45), .A (n_99_47), .B (n_93_50), .C1 (n_89_52), .C2 (n_83_55) );
AOI211_X1 g_105_44 (.ZN (n_105_44), .A (n_101_46), .B (n_95_49), .C1 (n_91_51), .C2 (n_85_54) );
AOI211_X1 g_107_43 (.ZN (n_107_43), .A (n_103_45), .B (n_97_48), .C1 (n_93_50), .C2 (n_87_53) );
AOI211_X1 g_106_45 (.ZN (n_106_45), .A (n_105_44), .B (n_99_47), .C1 (n_95_49), .C2 (n_89_52) );
AOI211_X1 g_104_46 (.ZN (n_104_46), .A (n_107_43), .B (n_101_46), .C1 (n_97_48), .C2 (n_91_51) );
AOI211_X1 g_102_47 (.ZN (n_102_47), .A (n_106_45), .B (n_103_45), .C1 (n_99_47), .C2 (n_93_50) );
AOI211_X1 g_100_48 (.ZN (n_100_48), .A (n_104_46), .B (n_105_44), .C1 (n_101_46), .C2 (n_95_49) );
AOI211_X1 g_98_49 (.ZN (n_98_49), .A (n_102_47), .B (n_107_43), .C1 (n_103_45), .C2 (n_97_48) );
AOI211_X1 g_96_50 (.ZN (n_96_50), .A (n_100_48), .B (n_106_45), .C1 (n_105_44), .C2 (n_99_47) );
AOI211_X1 g_94_51 (.ZN (n_94_51), .A (n_98_49), .B (n_104_46), .C1 (n_107_43), .C2 (n_101_46) );
AOI211_X1 g_92_52 (.ZN (n_92_52), .A (n_96_50), .B (n_102_47), .C1 (n_106_45), .C2 (n_103_45) );
AOI211_X1 g_90_53 (.ZN (n_90_53), .A (n_94_51), .B (n_100_48), .C1 (n_104_46), .C2 (n_105_44) );
AOI211_X1 g_88_54 (.ZN (n_88_54), .A (n_92_52), .B (n_98_49), .C1 (n_102_47), .C2 (n_107_43) );
AOI211_X1 g_86_55 (.ZN (n_86_55), .A (n_90_53), .B (n_96_50), .C1 (n_100_48), .C2 (n_106_45) );
AOI211_X1 g_84_56 (.ZN (n_84_56), .A (n_88_54), .B (n_94_51), .C1 (n_98_49), .C2 (n_104_46) );
AOI211_X1 g_82_57 (.ZN (n_82_57), .A (n_86_55), .B (n_92_52), .C1 (n_96_50), .C2 (n_102_47) );
AOI211_X1 g_80_58 (.ZN (n_80_58), .A (n_84_56), .B (n_90_53), .C1 (n_94_51), .C2 (n_100_48) );
AOI211_X1 g_78_59 (.ZN (n_78_59), .A (n_82_57), .B (n_88_54), .C1 (n_92_52), .C2 (n_98_49) );
AOI211_X1 g_76_60 (.ZN (n_76_60), .A (n_80_58), .B (n_86_55), .C1 (n_90_53), .C2 (n_96_50) );
AOI211_X1 g_74_61 (.ZN (n_74_61), .A (n_78_59), .B (n_84_56), .C1 (n_88_54), .C2 (n_94_51) );
AOI211_X1 g_72_62 (.ZN (n_72_62), .A (n_76_60), .B (n_82_57), .C1 (n_86_55), .C2 (n_92_52) );
AOI211_X1 g_70_63 (.ZN (n_70_63), .A (n_74_61), .B (n_80_58), .C1 (n_84_56), .C2 (n_90_53) );
AOI211_X1 g_68_64 (.ZN (n_68_64), .A (n_72_62), .B (n_78_59), .C1 (n_82_57), .C2 (n_88_54) );
AOI211_X1 g_66_65 (.ZN (n_66_65), .A (n_70_63), .B (n_76_60), .C1 (n_80_58), .C2 (n_86_55) );
AOI211_X1 g_64_66 (.ZN (n_64_66), .A (n_68_64), .B (n_74_61), .C1 (n_78_59), .C2 (n_84_56) );
AOI211_X1 g_62_67 (.ZN (n_62_67), .A (n_66_65), .B (n_72_62), .C1 (n_76_60), .C2 (n_82_57) );
AOI211_X1 g_60_68 (.ZN (n_60_68), .A (n_64_66), .B (n_70_63), .C1 (n_74_61), .C2 (n_80_58) );
AOI211_X1 g_58_69 (.ZN (n_58_69), .A (n_62_67), .B (n_68_64), .C1 (n_72_62), .C2 (n_78_59) );
AOI211_X1 g_59_67 (.ZN (n_59_67), .A (n_60_68), .B (n_66_65), .C1 (n_70_63), .C2 (n_76_60) );
AOI211_X1 g_57_68 (.ZN (n_57_68), .A (n_58_69), .B (n_64_66), .C1 (n_68_64), .C2 (n_74_61) );
AOI211_X1 g_55_69 (.ZN (n_55_69), .A (n_59_67), .B (n_62_67), .C1 (n_66_65), .C2 (n_72_62) );
AOI211_X1 g_53_70 (.ZN (n_53_70), .A (n_57_68), .B (n_60_68), .C1 (n_64_66), .C2 (n_70_63) );
AOI211_X1 g_51_71 (.ZN (n_51_71), .A (n_55_69), .B (n_58_69), .C1 (n_62_67), .C2 (n_68_64) );
AOI211_X1 g_49_72 (.ZN (n_49_72), .A (n_53_70), .B (n_59_67), .C1 (n_60_68), .C2 (n_66_65) );
AOI211_X1 g_47_73 (.ZN (n_47_73), .A (n_51_71), .B (n_57_68), .C1 (n_58_69), .C2 (n_64_66) );
AOI211_X1 g_45_74 (.ZN (n_45_74), .A (n_49_72), .B (n_55_69), .C1 (n_59_67), .C2 (n_62_67) );
AOI211_X1 g_43_75 (.ZN (n_43_75), .A (n_47_73), .B (n_53_70), .C1 (n_57_68), .C2 (n_60_68) );
AOI211_X1 g_41_76 (.ZN (n_41_76), .A (n_45_74), .B (n_51_71), .C1 (n_55_69), .C2 (n_58_69) );
AOI211_X1 g_39_77 (.ZN (n_39_77), .A (n_43_75), .B (n_49_72), .C1 (n_53_70), .C2 (n_59_67) );
AOI211_X1 g_38_79 (.ZN (n_38_79), .A (n_41_76), .B (n_47_73), .C1 (n_51_71), .C2 (n_57_68) );
AOI211_X1 g_40_78 (.ZN (n_40_78), .A (n_39_77), .B (n_45_74), .C1 (n_49_72), .C2 (n_55_69) );
AOI211_X1 g_42_77 (.ZN (n_42_77), .A (n_38_79), .B (n_43_75), .C1 (n_47_73), .C2 (n_53_70) );
AOI211_X1 g_44_76 (.ZN (n_44_76), .A (n_40_78), .B (n_41_76), .C1 (n_45_74), .C2 (n_51_71) );
AOI211_X1 g_46_75 (.ZN (n_46_75), .A (n_42_77), .B (n_39_77), .C1 (n_43_75), .C2 (n_49_72) );
AOI211_X1 g_48_74 (.ZN (n_48_74), .A (n_44_76), .B (n_38_79), .C1 (n_41_76), .C2 (n_47_73) );
AOI211_X1 g_50_73 (.ZN (n_50_73), .A (n_46_75), .B (n_40_78), .C1 (n_39_77), .C2 (n_45_74) );
AOI211_X1 g_52_72 (.ZN (n_52_72), .A (n_48_74), .B (n_42_77), .C1 (n_38_79), .C2 (n_43_75) );
AOI211_X1 g_54_71 (.ZN (n_54_71), .A (n_50_73), .B (n_44_76), .C1 (n_40_78), .C2 (n_41_76) );
AOI211_X1 g_56_70 (.ZN (n_56_70), .A (n_52_72), .B (n_46_75), .C1 (n_42_77), .C2 (n_39_77) );
AOI211_X1 g_58_71 (.ZN (n_58_71), .A (n_54_71), .B (n_48_74), .C1 (n_44_76), .C2 (n_38_79) );
AOI211_X1 g_60_70 (.ZN (n_60_70), .A (n_56_70), .B (n_50_73), .C1 (n_46_75), .C2 (n_40_78) );
AOI211_X1 g_62_69 (.ZN (n_62_69), .A (n_58_71), .B (n_52_72), .C1 (n_48_74), .C2 (n_42_77) );
AOI211_X1 g_64_68 (.ZN (n_64_68), .A (n_60_70), .B (n_54_71), .C1 (n_50_73), .C2 (n_44_76) );
AOI211_X1 g_66_67 (.ZN (n_66_67), .A (n_62_69), .B (n_56_70), .C1 (n_52_72), .C2 (n_46_75) );
AOI211_X1 g_68_66 (.ZN (n_68_66), .A (n_64_68), .B (n_58_71), .C1 (n_54_71), .C2 (n_48_74) );
AOI211_X1 g_70_65 (.ZN (n_70_65), .A (n_66_67), .B (n_60_70), .C1 (n_56_70), .C2 (n_50_73) );
AOI211_X1 g_72_64 (.ZN (n_72_64), .A (n_68_66), .B (n_62_69), .C1 (n_58_71), .C2 (n_52_72) );
AOI211_X1 g_74_63 (.ZN (n_74_63), .A (n_70_65), .B (n_64_68), .C1 (n_60_70), .C2 (n_54_71) );
AOI211_X1 g_76_62 (.ZN (n_76_62), .A (n_72_64), .B (n_66_67), .C1 (n_62_69), .C2 (n_56_70) );
AOI211_X1 g_78_61 (.ZN (n_78_61), .A (n_74_63), .B (n_68_66), .C1 (n_64_68), .C2 (n_58_71) );
AOI211_X1 g_80_60 (.ZN (n_80_60), .A (n_76_62), .B (n_70_65), .C1 (n_66_67), .C2 (n_60_70) );
AOI211_X1 g_82_59 (.ZN (n_82_59), .A (n_78_61), .B (n_72_64), .C1 (n_68_66), .C2 (n_62_69) );
AOI211_X1 g_84_58 (.ZN (n_84_58), .A (n_80_60), .B (n_74_63), .C1 (n_70_65), .C2 (n_64_68) );
AOI211_X1 g_86_57 (.ZN (n_86_57), .A (n_82_59), .B (n_76_62), .C1 (n_72_64), .C2 (n_66_67) );
AOI211_X1 g_88_56 (.ZN (n_88_56), .A (n_84_58), .B (n_78_61), .C1 (n_74_63), .C2 (n_68_66) );
AOI211_X1 g_90_55 (.ZN (n_90_55), .A (n_86_57), .B (n_80_60), .C1 (n_76_62), .C2 (n_70_65) );
AOI211_X1 g_92_54 (.ZN (n_92_54), .A (n_88_56), .B (n_82_59), .C1 (n_78_61), .C2 (n_72_64) );
AOI211_X1 g_93_52 (.ZN (n_93_52), .A (n_90_55), .B (n_84_58), .C1 (n_80_60), .C2 (n_74_63) );
AOI211_X1 g_94_50 (.ZN (n_94_50), .A (n_92_54), .B (n_86_57), .C1 (n_82_59), .C2 (n_76_62) );
AOI211_X1 g_96_49 (.ZN (n_96_49), .A (n_93_52), .B (n_88_56), .C1 (n_84_58), .C2 (n_78_61) );
AOI211_X1 g_98_48 (.ZN (n_98_48), .A (n_94_50), .B (n_90_55), .C1 (n_86_57), .C2 (n_80_60) );
AOI211_X1 g_100_47 (.ZN (n_100_47), .A (n_96_49), .B (n_92_54), .C1 (n_88_56), .C2 (n_82_59) );
AOI211_X1 g_102_46 (.ZN (n_102_46), .A (n_98_48), .B (n_93_52), .C1 (n_90_55), .C2 (n_84_58) );
AOI211_X1 g_104_45 (.ZN (n_104_45), .A (n_100_47), .B (n_94_50), .C1 (n_92_54), .C2 (n_86_57) );
AOI211_X1 g_106_44 (.ZN (n_106_44), .A (n_102_46), .B (n_96_49), .C1 (n_93_52), .C2 (n_88_56) );
AOI211_X1 g_108_43 (.ZN (n_108_43), .A (n_104_45), .B (n_98_48), .C1 (n_94_50), .C2 (n_90_55) );
AOI211_X1 g_110_42 (.ZN (n_110_42), .A (n_106_44), .B (n_100_47), .C1 (n_96_49), .C2 (n_92_54) );
AOI211_X1 g_109_40 (.ZN (n_109_40), .A (n_108_43), .B (n_102_46), .C1 (n_98_48), .C2 (n_93_52) );
AOI211_X1 g_111_39 (.ZN (n_111_39), .A (n_110_42), .B (n_104_45), .C1 (n_100_47), .C2 (n_94_50) );
AOI211_X1 g_113_38 (.ZN (n_113_38), .A (n_109_40), .B (n_106_44), .C1 (n_102_46), .C2 (n_96_49) );
AOI211_X1 g_115_37 (.ZN (n_115_37), .A (n_111_39), .B (n_108_43), .C1 (n_104_45), .C2 (n_98_48) );
AOI211_X1 g_117_36 (.ZN (n_117_36), .A (n_113_38), .B (n_110_42), .C1 (n_106_44), .C2 (n_100_47) );
AOI211_X1 g_119_37 (.ZN (n_119_37), .A (n_115_37), .B (n_109_40), .C1 (n_108_43), .C2 (n_102_46) );
AOI211_X1 g_117_38 (.ZN (n_117_38), .A (n_117_36), .B (n_111_39), .C1 (n_110_42), .C2 (n_104_45) );
AOI211_X1 g_115_39 (.ZN (n_115_39), .A (n_119_37), .B (n_113_38), .C1 (n_109_40), .C2 (n_106_44) );
AOI211_X1 g_113_40 (.ZN (n_113_40), .A (n_117_38), .B (n_115_37), .C1 (n_111_39), .C2 (n_108_43) );
AOI211_X1 g_111_41 (.ZN (n_111_41), .A (n_115_39), .B (n_117_36), .C1 (n_113_38), .C2 (n_110_42) );
AOI211_X1 g_110_43 (.ZN (n_110_43), .A (n_113_40), .B (n_119_37), .C1 (n_115_37), .C2 (n_109_40) );
AOI211_X1 g_108_42 (.ZN (n_108_42), .A (n_111_41), .B (n_117_38), .C1 (n_117_36), .C2 (n_111_39) );
AOI211_X1 g_106_43 (.ZN (n_106_43), .A (n_110_43), .B (n_115_39), .C1 (n_119_37), .C2 (n_113_38) );
AOI211_X1 g_108_44 (.ZN (n_108_44), .A (n_108_42), .B (n_113_40), .C1 (n_117_38), .C2 (n_115_37) );
AOI211_X1 g_107_46 (.ZN (n_107_46), .A (n_106_43), .B (n_111_41), .C1 (n_115_39), .C2 (n_117_36) );
AOI211_X1 g_105_45 (.ZN (n_105_45), .A (n_108_44), .B (n_110_43), .C1 (n_113_40), .C2 (n_119_37) );
AOI211_X1 g_107_44 (.ZN (n_107_44), .A (n_107_46), .B (n_108_42), .C1 (n_111_41), .C2 (n_117_38) );
AOI211_X1 g_109_45 (.ZN (n_109_45), .A (n_105_45), .B (n_106_43), .C1 (n_110_43), .C2 (n_115_39) );
AOI211_X1 g_111_44 (.ZN (n_111_44), .A (n_107_44), .B (n_108_44), .C1 (n_108_42), .C2 (n_113_40) );
AOI211_X1 g_112_42 (.ZN (n_112_42), .A (n_109_45), .B (n_107_46), .C1 (n_106_43), .C2 (n_111_41) );
AOI211_X1 g_110_41 (.ZN (n_110_41), .A (n_111_44), .B (n_105_45), .C1 (n_108_44), .C2 (n_110_43) );
AOI211_X1 g_109_43 (.ZN (n_109_43), .A (n_112_42), .B (n_107_44), .C1 (n_107_46), .C2 (n_108_42) );
AOI211_X1 g_111_42 (.ZN (n_111_42), .A (n_110_41), .B (n_109_45), .C1 (n_105_45), .C2 (n_106_43) );
AOI211_X1 g_112_40 (.ZN (n_112_40), .A (n_109_43), .B (n_111_44), .C1 (n_107_44), .C2 (n_108_44) );
AOI211_X1 g_114_39 (.ZN (n_114_39), .A (n_111_42), .B (n_112_42), .C1 (n_109_45), .C2 (n_107_46) );
AOI211_X1 g_116_38 (.ZN (n_116_38), .A (n_112_40), .B (n_110_41), .C1 (n_111_44), .C2 (n_105_45) );
AOI211_X1 g_118_37 (.ZN (n_118_37), .A (n_114_39), .B (n_109_43), .C1 (n_112_42), .C2 (n_107_44) );
AOI211_X1 g_120_36 (.ZN (n_120_36), .A (n_116_38), .B (n_111_42), .C1 (n_110_41), .C2 (n_109_45) );
AOI211_X1 g_122_35 (.ZN (n_122_35), .A (n_118_37), .B (n_112_40), .C1 (n_109_43), .C2 (n_111_44) );
AOI211_X1 g_124_34 (.ZN (n_124_34), .A (n_120_36), .B (n_114_39), .C1 (n_111_42), .C2 (n_112_42) );
AOI211_X1 g_123_36 (.ZN (n_123_36), .A (n_122_35), .B (n_116_38), .C1 (n_112_40), .C2 (n_110_41) );
AOI211_X1 g_125_35 (.ZN (n_125_35), .A (n_124_34), .B (n_118_37), .C1 (n_114_39), .C2 (n_109_43) );
AOI211_X1 g_127_34 (.ZN (n_127_34), .A (n_123_36), .B (n_120_36), .C1 (n_116_38), .C2 (n_111_42) );
AOI211_X1 g_129_33 (.ZN (n_129_33), .A (n_125_35), .B (n_122_35), .C1 (n_118_37), .C2 (n_112_40) );
AOI211_X1 g_131_32 (.ZN (n_131_32), .A (n_127_34), .B (n_124_34), .C1 (n_120_36), .C2 (n_114_39) );
AOI211_X1 g_133_31 (.ZN (n_133_31), .A (n_129_33), .B (n_123_36), .C1 (n_122_35), .C2 (n_116_38) );
AOI211_X1 g_132_33 (.ZN (n_132_33), .A (n_131_32), .B (n_125_35), .C1 (n_124_34), .C2 (n_118_37) );
AOI211_X1 g_130_34 (.ZN (n_130_34), .A (n_133_31), .B (n_127_34), .C1 (n_123_36), .C2 (n_120_36) );
AOI211_X1 g_128_33 (.ZN (n_128_33), .A (n_132_33), .B (n_129_33), .C1 (n_125_35), .C2 (n_122_35) );
AOI211_X1 g_126_34 (.ZN (n_126_34), .A (n_130_34), .B (n_131_32), .C1 (n_127_34), .C2 (n_124_34) );
AOI211_X1 g_124_35 (.ZN (n_124_35), .A (n_128_33), .B (n_133_31), .C1 (n_129_33), .C2 (n_123_36) );
AOI211_X1 g_122_36 (.ZN (n_122_36), .A (n_126_34), .B (n_132_33), .C1 (n_131_32), .C2 (n_125_35) );
AOI211_X1 g_120_37 (.ZN (n_120_37), .A (n_124_35), .B (n_130_34), .C1 (n_133_31), .C2 (n_127_34) );
AOI211_X1 g_118_38 (.ZN (n_118_38), .A (n_122_36), .B (n_128_33), .C1 (n_132_33), .C2 (n_129_33) );
AOI211_X1 g_116_39 (.ZN (n_116_39), .A (n_120_37), .B (n_126_34), .C1 (n_130_34), .C2 (n_131_32) );
AOI211_X1 g_114_40 (.ZN (n_114_40), .A (n_118_38), .B (n_124_35), .C1 (n_128_33), .C2 (n_133_31) );
AOI211_X1 g_112_41 (.ZN (n_112_41), .A (n_116_39), .B (n_122_36), .C1 (n_126_34), .C2 (n_132_33) );
AOI211_X1 g_111_43 (.ZN (n_111_43), .A (n_114_40), .B (n_120_37), .C1 (n_124_35), .C2 (n_130_34) );
AOI211_X1 g_113_42 (.ZN (n_113_42), .A (n_112_41), .B (n_118_38), .C1 (n_122_36), .C2 (n_128_33) );
AOI211_X1 g_115_41 (.ZN (n_115_41), .A (n_111_43), .B (n_116_39), .C1 (n_120_37), .C2 (n_126_34) );
AOI211_X1 g_117_40 (.ZN (n_117_40), .A (n_113_42), .B (n_114_40), .C1 (n_118_38), .C2 (n_124_35) );
AOI211_X1 g_119_39 (.ZN (n_119_39), .A (n_115_41), .B (n_112_41), .C1 (n_116_39), .C2 (n_122_36) );
AOI211_X1 g_121_38 (.ZN (n_121_38), .A (n_117_40), .B (n_111_43), .C1 (n_114_40), .C2 (n_120_37) );
AOI211_X1 g_123_37 (.ZN (n_123_37), .A (n_119_39), .B (n_113_42), .C1 (n_112_41), .C2 (n_118_38) );
AOI211_X1 g_125_36 (.ZN (n_125_36), .A (n_121_38), .B (n_115_41), .C1 (n_111_43), .C2 (n_116_39) );
AOI211_X1 g_127_35 (.ZN (n_127_35), .A (n_123_37), .B (n_117_40), .C1 (n_113_42), .C2 (n_114_40) );
AOI211_X1 g_126_37 (.ZN (n_126_37), .A (n_125_36), .B (n_119_39), .C1 (n_115_41), .C2 (n_112_41) );
AOI211_X1 g_124_36 (.ZN (n_124_36), .A (n_127_35), .B (n_121_38), .C1 (n_117_40), .C2 (n_111_43) );
AOI211_X1 g_126_35 (.ZN (n_126_35), .A (n_126_37), .B (n_123_37), .C1 (n_119_39), .C2 (n_113_42) );
AOI211_X1 g_128_34 (.ZN (n_128_34), .A (n_124_36), .B (n_125_36), .C1 (n_121_38), .C2 (n_115_41) );
AOI211_X1 g_130_33 (.ZN (n_130_33), .A (n_126_35), .B (n_127_35), .C1 (n_123_37), .C2 (n_117_40) );
AOI211_X1 g_132_32 (.ZN (n_132_32), .A (n_128_34), .B (n_126_37), .C1 (n_125_36), .C2 (n_119_39) );
AOI211_X1 g_134_31 (.ZN (n_134_31), .A (n_130_33), .B (n_124_36), .C1 (n_127_35), .C2 (n_121_38) );
AOI211_X1 g_136_30 (.ZN (n_136_30), .A (n_132_32), .B (n_126_35), .C1 (n_126_37), .C2 (n_123_37) );
AOI211_X1 g_138_29 (.ZN (n_138_29), .A (n_134_31), .B (n_128_34), .C1 (n_124_36), .C2 (n_125_36) );
AOI211_X1 g_140_28 (.ZN (n_140_28), .A (n_136_30), .B (n_130_33), .C1 (n_126_35), .C2 (n_127_35) );
AOI211_X1 g_139_30 (.ZN (n_139_30), .A (n_138_29), .B (n_132_32), .C1 (n_128_34), .C2 (n_126_37) );
AOI211_X1 g_137_31 (.ZN (n_137_31), .A (n_140_28), .B (n_134_31), .C1 (n_130_33), .C2 (n_124_36) );
AOI211_X1 g_135_32 (.ZN (n_135_32), .A (n_139_30), .B (n_136_30), .C1 (n_132_32), .C2 (n_126_35) );
AOI211_X1 g_133_33 (.ZN (n_133_33), .A (n_137_31), .B (n_138_29), .C1 (n_134_31), .C2 (n_128_34) );
AOI211_X1 g_131_34 (.ZN (n_131_34), .A (n_135_32), .B (n_140_28), .C1 (n_136_30), .C2 (n_130_33) );
AOI211_X1 g_129_35 (.ZN (n_129_35), .A (n_133_33), .B (n_139_30), .C1 (n_138_29), .C2 (n_132_32) );
AOI211_X1 g_127_36 (.ZN (n_127_36), .A (n_131_34), .B (n_137_31), .C1 (n_140_28), .C2 (n_134_31) );
AOI211_X1 g_125_37 (.ZN (n_125_37), .A (n_129_35), .B (n_135_32), .C1 (n_139_30), .C2 (n_136_30) );
AOI211_X1 g_123_38 (.ZN (n_123_38), .A (n_127_36), .B (n_133_33), .C1 (n_137_31), .C2 (n_138_29) );
AOI211_X1 g_121_37 (.ZN (n_121_37), .A (n_125_37), .B (n_131_34), .C1 (n_135_32), .C2 (n_140_28) );
AOI211_X1 g_119_38 (.ZN (n_119_38), .A (n_123_38), .B (n_129_35), .C1 (n_133_33), .C2 (n_139_30) );
AOI211_X1 g_117_39 (.ZN (n_117_39), .A (n_121_37), .B (n_127_36), .C1 (n_131_34), .C2 (n_137_31) );
AOI211_X1 g_115_40 (.ZN (n_115_40), .A (n_119_38), .B (n_125_37), .C1 (n_129_35), .C2 (n_135_32) );
AOI211_X1 g_113_41 (.ZN (n_113_41), .A (n_117_39), .B (n_123_38), .C1 (n_127_36), .C2 (n_133_33) );
AOI211_X1 g_112_43 (.ZN (n_112_43), .A (n_115_40), .B (n_121_37), .C1 (n_125_37), .C2 (n_131_34) );
AOI211_X1 g_114_42 (.ZN (n_114_42), .A (n_113_41), .B (n_119_38), .C1 (n_123_38), .C2 (n_129_35) );
AOI211_X1 g_116_41 (.ZN (n_116_41), .A (n_112_43), .B (n_117_39), .C1 (n_121_37), .C2 (n_127_36) );
AOI211_X1 g_118_40 (.ZN (n_118_40), .A (n_114_42), .B (n_115_40), .C1 (n_119_38), .C2 (n_125_37) );
AOI211_X1 g_120_39 (.ZN (n_120_39), .A (n_116_41), .B (n_113_41), .C1 (n_117_39), .C2 (n_123_38) );
AOI211_X1 g_122_38 (.ZN (n_122_38), .A (n_118_40), .B (n_112_43), .C1 (n_115_40), .C2 (n_121_37) );
AOI211_X1 g_124_37 (.ZN (n_124_37), .A (n_120_39), .B (n_114_42), .C1 (n_113_41), .C2 (n_119_38) );
AOI211_X1 g_126_36 (.ZN (n_126_36), .A (n_122_38), .B (n_116_41), .C1 (n_112_43), .C2 (n_117_39) );
AOI211_X1 g_128_35 (.ZN (n_128_35), .A (n_124_37), .B (n_118_40), .C1 (n_114_42), .C2 (n_115_40) );
AOI211_X1 g_127_37 (.ZN (n_127_37), .A (n_126_36), .B (n_120_39), .C1 (n_116_41), .C2 (n_113_41) );
AOI211_X1 g_129_36 (.ZN (n_129_36), .A (n_128_35), .B (n_122_38), .C1 (n_118_40), .C2 (n_112_43) );
AOI211_X1 g_131_35 (.ZN (n_131_35), .A (n_127_37), .B (n_124_37), .C1 (n_120_39), .C2 (n_114_42) );
AOI211_X1 g_133_34 (.ZN (n_133_34), .A (n_129_36), .B (n_126_36), .C1 (n_122_38), .C2 (n_116_41) );
AOI211_X1 g_135_33 (.ZN (n_135_33), .A (n_131_35), .B (n_128_35), .C1 (n_124_37), .C2 (n_118_40) );
AOI211_X1 g_137_32 (.ZN (n_137_32), .A (n_133_34), .B (n_127_37), .C1 (n_126_36), .C2 (n_120_39) );
AOI211_X1 g_139_31 (.ZN (n_139_31), .A (n_135_33), .B (n_129_36), .C1 (n_128_35), .C2 (n_122_38) );
AOI211_X1 g_141_30 (.ZN (n_141_30), .A (n_137_32), .B (n_131_35), .C1 (n_127_37), .C2 (n_124_37) );
AOI211_X1 g_143_29 (.ZN (n_143_29), .A (n_139_31), .B (n_133_34), .C1 (n_129_36), .C2 (n_126_36) );
AOI211_X1 g_145_28 (.ZN (n_145_28), .A (n_141_30), .B (n_135_33), .C1 (n_131_35), .C2 (n_128_35) );
AOI211_X1 g_147_29 (.ZN (n_147_29), .A (n_143_29), .B (n_137_32), .C1 (n_133_34), .C2 (n_127_37) );
AOI211_X1 g_145_30 (.ZN (n_145_30), .A (n_145_28), .B (n_139_31), .C1 (n_135_33), .C2 (n_129_36) );
AOI211_X1 g_143_31 (.ZN (n_143_31), .A (n_147_29), .B (n_141_30), .C1 (n_137_32), .C2 (n_131_35) );
AOI211_X1 g_141_32 (.ZN (n_141_32), .A (n_145_30), .B (n_143_29), .C1 (n_139_31), .C2 (n_133_34) );
AOI211_X1 g_140_30 (.ZN (n_140_30), .A (n_143_31), .B (n_145_28), .C1 (n_141_30), .C2 (n_135_33) );
AOI211_X1 g_138_31 (.ZN (n_138_31), .A (n_141_32), .B (n_147_29), .C1 (n_143_29), .C2 (n_137_32) );
AOI211_X1 g_136_32 (.ZN (n_136_32), .A (n_140_30), .B (n_145_30), .C1 (n_145_28), .C2 (n_139_31) );
AOI211_X1 g_134_33 (.ZN (n_134_33), .A (n_138_31), .B (n_143_31), .C1 (n_147_29), .C2 (n_141_30) );
AOI211_X1 g_132_34 (.ZN (n_132_34), .A (n_136_32), .B (n_141_32), .C1 (n_145_30), .C2 (n_143_29) );
AOI211_X1 g_130_35 (.ZN (n_130_35), .A (n_134_33), .B (n_140_30), .C1 (n_143_31), .C2 (n_145_28) );
AOI211_X1 g_128_36 (.ZN (n_128_36), .A (n_132_34), .B (n_138_31), .C1 (n_141_32), .C2 (n_147_29) );
AOI211_X1 g_127_38 (.ZN (n_127_38), .A (n_130_35), .B (n_136_32), .C1 (n_140_30), .C2 (n_145_30) );
AOI211_X1 g_129_37 (.ZN (n_129_37), .A (n_128_36), .B (n_134_33), .C1 (n_138_31), .C2 (n_143_31) );
AOI211_X1 g_131_36 (.ZN (n_131_36), .A (n_127_38), .B (n_132_34), .C1 (n_136_32), .C2 (n_141_32) );
AOI211_X1 g_133_35 (.ZN (n_133_35), .A (n_129_37), .B (n_130_35), .C1 (n_134_33), .C2 (n_140_30) );
AOI211_X1 g_135_34 (.ZN (n_135_34), .A (n_131_36), .B (n_128_36), .C1 (n_132_34), .C2 (n_138_31) );
AOI211_X1 g_137_33 (.ZN (n_137_33), .A (n_133_35), .B (n_127_38), .C1 (n_130_35), .C2 (n_136_32) );
AOI211_X1 g_139_32 (.ZN (n_139_32), .A (n_135_34), .B (n_129_37), .C1 (n_128_36), .C2 (n_134_33) );
AOI211_X1 g_141_31 (.ZN (n_141_31), .A (n_137_33), .B (n_131_36), .C1 (n_127_38), .C2 (n_132_34) );
AOI211_X1 g_143_32 (.ZN (n_143_32), .A (n_139_32), .B (n_133_35), .C1 (n_129_37), .C2 (n_130_35) );
AOI211_X1 g_144_30 (.ZN (n_144_30), .A (n_141_31), .B (n_135_34), .C1 (n_131_36), .C2 (n_128_36) );
AOI211_X1 g_146_31 (.ZN (n_146_31), .A (n_143_32), .B (n_137_33), .C1 (n_133_35), .C2 (n_127_38) );
AOI211_X1 g_144_32 (.ZN (n_144_32), .A (n_144_30), .B (n_139_32), .C1 (n_135_34), .C2 (n_129_37) );
AOI211_X1 g_142_31 (.ZN (n_142_31), .A (n_146_31), .B (n_141_31), .C1 (n_137_33), .C2 (n_131_36) );
AOI211_X1 g_140_32 (.ZN (n_140_32), .A (n_144_32), .B (n_143_32), .C1 (n_139_32), .C2 (n_133_35) );
AOI211_X1 g_138_33 (.ZN (n_138_33), .A (n_142_31), .B (n_144_30), .C1 (n_141_31), .C2 (n_135_34) );
AOI211_X1 g_136_34 (.ZN (n_136_34), .A (n_140_32), .B (n_146_31), .C1 (n_143_32), .C2 (n_137_33) );
AOI211_X1 g_134_35 (.ZN (n_134_35), .A (n_138_33), .B (n_144_32), .C1 (n_144_30), .C2 (n_139_32) );
AOI211_X1 g_132_36 (.ZN (n_132_36), .A (n_136_34), .B (n_142_31), .C1 (n_146_31), .C2 (n_141_31) );
AOI211_X1 g_130_37 (.ZN (n_130_37), .A (n_134_35), .B (n_140_32), .C1 (n_144_32), .C2 (n_143_32) );
AOI211_X1 g_128_38 (.ZN (n_128_38), .A (n_132_36), .B (n_138_33), .C1 (n_142_31), .C2 (n_144_30) );
AOI211_X1 g_126_39 (.ZN (n_126_39), .A (n_130_37), .B (n_136_34), .C1 (n_140_32), .C2 (n_146_31) );
AOI211_X1 g_124_38 (.ZN (n_124_38), .A (n_128_38), .B (n_134_35), .C1 (n_138_33), .C2 (n_144_32) );
AOI211_X1 g_122_37 (.ZN (n_122_37), .A (n_126_39), .B (n_132_36), .C1 (n_136_34), .C2 (n_142_31) );
AOI211_X1 g_120_38 (.ZN (n_120_38), .A (n_124_38), .B (n_130_37), .C1 (n_134_35), .C2 (n_140_32) );
AOI211_X1 g_118_39 (.ZN (n_118_39), .A (n_122_37), .B (n_128_38), .C1 (n_132_36), .C2 (n_138_33) );
AOI211_X1 g_116_40 (.ZN (n_116_40), .A (n_120_38), .B (n_126_39), .C1 (n_130_37), .C2 (n_136_34) );
AOI211_X1 g_114_41 (.ZN (n_114_41), .A (n_118_39), .B (n_124_38), .C1 (n_128_38), .C2 (n_134_35) );
AOI211_X1 g_113_43 (.ZN (n_113_43), .A (n_116_40), .B (n_122_37), .C1 (n_126_39), .C2 (n_132_36) );
AOI211_X1 g_115_42 (.ZN (n_115_42), .A (n_114_41), .B (n_120_38), .C1 (n_124_38), .C2 (n_130_37) );
AOI211_X1 g_117_41 (.ZN (n_117_41), .A (n_113_43), .B (n_118_39), .C1 (n_122_37), .C2 (n_128_38) );
AOI211_X1 g_119_40 (.ZN (n_119_40), .A (n_115_42), .B (n_116_40), .C1 (n_120_38), .C2 (n_126_39) );
AOI211_X1 g_121_39 (.ZN (n_121_39), .A (n_117_41), .B (n_114_41), .C1 (n_118_39), .C2 (n_124_38) );
AOI211_X1 g_120_41 (.ZN (n_120_41), .A (n_119_40), .B (n_113_43), .C1 (n_116_40), .C2 (n_122_37) );
AOI211_X1 g_122_40 (.ZN (n_122_40), .A (n_121_39), .B (n_115_42), .C1 (n_114_41), .C2 (n_120_38) );
AOI211_X1 g_124_39 (.ZN (n_124_39), .A (n_120_41), .B (n_117_41), .C1 (n_113_43), .C2 (n_118_39) );
AOI211_X1 g_126_38 (.ZN (n_126_38), .A (n_122_40), .B (n_119_40), .C1 (n_115_42), .C2 (n_116_40) );
AOI211_X1 g_128_37 (.ZN (n_128_37), .A (n_124_39), .B (n_121_39), .C1 (n_117_41), .C2 (n_114_41) );
AOI211_X1 g_130_36 (.ZN (n_130_36), .A (n_126_38), .B (n_120_41), .C1 (n_119_40), .C2 (n_113_43) );
AOI211_X1 g_132_35 (.ZN (n_132_35), .A (n_128_37), .B (n_122_40), .C1 (n_121_39), .C2 (n_115_42) );
AOI211_X1 g_134_34 (.ZN (n_134_34), .A (n_130_36), .B (n_124_39), .C1 (n_120_41), .C2 (n_117_41) );
AOI211_X1 g_136_33 (.ZN (n_136_33), .A (n_132_35), .B (n_126_38), .C1 (n_122_40), .C2 (n_119_40) );
AOI211_X1 g_138_32 (.ZN (n_138_32), .A (n_134_34), .B (n_128_37), .C1 (n_124_39), .C2 (n_121_39) );
AOI211_X1 g_140_31 (.ZN (n_140_31), .A (n_136_33), .B (n_130_36), .C1 (n_126_38), .C2 (n_120_41) );
AOI211_X1 g_139_33 (.ZN (n_139_33), .A (n_138_32), .B (n_132_35), .C1 (n_128_37), .C2 (n_122_40) );
AOI211_X1 g_137_34 (.ZN (n_137_34), .A (n_140_31), .B (n_134_34), .C1 (n_130_36), .C2 (n_124_39) );
AOI211_X1 g_135_35 (.ZN (n_135_35), .A (n_139_33), .B (n_136_33), .C1 (n_132_35), .C2 (n_126_38) );
AOI211_X1 g_133_36 (.ZN (n_133_36), .A (n_137_34), .B (n_138_32), .C1 (n_134_34), .C2 (n_128_37) );
AOI211_X1 g_131_37 (.ZN (n_131_37), .A (n_135_35), .B (n_140_31), .C1 (n_136_33), .C2 (n_130_36) );
AOI211_X1 g_129_38 (.ZN (n_129_38), .A (n_133_36), .B (n_139_33), .C1 (n_138_32), .C2 (n_132_35) );
AOI211_X1 g_127_39 (.ZN (n_127_39), .A (n_131_37), .B (n_137_34), .C1 (n_140_31), .C2 (n_134_34) );
AOI211_X1 g_125_38 (.ZN (n_125_38), .A (n_129_38), .B (n_135_35), .C1 (n_139_33), .C2 (n_136_33) );
AOI211_X1 g_123_39 (.ZN (n_123_39), .A (n_127_39), .B (n_133_36), .C1 (n_137_34), .C2 (n_138_32) );
AOI211_X1 g_121_40 (.ZN (n_121_40), .A (n_125_38), .B (n_131_37), .C1 (n_135_35), .C2 (n_140_31) );
AOI211_X1 g_119_41 (.ZN (n_119_41), .A (n_123_39), .B (n_129_38), .C1 (n_133_36), .C2 (n_139_33) );
AOI211_X1 g_117_42 (.ZN (n_117_42), .A (n_121_40), .B (n_127_39), .C1 (n_131_37), .C2 (n_137_34) );
AOI211_X1 g_115_43 (.ZN (n_115_43), .A (n_119_41), .B (n_125_38), .C1 (n_129_38), .C2 (n_135_35) );
AOI211_X1 g_113_44 (.ZN (n_113_44), .A (n_117_42), .B (n_123_39), .C1 (n_127_39), .C2 (n_133_36) );
AOI211_X1 g_111_45 (.ZN (n_111_45), .A (n_115_43), .B (n_121_40), .C1 (n_125_38), .C2 (n_131_37) );
AOI211_X1 g_109_44 (.ZN (n_109_44), .A (n_113_44), .B (n_119_41), .C1 (n_123_39), .C2 (n_129_38) );
AOI211_X1 g_107_45 (.ZN (n_107_45), .A (n_111_45), .B (n_117_42), .C1 (n_121_40), .C2 (n_127_39) );
AOI211_X1 g_105_46 (.ZN (n_105_46), .A (n_109_44), .B (n_115_43), .C1 (n_119_41), .C2 (n_125_38) );
AOI211_X1 g_103_47 (.ZN (n_103_47), .A (n_107_45), .B (n_113_44), .C1 (n_117_42), .C2 (n_123_39) );
AOI211_X1 g_101_48 (.ZN (n_101_48), .A (n_105_46), .B (n_111_45), .C1 (n_115_43), .C2 (n_121_40) );
AOI211_X1 g_99_49 (.ZN (n_99_49), .A (n_103_47), .B (n_109_44), .C1 (n_113_44), .C2 (n_119_41) );
AOI211_X1 g_97_50 (.ZN (n_97_50), .A (n_101_48), .B (n_107_45), .C1 (n_111_45), .C2 (n_117_42) );
AOI211_X1 g_95_51 (.ZN (n_95_51), .A (n_99_49), .B (n_105_46), .C1 (n_109_44), .C2 (n_115_43) );
AOI211_X1 g_94_53 (.ZN (n_94_53), .A (n_97_50), .B (n_103_47), .C1 (n_107_45), .C2 (n_113_44) );
AOI211_X1 g_93_51 (.ZN (n_93_51), .A (n_95_51), .B (n_101_48), .C1 (n_105_46), .C2 (n_111_45) );
AOI211_X1 g_95_50 (.ZN (n_95_50), .A (n_94_53), .B (n_99_49), .C1 (n_103_47), .C2 (n_109_44) );
AOI211_X1 g_97_49 (.ZN (n_97_49), .A (n_93_51), .B (n_97_50), .C1 (n_101_48), .C2 (n_107_45) );
AOI211_X1 g_99_48 (.ZN (n_99_48), .A (n_95_50), .B (n_95_51), .C1 (n_99_49), .C2 (n_105_46) );
AOI211_X1 g_101_47 (.ZN (n_101_47), .A (n_97_49), .B (n_94_53), .C1 (n_97_50), .C2 (n_103_47) );
AOI211_X1 g_103_46 (.ZN (n_103_46), .A (n_99_48), .B (n_93_51), .C1 (n_95_51), .C2 (n_101_48) );
AOI211_X1 g_105_47 (.ZN (n_105_47), .A (n_101_47), .B (n_95_50), .C1 (n_94_53), .C2 (n_99_49) );
AOI211_X1 g_103_48 (.ZN (n_103_48), .A (n_103_46), .B (n_97_49), .C1 (n_93_51), .C2 (n_97_50) );
AOI211_X1 g_101_49 (.ZN (n_101_49), .A (n_105_47), .B (n_99_48), .C1 (n_95_50), .C2 (n_95_51) );
AOI211_X1 g_99_50 (.ZN (n_99_50), .A (n_103_48), .B (n_101_47), .C1 (n_97_49), .C2 (n_94_53) );
AOI211_X1 g_97_51 (.ZN (n_97_51), .A (n_101_49), .B (n_103_46), .C1 (n_99_48), .C2 (n_93_51) );
AOI211_X1 g_95_52 (.ZN (n_95_52), .A (n_99_50), .B (n_105_47), .C1 (n_101_47), .C2 (n_95_50) );
AOI211_X1 g_93_53 (.ZN (n_93_53), .A (n_97_51), .B (n_103_48), .C1 (n_103_46), .C2 (n_97_49) );
AOI211_X1 g_92_51 (.ZN (n_92_51), .A (n_95_52), .B (n_101_49), .C1 (n_105_47), .C2 (n_99_48) );
AOI211_X1 g_91_53 (.ZN (n_91_53), .A (n_93_53), .B (n_99_50), .C1 (n_103_48), .C2 (n_101_47) );
AOI211_X1 g_89_54 (.ZN (n_89_54), .A (n_92_51), .B (n_97_51), .C1 (n_101_49), .C2 (n_103_46) );
AOI211_X1 g_90_52 (.ZN (n_90_52), .A (n_91_53), .B (n_95_52), .C1 (n_99_50), .C2 (n_105_47) );
AOI211_X1 g_88_53 (.ZN (n_88_53), .A (n_89_54), .B (n_93_53), .C1 (n_97_51), .C2 (n_103_48) );
AOI211_X1 g_87_55 (.ZN (n_87_55), .A (n_90_52), .B (n_92_51), .C1 (n_95_52), .C2 (n_101_49) );
AOI211_X1 g_85_56 (.ZN (n_85_56), .A (n_88_53), .B (n_91_53), .C1 (n_93_53), .C2 (n_99_50) );
AOI211_X1 g_86_54 (.ZN (n_86_54), .A (n_87_55), .B (n_89_54), .C1 (n_92_51), .C2 (n_97_51) );
AOI211_X1 g_84_55 (.ZN (n_84_55), .A (n_85_56), .B (n_90_52), .C1 (n_91_53), .C2 (n_95_52) );
AOI211_X1 g_83_57 (.ZN (n_83_57), .A (n_86_54), .B (n_88_53), .C1 (n_89_54), .C2 (n_93_53) );
AOI211_X1 g_81_58 (.ZN (n_81_58), .A (n_84_55), .B (n_87_55), .C1 (n_90_52), .C2 (n_92_51) );
AOI211_X1 g_82_56 (.ZN (n_82_56), .A (n_83_57), .B (n_85_56), .C1 (n_88_53), .C2 (n_91_53) );
AOI211_X1 g_80_57 (.ZN (n_80_57), .A (n_81_58), .B (n_86_54), .C1 (n_87_55), .C2 (n_89_54) );
AOI211_X1 g_79_59 (.ZN (n_79_59), .A (n_82_56), .B (n_84_55), .C1 (n_85_56), .C2 (n_90_52) );
AOI211_X1 g_77_60 (.ZN (n_77_60), .A (n_80_57), .B (n_83_57), .C1 (n_86_54), .C2 (n_88_53) );
AOI211_X1 g_78_58 (.ZN (n_78_58), .A (n_79_59), .B (n_81_58), .C1 (n_84_55), .C2 (n_87_55) );
AOI211_X1 g_76_59 (.ZN (n_76_59), .A (n_77_60), .B (n_82_56), .C1 (n_83_57), .C2 (n_85_56) );
AOI211_X1 g_75_61 (.ZN (n_75_61), .A (n_78_58), .B (n_80_57), .C1 (n_81_58), .C2 (n_86_54) );
AOI211_X1 g_73_62 (.ZN (n_73_62), .A (n_76_59), .B (n_79_59), .C1 (n_82_56), .C2 (n_84_55) );
AOI211_X1 g_74_60 (.ZN (n_74_60), .A (n_75_61), .B (n_77_60), .C1 (n_80_57), .C2 (n_83_57) );
AOI211_X1 g_72_61 (.ZN (n_72_61), .A (n_73_62), .B (n_78_58), .C1 (n_79_59), .C2 (n_81_58) );
AOI211_X1 g_71_63 (.ZN (n_71_63), .A (n_74_60), .B (n_76_59), .C1 (n_77_60), .C2 (n_82_56) );
AOI211_X1 g_69_64 (.ZN (n_69_64), .A (n_72_61), .B (n_75_61), .C1 (n_78_58), .C2 (n_80_57) );
AOI211_X1 g_70_62 (.ZN (n_70_62), .A (n_71_63), .B (n_73_62), .C1 (n_76_59), .C2 (n_79_59) );
AOI211_X1 g_68_63 (.ZN (n_68_63), .A (n_69_64), .B (n_74_60), .C1 (n_75_61), .C2 (n_77_60) );
AOI211_X1 g_67_65 (.ZN (n_67_65), .A (n_70_62), .B (n_72_61), .C1 (n_73_62), .C2 (n_78_58) );
AOI211_X1 g_65_66 (.ZN (n_65_66), .A (n_68_63), .B (n_71_63), .C1 (n_74_60), .C2 (n_76_59) );
AOI211_X1 g_66_64 (.ZN (n_66_64), .A (n_67_65), .B (n_69_64), .C1 (n_72_61), .C2 (n_75_61) );
AOI211_X1 g_64_65 (.ZN (n_64_65), .A (n_65_66), .B (n_70_62), .C1 (n_71_63), .C2 (n_73_62) );
AOI211_X1 g_63_67 (.ZN (n_63_67), .A (n_66_64), .B (n_68_63), .C1 (n_69_64), .C2 (n_74_60) );
AOI211_X1 g_61_68 (.ZN (n_61_68), .A (n_64_65), .B (n_67_65), .C1 (n_70_62), .C2 (n_72_61) );
AOI211_X1 g_62_66 (.ZN (n_62_66), .A (n_63_67), .B (n_65_66), .C1 (n_68_63), .C2 (n_71_63) );
AOI211_X1 g_60_67 (.ZN (n_60_67), .A (n_61_68), .B (n_66_64), .C1 (n_67_65), .C2 (n_69_64) );
AOI211_X1 g_59_69 (.ZN (n_59_69), .A (n_62_66), .B (n_64_65), .C1 (n_65_66), .C2 (n_70_62) );
AOI211_X1 g_57_70 (.ZN (n_57_70), .A (n_60_67), .B (n_63_67), .C1 (n_66_64), .C2 (n_68_63) );
AOI211_X1 g_58_68 (.ZN (n_58_68), .A (n_59_69), .B (n_61_68), .C1 (n_64_65), .C2 (n_67_65) );
AOI211_X1 g_56_69 (.ZN (n_56_69), .A (n_57_70), .B (n_62_66), .C1 (n_63_67), .C2 (n_65_66) );
AOI211_X1 g_54_70 (.ZN (n_54_70), .A (n_58_68), .B (n_60_67), .C1 (n_61_68), .C2 (n_66_64) );
AOI211_X1 g_52_71 (.ZN (n_52_71), .A (n_56_69), .B (n_59_69), .C1 (n_62_66), .C2 (n_64_65) );
AOI211_X1 g_50_72 (.ZN (n_50_72), .A (n_54_70), .B (n_57_70), .C1 (n_60_67), .C2 (n_63_67) );
AOI211_X1 g_48_73 (.ZN (n_48_73), .A (n_52_71), .B (n_58_68), .C1 (n_59_69), .C2 (n_61_68) );
AOI211_X1 g_46_74 (.ZN (n_46_74), .A (n_50_72), .B (n_56_69), .C1 (n_57_70), .C2 (n_62_66) );
AOI211_X1 g_44_75 (.ZN (n_44_75), .A (n_48_73), .B (n_54_70), .C1 (n_58_68), .C2 (n_60_67) );
AOI211_X1 g_42_76 (.ZN (n_42_76), .A (n_46_74), .B (n_52_71), .C1 (n_56_69), .C2 (n_59_69) );
AOI211_X1 g_40_77 (.ZN (n_40_77), .A (n_44_75), .B (n_50_72), .C1 (n_54_70), .C2 (n_57_70) );
AOI211_X1 g_38_78 (.ZN (n_38_78), .A (n_42_76), .B (n_48_73), .C1 (n_52_71), .C2 (n_58_68) );
AOI211_X1 g_36_79 (.ZN (n_36_79), .A (n_40_77), .B (n_46_74), .C1 (n_50_72), .C2 (n_56_69) );
AOI211_X1 g_34_80 (.ZN (n_34_80), .A (n_38_78), .B (n_44_75), .C1 (n_48_73), .C2 (n_54_70) );
AOI211_X1 g_33_82 (.ZN (n_33_82), .A (n_36_79), .B (n_42_76), .C1 (n_46_74), .C2 (n_52_71) );
AOI211_X1 g_31_81 (.ZN (n_31_81), .A (n_34_80), .B (n_40_77), .C1 (n_44_75), .C2 (n_50_72) );
AOI211_X1 g_29_82 (.ZN (n_29_82), .A (n_33_82), .B (n_38_78), .C1 (n_42_76), .C2 (n_48_73) );
AOI211_X1 g_27_83 (.ZN (n_27_83), .A (n_31_81), .B (n_36_79), .C1 (n_40_77), .C2 (n_46_74) );
AOI211_X1 g_25_84 (.ZN (n_25_84), .A (n_29_82), .B (n_34_80), .C1 (n_38_78), .C2 (n_44_75) );
AOI211_X1 g_23_85 (.ZN (n_23_85), .A (n_27_83), .B (n_33_82), .C1 (n_36_79), .C2 (n_42_76) );
AOI211_X1 g_21_86 (.ZN (n_21_86), .A (n_25_84), .B (n_31_81), .C1 (n_34_80), .C2 (n_40_77) );
AOI211_X1 g_19_87 (.ZN (n_19_87), .A (n_23_85), .B (n_29_82), .C1 (n_33_82), .C2 (n_38_78) );
AOI211_X1 g_17_88 (.ZN (n_17_88), .A (n_21_86), .B (n_27_83), .C1 (n_31_81), .C2 (n_36_79) );
AOI211_X1 g_15_89 (.ZN (n_15_89), .A (n_19_87), .B (n_25_84), .C1 (n_29_82), .C2 (n_34_80) );
AOI211_X1 g_13_90 (.ZN (n_13_90), .A (n_17_88), .B (n_23_85), .C1 (n_27_83), .C2 (n_33_82) );
AOI211_X1 g_11_91 (.ZN (n_11_91), .A (n_15_89), .B (n_21_86), .C1 (n_25_84), .C2 (n_31_81) );
AOI211_X1 g_9_92 (.ZN (n_9_92), .A (n_13_90), .B (n_19_87), .C1 (n_23_85), .C2 (n_29_82) );
AOI211_X1 g_7_93 (.ZN (n_7_93), .A (n_11_91), .B (n_17_88), .C1 (n_21_86), .C2 (n_27_83) );
AOI211_X1 g_6_95 (.ZN (n_6_95), .A (n_9_92), .B (n_15_89), .C1 (n_19_87), .C2 (n_25_84) );
AOI211_X1 g_5_93 (.ZN (n_5_93), .A (n_7_93), .B (n_13_90), .C1 (n_17_88), .C2 (n_23_85) );
AOI211_X1 g_7_92 (.ZN (n_7_92), .A (n_6_95), .B (n_11_91), .C1 (n_15_89), .C2 (n_21_86) );
AOI211_X1 g_9_91 (.ZN (n_9_91), .A (n_5_93), .B (n_9_92), .C1 (n_13_90), .C2 (n_19_87) );
AOI211_X1 g_11_90 (.ZN (n_11_90), .A (n_7_92), .B (n_7_93), .C1 (n_11_91), .C2 (n_17_88) );
AOI211_X1 g_10_92 (.ZN (n_10_92), .A (n_9_91), .B (n_6_95), .C1 (n_9_92), .C2 (n_15_89) );
AOI211_X1 g_12_91 (.ZN (n_12_91), .A (n_11_90), .B (n_5_93), .C1 (n_7_93), .C2 (n_13_90) );
AOI211_X1 g_14_90 (.ZN (n_14_90), .A (n_10_92), .B (n_7_92), .C1 (n_6_95), .C2 (n_11_91) );
AOI211_X1 g_16_89 (.ZN (n_16_89), .A (n_12_91), .B (n_9_91), .C1 (n_5_93), .C2 (n_9_92) );
AOI211_X1 g_18_88 (.ZN (n_18_88), .A (n_14_90), .B (n_11_90), .C1 (n_7_92), .C2 (n_7_93) );
AOI211_X1 g_20_87 (.ZN (n_20_87), .A (n_16_89), .B (n_10_92), .C1 (n_9_91), .C2 (n_6_95) );
AOI211_X1 g_22_86 (.ZN (n_22_86), .A (n_18_88), .B (n_12_91), .C1 (n_11_90), .C2 (n_5_93) );
AOI211_X1 g_23_84 (.ZN (n_23_84), .A (n_20_87), .B (n_14_90), .C1 (n_10_92), .C2 (n_7_92) );
AOI211_X1 g_25_85 (.ZN (n_25_85), .A (n_22_86), .B (n_16_89), .C1 (n_12_91), .C2 (n_9_91) );
AOI211_X1 g_27_84 (.ZN (n_27_84), .A (n_23_84), .B (n_18_88), .C1 (n_14_90), .C2 (n_11_90) );
AOI211_X1 g_29_83 (.ZN (n_29_83), .A (n_25_85), .B (n_20_87), .C1 (n_16_89), .C2 (n_10_92) );
AOI211_X1 g_31_82 (.ZN (n_31_82), .A (n_27_84), .B (n_22_86), .C1 (n_18_88), .C2 (n_12_91) );
AOI211_X1 g_33_81 (.ZN (n_33_81), .A (n_29_83), .B (n_23_84), .C1 (n_20_87), .C2 (n_14_90) );
AOI211_X1 g_35_80 (.ZN (n_35_80), .A (n_31_82), .B (n_25_85), .C1 (n_22_86), .C2 (n_16_89) );
AOI211_X1 g_37_79 (.ZN (n_37_79), .A (n_33_81), .B (n_27_84), .C1 (n_23_84), .C2 (n_18_88) );
AOI211_X1 g_39_78 (.ZN (n_39_78), .A (n_35_80), .B (n_29_83), .C1 (n_25_85), .C2 (n_20_87) );
AOI211_X1 g_41_77 (.ZN (n_41_77), .A (n_37_79), .B (n_31_82), .C1 (n_27_84), .C2 (n_22_86) );
AOI211_X1 g_43_76 (.ZN (n_43_76), .A (n_39_78), .B (n_33_81), .C1 (n_29_83), .C2 (n_23_84) );
AOI211_X1 g_45_75 (.ZN (n_45_75), .A (n_41_77), .B (n_35_80), .C1 (n_31_82), .C2 (n_25_85) );
AOI211_X1 g_47_74 (.ZN (n_47_74), .A (n_43_76), .B (n_37_79), .C1 (n_33_81), .C2 (n_27_84) );
AOI211_X1 g_49_73 (.ZN (n_49_73), .A (n_45_75), .B (n_39_78), .C1 (n_35_80), .C2 (n_29_83) );
AOI211_X1 g_51_72 (.ZN (n_51_72), .A (n_47_74), .B (n_41_77), .C1 (n_37_79), .C2 (n_31_82) );
AOI211_X1 g_53_71 (.ZN (n_53_71), .A (n_49_73), .B (n_43_76), .C1 (n_39_78), .C2 (n_33_81) );
AOI211_X1 g_52_73 (.ZN (n_52_73), .A (n_51_72), .B (n_45_75), .C1 (n_41_77), .C2 (n_35_80) );
AOI211_X1 g_54_72 (.ZN (n_54_72), .A (n_53_71), .B (n_47_74), .C1 (n_43_76), .C2 (n_37_79) );
AOI211_X1 g_56_71 (.ZN (n_56_71), .A (n_52_73), .B (n_49_73), .C1 (n_45_75), .C2 (n_39_78) );
AOI211_X1 g_58_70 (.ZN (n_58_70), .A (n_54_72), .B (n_51_72), .C1 (n_47_74), .C2 (n_41_77) );
AOI211_X1 g_60_69 (.ZN (n_60_69), .A (n_56_71), .B (n_53_71), .C1 (n_49_73), .C2 (n_43_76) );
AOI211_X1 g_59_71 (.ZN (n_59_71), .A (n_58_70), .B (n_52_73), .C1 (n_51_72), .C2 (n_45_75) );
AOI211_X1 g_61_70 (.ZN (n_61_70), .A (n_60_69), .B (n_54_72), .C1 (n_53_71), .C2 (n_47_74) );
AOI211_X1 g_63_69 (.ZN (n_63_69), .A (n_59_71), .B (n_56_71), .C1 (n_52_73), .C2 (n_49_73) );
AOI211_X1 g_64_67 (.ZN (n_64_67), .A (n_61_70), .B (n_58_70), .C1 (n_54_72), .C2 (n_51_72) );
AOI211_X1 g_66_66 (.ZN (n_66_66), .A (n_63_69), .B (n_60_69), .C1 (n_56_71), .C2 (n_53_71) );
AOI211_X1 g_68_65 (.ZN (n_68_65), .A (n_64_67), .B (n_59_71), .C1 (n_58_70), .C2 (n_52_73) );
AOI211_X1 g_70_64 (.ZN (n_70_64), .A (n_66_66), .B (n_61_70), .C1 (n_60_69), .C2 (n_54_72) );
AOI211_X1 g_72_63 (.ZN (n_72_63), .A (n_68_65), .B (n_63_69), .C1 (n_59_71), .C2 (n_56_71) );
AOI211_X1 g_74_62 (.ZN (n_74_62), .A (n_70_64), .B (n_64_67), .C1 (n_61_70), .C2 (n_58_70) );
AOI211_X1 g_76_61 (.ZN (n_76_61), .A (n_72_63), .B (n_66_66), .C1 (n_63_69), .C2 (n_60_69) );
AOI211_X1 g_78_60 (.ZN (n_78_60), .A (n_74_62), .B (n_68_65), .C1 (n_64_67), .C2 (n_59_71) );
AOI211_X1 g_80_59 (.ZN (n_80_59), .A (n_76_61), .B (n_70_64), .C1 (n_66_66), .C2 (n_61_70) );
AOI211_X1 g_82_58 (.ZN (n_82_58), .A (n_78_60), .B (n_72_63), .C1 (n_68_65), .C2 (n_63_69) );
AOI211_X1 g_84_57 (.ZN (n_84_57), .A (n_80_59), .B (n_74_62), .C1 (n_70_64), .C2 (n_64_67) );
AOI211_X1 g_86_56 (.ZN (n_86_56), .A (n_82_58), .B (n_76_61), .C1 (n_72_63), .C2 (n_66_66) );
AOI211_X1 g_88_55 (.ZN (n_88_55), .A (n_84_57), .B (n_78_60), .C1 (n_74_62), .C2 (n_68_65) );
AOI211_X1 g_90_54 (.ZN (n_90_54), .A (n_86_56), .B (n_80_59), .C1 (n_76_61), .C2 (n_70_64) );
AOI211_X1 g_92_53 (.ZN (n_92_53), .A (n_88_55), .B (n_82_58), .C1 (n_78_60), .C2 (n_72_63) );
AOI211_X1 g_94_52 (.ZN (n_94_52), .A (n_90_54), .B (n_84_57), .C1 (n_80_59), .C2 (n_74_62) );
AOI211_X1 g_96_51 (.ZN (n_96_51), .A (n_92_53), .B (n_86_56), .C1 (n_82_58), .C2 (n_76_61) );
AOI211_X1 g_98_50 (.ZN (n_98_50), .A (n_94_52), .B (n_88_55), .C1 (n_84_57), .C2 (n_78_60) );
AOI211_X1 g_100_49 (.ZN (n_100_49), .A (n_96_51), .B (n_90_54), .C1 (n_86_56), .C2 (n_80_59) );
AOI211_X1 g_102_48 (.ZN (n_102_48), .A (n_98_50), .B (n_92_53), .C1 (n_88_55), .C2 (n_82_58) );
AOI211_X1 g_104_47 (.ZN (n_104_47), .A (n_100_49), .B (n_94_52), .C1 (n_90_54), .C2 (n_84_57) );
AOI211_X1 g_106_46 (.ZN (n_106_46), .A (n_102_48), .B (n_96_51), .C1 (n_92_53), .C2 (n_86_56) );
AOI211_X1 g_108_45 (.ZN (n_108_45), .A (n_104_47), .B (n_98_50), .C1 (n_94_52), .C2 (n_88_55) );
AOI211_X1 g_110_44 (.ZN (n_110_44), .A (n_106_46), .B (n_100_49), .C1 (n_96_51), .C2 (n_90_54) );
AOI211_X1 g_109_46 (.ZN (n_109_46), .A (n_108_45), .B (n_102_48), .C1 (n_98_50), .C2 (n_92_53) );
AOI211_X1 g_107_47 (.ZN (n_107_47), .A (n_110_44), .B (n_104_47), .C1 (n_100_49), .C2 (n_94_52) );
AOI211_X1 g_105_48 (.ZN (n_105_48), .A (n_109_46), .B (n_106_46), .C1 (n_102_48), .C2 (n_96_51) );
AOI211_X1 g_103_49 (.ZN (n_103_49), .A (n_107_47), .B (n_108_45), .C1 (n_104_47), .C2 (n_98_50) );
AOI211_X1 g_101_50 (.ZN (n_101_50), .A (n_105_48), .B (n_110_44), .C1 (n_106_46), .C2 (n_100_49) );
AOI211_X1 g_99_51 (.ZN (n_99_51), .A (n_103_49), .B (n_109_46), .C1 (n_108_45), .C2 (n_102_48) );
AOI211_X1 g_97_52 (.ZN (n_97_52), .A (n_101_50), .B (n_107_47), .C1 (n_110_44), .C2 (n_104_47) );
AOI211_X1 g_95_53 (.ZN (n_95_53), .A (n_99_51), .B (n_105_48), .C1 (n_109_46), .C2 (n_106_46) );
AOI211_X1 g_93_54 (.ZN (n_93_54), .A (n_97_52), .B (n_103_49), .C1 (n_107_47), .C2 (n_108_45) );
AOI211_X1 g_91_55 (.ZN (n_91_55), .A (n_95_53), .B (n_101_50), .C1 (n_105_48), .C2 (n_110_44) );
AOI211_X1 g_89_56 (.ZN (n_89_56), .A (n_93_54), .B (n_99_51), .C1 (n_103_49), .C2 (n_109_46) );
AOI211_X1 g_87_57 (.ZN (n_87_57), .A (n_91_55), .B (n_97_52), .C1 (n_101_50), .C2 (n_107_47) );
AOI211_X1 g_85_58 (.ZN (n_85_58), .A (n_89_56), .B (n_95_53), .C1 (n_99_51), .C2 (n_105_48) );
AOI211_X1 g_83_59 (.ZN (n_83_59), .A (n_87_57), .B (n_93_54), .C1 (n_97_52), .C2 (n_103_49) );
AOI211_X1 g_81_60 (.ZN (n_81_60), .A (n_85_58), .B (n_91_55), .C1 (n_95_53), .C2 (n_101_50) );
AOI211_X1 g_79_61 (.ZN (n_79_61), .A (n_83_59), .B (n_89_56), .C1 (n_93_54), .C2 (n_99_51) );
AOI211_X1 g_77_62 (.ZN (n_77_62), .A (n_81_60), .B (n_87_57), .C1 (n_91_55), .C2 (n_97_52) );
AOI211_X1 g_75_63 (.ZN (n_75_63), .A (n_79_61), .B (n_85_58), .C1 (n_89_56), .C2 (n_95_53) );
AOI211_X1 g_73_64 (.ZN (n_73_64), .A (n_77_62), .B (n_83_59), .C1 (n_87_57), .C2 (n_93_54) );
AOI211_X1 g_71_65 (.ZN (n_71_65), .A (n_75_63), .B (n_81_60), .C1 (n_85_58), .C2 (n_91_55) );
AOI211_X1 g_69_66 (.ZN (n_69_66), .A (n_73_64), .B (n_79_61), .C1 (n_83_59), .C2 (n_89_56) );
AOI211_X1 g_67_67 (.ZN (n_67_67), .A (n_71_65), .B (n_77_62), .C1 (n_81_60), .C2 (n_87_57) );
AOI211_X1 g_65_68 (.ZN (n_65_68), .A (n_69_66), .B (n_75_63), .C1 (n_79_61), .C2 (n_85_58) );
AOI211_X1 g_64_70 (.ZN (n_64_70), .A (n_67_67), .B (n_73_64), .C1 (n_77_62), .C2 (n_83_59) );
AOI211_X1 g_63_68 (.ZN (n_63_68), .A (n_65_68), .B (n_71_65), .C1 (n_75_63), .C2 (n_81_60) );
AOI211_X1 g_65_67 (.ZN (n_65_67), .A (n_64_70), .B (n_69_66), .C1 (n_73_64), .C2 (n_79_61) );
AOI211_X1 g_67_66 (.ZN (n_67_66), .A (n_63_68), .B (n_67_67), .C1 (n_71_65), .C2 (n_77_62) );
AOI211_X1 g_69_65 (.ZN (n_69_65), .A (n_65_67), .B (n_65_68), .C1 (n_69_66), .C2 (n_75_63) );
AOI211_X1 g_71_64 (.ZN (n_71_64), .A (n_67_66), .B (n_64_70), .C1 (n_67_67), .C2 (n_73_64) );
AOI211_X1 g_73_63 (.ZN (n_73_63), .A (n_69_65), .B (n_63_68), .C1 (n_65_68), .C2 (n_71_65) );
AOI211_X1 g_75_62 (.ZN (n_75_62), .A (n_71_64), .B (n_65_67), .C1 (n_64_70), .C2 (n_69_66) );
AOI211_X1 g_77_61 (.ZN (n_77_61), .A (n_73_63), .B (n_67_66), .C1 (n_63_68), .C2 (n_67_67) );
AOI211_X1 g_79_60 (.ZN (n_79_60), .A (n_75_62), .B (n_69_65), .C1 (n_65_67), .C2 (n_65_68) );
AOI211_X1 g_81_59 (.ZN (n_81_59), .A (n_77_61), .B (n_71_64), .C1 (n_67_66), .C2 (n_64_70) );
AOI211_X1 g_83_58 (.ZN (n_83_58), .A (n_79_60), .B (n_73_63), .C1 (n_69_65), .C2 (n_63_68) );
AOI211_X1 g_85_57 (.ZN (n_85_57), .A (n_81_59), .B (n_75_62), .C1 (n_71_64), .C2 (n_65_67) );
AOI211_X1 g_87_56 (.ZN (n_87_56), .A (n_83_58), .B (n_77_61), .C1 (n_73_63), .C2 (n_67_66) );
AOI211_X1 g_89_55 (.ZN (n_89_55), .A (n_85_57), .B (n_79_60), .C1 (n_75_62), .C2 (n_69_65) );
AOI211_X1 g_91_54 (.ZN (n_91_54), .A (n_87_56), .B (n_81_59), .C1 (n_77_61), .C2 (n_71_64) );
AOI211_X1 g_90_56 (.ZN (n_90_56), .A (n_89_55), .B (n_83_58), .C1 (n_79_60), .C2 (n_73_63) );
AOI211_X1 g_92_55 (.ZN (n_92_55), .A (n_91_54), .B (n_85_57), .C1 (n_81_59), .C2 (n_75_62) );
AOI211_X1 g_94_54 (.ZN (n_94_54), .A (n_90_56), .B (n_87_56), .C1 (n_83_58), .C2 (n_77_61) );
AOI211_X1 g_96_53 (.ZN (n_96_53), .A (n_92_55), .B (n_89_55), .C1 (n_85_57), .C2 (n_79_60) );
AOI211_X1 g_98_52 (.ZN (n_98_52), .A (n_94_54), .B (n_91_54), .C1 (n_87_56), .C2 (n_81_59) );
AOI211_X1 g_100_51 (.ZN (n_100_51), .A (n_96_53), .B (n_90_56), .C1 (n_89_55), .C2 (n_83_58) );
AOI211_X1 g_102_50 (.ZN (n_102_50), .A (n_98_52), .B (n_92_55), .C1 (n_91_54), .C2 (n_85_57) );
AOI211_X1 g_104_49 (.ZN (n_104_49), .A (n_100_51), .B (n_94_54), .C1 (n_90_56), .C2 (n_87_56) );
AOI211_X1 g_106_48 (.ZN (n_106_48), .A (n_102_50), .B (n_96_53), .C1 (n_92_55), .C2 (n_89_55) );
AOI211_X1 g_108_47 (.ZN (n_108_47), .A (n_104_49), .B (n_98_52), .C1 (n_94_54), .C2 (n_91_54) );
AOI211_X1 g_110_46 (.ZN (n_110_46), .A (n_106_48), .B (n_100_51), .C1 (n_96_53), .C2 (n_90_56) );
AOI211_X1 g_112_45 (.ZN (n_112_45), .A (n_108_47), .B (n_102_50), .C1 (n_98_52), .C2 (n_92_55) );
AOI211_X1 g_114_44 (.ZN (n_114_44), .A (n_110_46), .B (n_104_49), .C1 (n_100_51), .C2 (n_94_54) );
AOI211_X1 g_116_43 (.ZN (n_116_43), .A (n_112_45), .B (n_106_48), .C1 (n_102_50), .C2 (n_96_53) );
AOI211_X1 g_118_42 (.ZN (n_118_42), .A (n_114_44), .B (n_108_47), .C1 (n_104_49), .C2 (n_98_52) );
AOI211_X1 g_117_44 (.ZN (n_117_44), .A (n_116_43), .B (n_110_46), .C1 (n_106_48), .C2 (n_100_51) );
AOI211_X1 g_116_42 (.ZN (n_116_42), .A (n_118_42), .B (n_112_45), .C1 (n_108_47), .C2 (n_102_50) );
AOI211_X1 g_118_41 (.ZN (n_118_41), .A (n_117_44), .B (n_114_44), .C1 (n_110_46), .C2 (n_104_49) );
AOI211_X1 g_120_40 (.ZN (n_120_40), .A (n_116_42), .B (n_116_43), .C1 (n_112_45), .C2 (n_106_48) );
AOI211_X1 g_122_39 (.ZN (n_122_39), .A (n_118_41), .B (n_118_42), .C1 (n_114_44), .C2 (n_108_47) );
AOI211_X1 g_124_40 (.ZN (n_124_40), .A (n_120_40), .B (n_117_44), .C1 (n_116_43), .C2 (n_110_46) );
AOI211_X1 g_122_41 (.ZN (n_122_41), .A (n_122_39), .B (n_116_42), .C1 (n_118_42), .C2 (n_112_45) );
AOI211_X1 g_120_42 (.ZN (n_120_42), .A (n_124_40), .B (n_118_41), .C1 (n_117_44), .C2 (n_114_44) );
AOI211_X1 g_118_43 (.ZN (n_118_43), .A (n_122_41), .B (n_120_40), .C1 (n_116_42), .C2 (n_116_43) );
AOI211_X1 g_116_44 (.ZN (n_116_44), .A (n_120_42), .B (n_122_39), .C1 (n_118_41), .C2 (n_118_42) );
AOI211_X1 g_114_43 (.ZN (n_114_43), .A (n_118_43), .B (n_124_40), .C1 (n_120_40), .C2 (n_117_44) );
AOI211_X1 g_112_44 (.ZN (n_112_44), .A (n_116_44), .B (n_122_41), .C1 (n_122_39), .C2 (n_116_42) );
AOI211_X1 g_110_45 (.ZN (n_110_45), .A (n_114_43), .B (n_120_42), .C1 (n_124_40), .C2 (n_118_41) );
AOI211_X1 g_108_46 (.ZN (n_108_46), .A (n_112_44), .B (n_118_43), .C1 (n_122_41), .C2 (n_120_40) );
AOI211_X1 g_106_47 (.ZN (n_106_47), .A (n_110_45), .B (n_116_44), .C1 (n_120_42), .C2 (n_122_39) );
AOI211_X1 g_104_48 (.ZN (n_104_48), .A (n_108_46), .B (n_114_43), .C1 (n_118_43), .C2 (n_124_40) );
AOI211_X1 g_102_49 (.ZN (n_102_49), .A (n_106_47), .B (n_112_44), .C1 (n_116_44), .C2 (n_122_41) );
AOI211_X1 g_100_50 (.ZN (n_100_50), .A (n_104_48), .B (n_110_45), .C1 (n_114_43), .C2 (n_120_42) );
AOI211_X1 g_98_51 (.ZN (n_98_51), .A (n_102_49), .B (n_108_46), .C1 (n_112_44), .C2 (n_118_43) );
AOI211_X1 g_96_52 (.ZN (n_96_52), .A (n_100_50), .B (n_106_47), .C1 (n_110_45), .C2 (n_116_44) );
AOI211_X1 g_95_54 (.ZN (n_95_54), .A (n_98_51), .B (n_104_48), .C1 (n_108_46), .C2 (n_114_43) );
AOI211_X1 g_97_53 (.ZN (n_97_53), .A (n_96_52), .B (n_102_49), .C1 (n_106_47), .C2 (n_112_44) );
AOI211_X1 g_99_52 (.ZN (n_99_52), .A (n_95_54), .B (n_100_50), .C1 (n_104_48), .C2 (n_110_45) );
AOI211_X1 g_101_51 (.ZN (n_101_51), .A (n_97_53), .B (n_98_51), .C1 (n_102_49), .C2 (n_108_46) );
AOI211_X1 g_103_50 (.ZN (n_103_50), .A (n_99_52), .B (n_96_52), .C1 (n_100_50), .C2 (n_106_47) );
AOI211_X1 g_105_49 (.ZN (n_105_49), .A (n_101_51), .B (n_95_54), .C1 (n_98_51), .C2 (n_104_48) );
AOI211_X1 g_107_48 (.ZN (n_107_48), .A (n_103_50), .B (n_97_53), .C1 (n_96_52), .C2 (n_102_49) );
AOI211_X1 g_109_47 (.ZN (n_109_47), .A (n_105_49), .B (n_99_52), .C1 (n_95_54), .C2 (n_100_50) );
AOI211_X1 g_111_46 (.ZN (n_111_46), .A (n_107_48), .B (n_101_51), .C1 (n_97_53), .C2 (n_98_51) );
AOI211_X1 g_113_45 (.ZN (n_113_45), .A (n_109_47), .B (n_103_50), .C1 (n_99_52), .C2 (n_96_52) );
AOI211_X1 g_115_44 (.ZN (n_115_44), .A (n_111_46), .B (n_105_49), .C1 (n_101_51), .C2 (n_95_54) );
AOI211_X1 g_117_43 (.ZN (n_117_43), .A (n_113_45), .B (n_107_48), .C1 (n_103_50), .C2 (n_97_53) );
AOI211_X1 g_119_42 (.ZN (n_119_42), .A (n_115_44), .B (n_109_47), .C1 (n_105_49), .C2 (n_99_52) );
AOI211_X1 g_121_41 (.ZN (n_121_41), .A (n_117_43), .B (n_111_46), .C1 (n_107_48), .C2 (n_101_51) );
AOI211_X1 g_123_40 (.ZN (n_123_40), .A (n_119_42), .B (n_113_45), .C1 (n_109_47), .C2 (n_103_50) );
AOI211_X1 g_125_39 (.ZN (n_125_39), .A (n_121_41), .B (n_115_44), .C1 (n_111_46), .C2 (n_105_49) );
AOI211_X1 g_124_41 (.ZN (n_124_41), .A (n_123_40), .B (n_117_43), .C1 (n_113_45), .C2 (n_107_48) );
AOI211_X1 g_126_40 (.ZN (n_126_40), .A (n_125_39), .B (n_119_42), .C1 (n_115_44), .C2 (n_109_47) );
AOI211_X1 g_128_39 (.ZN (n_128_39), .A (n_124_41), .B (n_121_41), .C1 (n_117_43), .C2 (n_111_46) );
AOI211_X1 g_130_38 (.ZN (n_130_38), .A (n_126_40), .B (n_123_40), .C1 (n_119_42), .C2 (n_113_45) );
AOI211_X1 g_132_37 (.ZN (n_132_37), .A (n_128_39), .B (n_125_39), .C1 (n_121_41), .C2 (n_115_44) );
AOI211_X1 g_134_36 (.ZN (n_134_36), .A (n_130_38), .B (n_124_41), .C1 (n_123_40), .C2 (n_117_43) );
AOI211_X1 g_136_35 (.ZN (n_136_35), .A (n_132_37), .B (n_126_40), .C1 (n_125_39), .C2 (n_119_42) );
AOI211_X1 g_138_34 (.ZN (n_138_34), .A (n_134_36), .B (n_128_39), .C1 (n_124_41), .C2 (n_121_41) );
AOI211_X1 g_140_33 (.ZN (n_140_33), .A (n_136_35), .B (n_130_38), .C1 (n_126_40), .C2 (n_123_40) );
AOI211_X1 g_142_32 (.ZN (n_142_32), .A (n_138_34), .B (n_132_37), .C1 (n_128_39), .C2 (n_125_39) );
AOI211_X1 g_144_31 (.ZN (n_144_31), .A (n_140_33), .B (n_134_36), .C1 (n_130_38), .C2 (n_124_41) );
AOI211_X1 g_146_30 (.ZN (n_146_30), .A (n_142_32), .B (n_136_35), .C1 (n_132_37), .C2 (n_126_40) );
AOI211_X1 g_147_32 (.ZN (n_147_32), .A (n_144_31), .B (n_138_34), .C1 (n_134_36), .C2 (n_128_39) );
AOI211_X1 g_149_33 (.ZN (n_149_33), .A (n_146_30), .B (n_140_33), .C1 (n_136_35), .C2 (n_130_38) );
AOI211_X1 g_148_31 (.ZN (n_148_31), .A (n_147_32), .B (n_142_32), .C1 (n_138_34), .C2 (n_132_37) );
AOI211_X1 g_146_32 (.ZN (n_146_32), .A (n_149_33), .B (n_144_31), .C1 (n_140_33), .C2 (n_134_36) );
AOI211_X1 g_147_34 (.ZN (n_147_34), .A (n_148_31), .B (n_146_30), .C1 (n_142_32), .C2 (n_136_35) );
AOI211_X1 g_145_33 (.ZN (n_145_33), .A (n_146_32), .B (n_147_32), .C1 (n_144_31), .C2 (n_138_34) );
AOI211_X1 g_143_34 (.ZN (n_143_34), .A (n_147_34), .B (n_149_33), .C1 (n_146_30), .C2 (n_140_33) );
AOI211_X1 g_141_33 (.ZN (n_141_33), .A (n_145_33), .B (n_148_31), .C1 (n_147_32), .C2 (n_142_32) );
AOI211_X1 g_139_34 (.ZN (n_139_34), .A (n_143_34), .B (n_146_32), .C1 (n_149_33), .C2 (n_144_31) );
AOI211_X1 g_137_35 (.ZN (n_137_35), .A (n_141_33), .B (n_147_34), .C1 (n_148_31), .C2 (n_146_30) );
AOI211_X1 g_135_36 (.ZN (n_135_36), .A (n_139_34), .B (n_145_33), .C1 (n_146_32), .C2 (n_147_32) );
AOI211_X1 g_133_37 (.ZN (n_133_37), .A (n_137_35), .B (n_143_34), .C1 (n_147_34), .C2 (n_149_33) );
AOI211_X1 g_131_38 (.ZN (n_131_38), .A (n_135_36), .B (n_141_33), .C1 (n_145_33), .C2 (n_148_31) );
AOI211_X1 g_129_39 (.ZN (n_129_39), .A (n_133_37), .B (n_139_34), .C1 (n_143_34), .C2 (n_146_32) );
AOI211_X1 g_127_40 (.ZN (n_127_40), .A (n_131_38), .B (n_137_35), .C1 (n_141_33), .C2 (n_147_34) );
AOI211_X1 g_125_41 (.ZN (n_125_41), .A (n_129_39), .B (n_135_36), .C1 (n_139_34), .C2 (n_145_33) );
AOI211_X1 g_123_42 (.ZN (n_123_42), .A (n_127_40), .B (n_133_37), .C1 (n_137_35), .C2 (n_143_34) );
AOI211_X1 g_121_43 (.ZN (n_121_43), .A (n_125_41), .B (n_131_38), .C1 (n_135_36), .C2 (n_141_33) );
AOI211_X1 g_119_44 (.ZN (n_119_44), .A (n_123_42), .B (n_129_39), .C1 (n_133_37), .C2 (n_139_34) );
AOI211_X1 g_117_45 (.ZN (n_117_45), .A (n_121_43), .B (n_127_40), .C1 (n_131_38), .C2 (n_137_35) );
AOI211_X1 g_115_46 (.ZN (n_115_46), .A (n_119_44), .B (n_125_41), .C1 (n_129_39), .C2 (n_135_36) );
AOI211_X1 g_113_47 (.ZN (n_113_47), .A (n_117_45), .B (n_123_42), .C1 (n_127_40), .C2 (n_133_37) );
AOI211_X1 g_114_45 (.ZN (n_114_45), .A (n_115_46), .B (n_121_43), .C1 (n_125_41), .C2 (n_131_38) );
AOI211_X1 g_112_46 (.ZN (n_112_46), .A (n_113_47), .B (n_119_44), .C1 (n_123_42), .C2 (n_129_39) );
AOI211_X1 g_110_47 (.ZN (n_110_47), .A (n_114_45), .B (n_117_45), .C1 (n_121_43), .C2 (n_127_40) );
AOI211_X1 g_108_48 (.ZN (n_108_48), .A (n_112_46), .B (n_115_46), .C1 (n_119_44), .C2 (n_125_41) );
AOI211_X1 g_106_49 (.ZN (n_106_49), .A (n_110_47), .B (n_113_47), .C1 (n_117_45), .C2 (n_123_42) );
AOI211_X1 g_104_50 (.ZN (n_104_50), .A (n_108_48), .B (n_114_45), .C1 (n_115_46), .C2 (n_121_43) );
AOI211_X1 g_102_51 (.ZN (n_102_51), .A (n_106_49), .B (n_112_46), .C1 (n_113_47), .C2 (n_119_44) );
AOI211_X1 g_100_52 (.ZN (n_100_52), .A (n_104_50), .B (n_110_47), .C1 (n_114_45), .C2 (n_117_45) );
AOI211_X1 g_98_53 (.ZN (n_98_53), .A (n_102_51), .B (n_108_48), .C1 (n_112_46), .C2 (n_115_46) );
AOI211_X1 g_96_54 (.ZN (n_96_54), .A (n_100_52), .B (n_106_49), .C1 (n_110_47), .C2 (n_113_47) );
AOI211_X1 g_94_55 (.ZN (n_94_55), .A (n_98_53), .B (n_104_50), .C1 (n_108_48), .C2 (n_114_45) );
AOI211_X1 g_92_56 (.ZN (n_92_56), .A (n_96_54), .B (n_102_51), .C1 (n_106_49), .C2 (n_112_46) );
AOI211_X1 g_90_57 (.ZN (n_90_57), .A (n_94_55), .B (n_100_52), .C1 (n_104_50), .C2 (n_110_47) );
AOI211_X1 g_88_58 (.ZN (n_88_58), .A (n_92_56), .B (n_98_53), .C1 (n_102_51), .C2 (n_108_48) );
AOI211_X1 g_86_59 (.ZN (n_86_59), .A (n_90_57), .B (n_96_54), .C1 (n_100_52), .C2 (n_106_49) );
AOI211_X1 g_84_60 (.ZN (n_84_60), .A (n_88_58), .B (n_94_55), .C1 (n_98_53), .C2 (n_104_50) );
AOI211_X1 g_82_61 (.ZN (n_82_61), .A (n_86_59), .B (n_92_56), .C1 (n_96_54), .C2 (n_102_51) );
AOI211_X1 g_80_62 (.ZN (n_80_62), .A (n_84_60), .B (n_90_57), .C1 (n_94_55), .C2 (n_100_52) );
AOI211_X1 g_78_63 (.ZN (n_78_63), .A (n_82_61), .B (n_88_58), .C1 (n_92_56), .C2 (n_98_53) );
AOI211_X1 g_76_64 (.ZN (n_76_64), .A (n_80_62), .B (n_86_59), .C1 (n_90_57), .C2 (n_96_54) );
AOI211_X1 g_74_65 (.ZN (n_74_65), .A (n_78_63), .B (n_84_60), .C1 (n_88_58), .C2 (n_94_55) );
AOI211_X1 g_72_66 (.ZN (n_72_66), .A (n_76_64), .B (n_82_61), .C1 (n_86_59), .C2 (n_92_56) );
AOI211_X1 g_70_67 (.ZN (n_70_67), .A (n_74_65), .B (n_80_62), .C1 (n_84_60), .C2 (n_90_57) );
AOI211_X1 g_68_68 (.ZN (n_68_68), .A (n_72_66), .B (n_78_63), .C1 (n_82_61), .C2 (n_88_58) );
AOI211_X1 g_66_69 (.ZN (n_66_69), .A (n_70_67), .B (n_76_64), .C1 (n_80_62), .C2 (n_86_59) );
AOI211_X1 g_65_71 (.ZN (n_65_71), .A (n_68_68), .B (n_74_65), .C1 (n_78_63), .C2 (n_84_60) );
AOI211_X1 g_64_69 (.ZN (n_64_69), .A (n_66_69), .B (n_72_66), .C1 (n_76_64), .C2 (n_82_61) );
AOI211_X1 g_66_68 (.ZN (n_66_68), .A (n_65_71), .B (n_70_67), .C1 (n_74_65), .C2 (n_80_62) );
AOI211_X1 g_68_67 (.ZN (n_68_67), .A (n_64_69), .B (n_68_68), .C1 (n_72_66), .C2 (n_78_63) );
AOI211_X1 g_70_66 (.ZN (n_70_66), .A (n_66_68), .B (n_66_69), .C1 (n_70_67), .C2 (n_76_64) );
AOI211_X1 g_72_65 (.ZN (n_72_65), .A (n_68_67), .B (n_65_71), .C1 (n_68_68), .C2 (n_74_65) );
AOI211_X1 g_74_64 (.ZN (n_74_64), .A (n_70_66), .B (n_64_69), .C1 (n_66_69), .C2 (n_72_66) );
AOI211_X1 g_76_63 (.ZN (n_76_63), .A (n_72_65), .B (n_66_68), .C1 (n_65_71), .C2 (n_70_67) );
AOI211_X1 g_78_62 (.ZN (n_78_62), .A (n_74_64), .B (n_68_67), .C1 (n_64_69), .C2 (n_68_68) );
AOI211_X1 g_80_61 (.ZN (n_80_61), .A (n_76_63), .B (n_70_66), .C1 (n_66_68), .C2 (n_66_69) );
AOI211_X1 g_82_60 (.ZN (n_82_60), .A (n_78_62), .B (n_72_65), .C1 (n_68_67), .C2 (n_65_71) );
AOI211_X1 g_84_59 (.ZN (n_84_59), .A (n_80_61), .B (n_74_64), .C1 (n_70_66), .C2 (n_64_69) );
AOI211_X1 g_86_58 (.ZN (n_86_58), .A (n_82_60), .B (n_76_63), .C1 (n_72_65), .C2 (n_66_68) );
AOI211_X1 g_88_57 (.ZN (n_88_57), .A (n_84_59), .B (n_78_62), .C1 (n_74_64), .C2 (n_68_67) );
AOI211_X1 g_87_59 (.ZN (n_87_59), .A (n_86_58), .B (n_80_61), .C1 (n_76_63), .C2 (n_70_66) );
AOI211_X1 g_89_58 (.ZN (n_89_58), .A (n_88_57), .B (n_82_60), .C1 (n_78_62), .C2 (n_72_65) );
AOI211_X1 g_91_57 (.ZN (n_91_57), .A (n_87_59), .B (n_84_59), .C1 (n_80_61), .C2 (n_74_64) );
AOI211_X1 g_93_56 (.ZN (n_93_56), .A (n_89_58), .B (n_86_58), .C1 (n_82_60), .C2 (n_76_63) );
AOI211_X1 g_95_55 (.ZN (n_95_55), .A (n_91_57), .B (n_88_57), .C1 (n_84_59), .C2 (n_78_62) );
AOI211_X1 g_97_54 (.ZN (n_97_54), .A (n_93_56), .B (n_87_59), .C1 (n_86_58), .C2 (n_80_61) );
AOI211_X1 g_99_53 (.ZN (n_99_53), .A (n_95_55), .B (n_89_58), .C1 (n_88_57), .C2 (n_82_60) );
AOI211_X1 g_101_52 (.ZN (n_101_52), .A (n_97_54), .B (n_91_57), .C1 (n_87_59), .C2 (n_84_59) );
AOI211_X1 g_103_51 (.ZN (n_103_51), .A (n_99_53), .B (n_93_56), .C1 (n_89_58), .C2 (n_86_58) );
AOI211_X1 g_105_50 (.ZN (n_105_50), .A (n_101_52), .B (n_95_55), .C1 (n_91_57), .C2 (n_88_57) );
AOI211_X1 g_107_49 (.ZN (n_107_49), .A (n_103_51), .B (n_97_54), .C1 (n_93_56), .C2 (n_87_59) );
AOI211_X1 g_109_48 (.ZN (n_109_48), .A (n_105_50), .B (n_99_53), .C1 (n_95_55), .C2 (n_89_58) );
AOI211_X1 g_111_47 (.ZN (n_111_47), .A (n_107_49), .B (n_101_52), .C1 (n_97_54), .C2 (n_91_57) );
AOI211_X1 g_113_46 (.ZN (n_113_46), .A (n_109_48), .B (n_103_51), .C1 (n_99_53), .C2 (n_93_56) );
AOI211_X1 g_115_45 (.ZN (n_115_45), .A (n_111_47), .B (n_105_50), .C1 (n_101_52), .C2 (n_95_55) );
AOI211_X1 g_114_47 (.ZN (n_114_47), .A (n_113_46), .B (n_107_49), .C1 (n_103_51), .C2 (n_97_54) );
AOI211_X1 g_116_46 (.ZN (n_116_46), .A (n_115_45), .B (n_109_48), .C1 (n_105_50), .C2 (n_99_53) );
AOI211_X1 g_118_45 (.ZN (n_118_45), .A (n_114_47), .B (n_111_47), .C1 (n_107_49), .C2 (n_101_52) );
AOI211_X1 g_119_43 (.ZN (n_119_43), .A (n_116_46), .B (n_113_46), .C1 (n_109_48), .C2 (n_103_51) );
AOI211_X1 g_121_42 (.ZN (n_121_42), .A (n_118_45), .B (n_115_45), .C1 (n_111_47), .C2 (n_105_50) );
AOI211_X1 g_123_41 (.ZN (n_123_41), .A (n_119_43), .B (n_114_47), .C1 (n_113_46), .C2 (n_107_49) );
AOI211_X1 g_125_40 (.ZN (n_125_40), .A (n_121_42), .B (n_116_46), .C1 (n_115_45), .C2 (n_109_48) );
AOI211_X1 g_124_42 (.ZN (n_124_42), .A (n_123_41), .B (n_118_45), .C1 (n_114_47), .C2 (n_111_47) );
AOI211_X1 g_126_41 (.ZN (n_126_41), .A (n_125_40), .B (n_119_43), .C1 (n_116_46), .C2 (n_113_46) );
AOI211_X1 g_128_40 (.ZN (n_128_40), .A (n_124_42), .B (n_121_42), .C1 (n_118_45), .C2 (n_115_45) );
AOI211_X1 g_130_39 (.ZN (n_130_39), .A (n_126_41), .B (n_123_41), .C1 (n_119_43), .C2 (n_114_47) );
AOI211_X1 g_132_38 (.ZN (n_132_38), .A (n_128_40), .B (n_125_40), .C1 (n_121_42), .C2 (n_116_46) );
AOI211_X1 g_134_37 (.ZN (n_134_37), .A (n_130_39), .B (n_124_42), .C1 (n_123_41), .C2 (n_118_45) );
AOI211_X1 g_136_36 (.ZN (n_136_36), .A (n_132_38), .B (n_126_41), .C1 (n_125_40), .C2 (n_119_43) );
AOI211_X1 g_138_35 (.ZN (n_138_35), .A (n_134_37), .B (n_128_40), .C1 (n_124_42), .C2 (n_121_42) );
AOI211_X1 g_140_34 (.ZN (n_140_34), .A (n_136_36), .B (n_130_39), .C1 (n_126_41), .C2 (n_123_41) );
AOI211_X1 g_142_33 (.ZN (n_142_33), .A (n_138_35), .B (n_132_38), .C1 (n_128_40), .C2 (n_125_40) );
AOI211_X1 g_141_35 (.ZN (n_141_35), .A (n_140_34), .B (n_134_37), .C1 (n_130_39), .C2 (n_124_42) );
AOI211_X1 g_139_36 (.ZN (n_139_36), .A (n_142_33), .B (n_136_36), .C1 (n_132_38), .C2 (n_126_41) );
AOI211_X1 g_137_37 (.ZN (n_137_37), .A (n_141_35), .B (n_138_35), .C1 (n_134_37), .C2 (n_128_40) );
AOI211_X1 g_135_38 (.ZN (n_135_38), .A (n_139_36), .B (n_140_34), .C1 (n_136_36), .C2 (n_130_39) );
AOI211_X1 g_133_39 (.ZN (n_133_39), .A (n_137_37), .B (n_142_33), .C1 (n_138_35), .C2 (n_132_38) );
AOI211_X1 g_131_40 (.ZN (n_131_40), .A (n_135_38), .B (n_141_35), .C1 (n_140_34), .C2 (n_134_37) );
AOI211_X1 g_129_41 (.ZN (n_129_41), .A (n_133_39), .B (n_139_36), .C1 (n_142_33), .C2 (n_136_36) );
AOI211_X1 g_127_42 (.ZN (n_127_42), .A (n_131_40), .B (n_137_37), .C1 (n_141_35), .C2 (n_138_35) );
AOI211_X1 g_125_43 (.ZN (n_125_43), .A (n_129_41), .B (n_135_38), .C1 (n_139_36), .C2 (n_140_34) );
AOI211_X1 g_123_44 (.ZN (n_123_44), .A (n_127_42), .B (n_133_39), .C1 (n_137_37), .C2 (n_142_33) );
AOI211_X1 g_122_42 (.ZN (n_122_42), .A (n_125_43), .B (n_131_40), .C1 (n_135_38), .C2 (n_141_35) );
AOI211_X1 g_120_43 (.ZN (n_120_43), .A (n_123_44), .B (n_129_41), .C1 (n_133_39), .C2 (n_139_36) );
AOI211_X1 g_118_44 (.ZN (n_118_44), .A (n_122_42), .B (n_127_42), .C1 (n_131_40), .C2 (n_137_37) );
AOI211_X1 g_116_45 (.ZN (n_116_45), .A (n_120_43), .B (n_125_43), .C1 (n_129_41), .C2 (n_135_38) );
AOI211_X1 g_114_46 (.ZN (n_114_46), .A (n_118_44), .B (n_123_44), .C1 (n_127_42), .C2 (n_133_39) );
AOI211_X1 g_112_47 (.ZN (n_112_47), .A (n_116_45), .B (n_122_42), .C1 (n_125_43), .C2 (n_131_40) );
AOI211_X1 g_110_48 (.ZN (n_110_48), .A (n_114_46), .B (n_120_43), .C1 (n_123_44), .C2 (n_129_41) );
AOI211_X1 g_108_49 (.ZN (n_108_49), .A (n_112_47), .B (n_118_44), .C1 (n_122_42), .C2 (n_127_42) );
AOI211_X1 g_106_50 (.ZN (n_106_50), .A (n_110_48), .B (n_116_45), .C1 (n_120_43), .C2 (n_125_43) );
AOI211_X1 g_104_51 (.ZN (n_104_51), .A (n_108_49), .B (n_114_46), .C1 (n_118_44), .C2 (n_123_44) );
AOI211_X1 g_102_52 (.ZN (n_102_52), .A (n_106_50), .B (n_112_47), .C1 (n_116_45), .C2 (n_122_42) );
AOI211_X1 g_100_53 (.ZN (n_100_53), .A (n_104_51), .B (n_110_48), .C1 (n_114_46), .C2 (n_120_43) );
AOI211_X1 g_98_54 (.ZN (n_98_54), .A (n_102_52), .B (n_108_49), .C1 (n_112_47), .C2 (n_118_44) );
AOI211_X1 g_96_55 (.ZN (n_96_55), .A (n_100_53), .B (n_106_50), .C1 (n_110_48), .C2 (n_116_45) );
AOI211_X1 g_94_56 (.ZN (n_94_56), .A (n_98_54), .B (n_104_51), .C1 (n_108_49), .C2 (n_114_46) );
AOI211_X1 g_92_57 (.ZN (n_92_57), .A (n_96_55), .B (n_102_52), .C1 (n_106_50), .C2 (n_112_47) );
AOI211_X1 g_93_55 (.ZN (n_93_55), .A (n_94_56), .B (n_100_53), .C1 (n_104_51), .C2 (n_110_48) );
AOI211_X1 g_91_56 (.ZN (n_91_56), .A (n_92_57), .B (n_98_54), .C1 (n_102_52), .C2 (n_108_49) );
AOI211_X1 g_89_57 (.ZN (n_89_57), .A (n_93_55), .B (n_96_55), .C1 (n_100_53), .C2 (n_106_50) );
AOI211_X1 g_87_58 (.ZN (n_87_58), .A (n_91_56), .B (n_94_56), .C1 (n_98_54), .C2 (n_104_51) );
AOI211_X1 g_85_59 (.ZN (n_85_59), .A (n_89_57), .B (n_92_57), .C1 (n_96_55), .C2 (n_102_52) );
AOI211_X1 g_83_60 (.ZN (n_83_60), .A (n_87_58), .B (n_93_55), .C1 (n_94_56), .C2 (n_100_53) );
AOI211_X1 g_81_61 (.ZN (n_81_61), .A (n_85_59), .B (n_91_56), .C1 (n_92_57), .C2 (n_98_54) );
AOI211_X1 g_79_62 (.ZN (n_79_62), .A (n_83_60), .B (n_89_57), .C1 (n_93_55), .C2 (n_96_55) );
AOI211_X1 g_77_63 (.ZN (n_77_63), .A (n_81_61), .B (n_87_58), .C1 (n_91_56), .C2 (n_94_56) );
AOI211_X1 g_75_64 (.ZN (n_75_64), .A (n_79_62), .B (n_85_59), .C1 (n_89_57), .C2 (n_92_57) );
AOI211_X1 g_73_65 (.ZN (n_73_65), .A (n_77_63), .B (n_83_60), .C1 (n_87_58), .C2 (n_93_55) );
AOI211_X1 g_71_66 (.ZN (n_71_66), .A (n_75_64), .B (n_81_61), .C1 (n_85_59), .C2 (n_91_56) );
AOI211_X1 g_69_67 (.ZN (n_69_67), .A (n_73_65), .B (n_79_62), .C1 (n_83_60), .C2 (n_89_57) );
AOI211_X1 g_67_68 (.ZN (n_67_68), .A (n_71_66), .B (n_77_63), .C1 (n_81_61), .C2 (n_87_58) );
AOI211_X1 g_65_69 (.ZN (n_65_69), .A (n_69_67), .B (n_75_64), .C1 (n_79_62), .C2 (n_85_59) );
AOI211_X1 g_63_70 (.ZN (n_63_70), .A (n_67_68), .B (n_73_65), .C1 (n_77_63), .C2 (n_83_60) );
AOI211_X1 g_61_69 (.ZN (n_61_69), .A (n_65_69), .B (n_71_66), .C1 (n_75_64), .C2 (n_81_61) );
AOI211_X1 g_59_70 (.ZN (n_59_70), .A (n_63_70), .B (n_69_67), .C1 (n_73_65), .C2 (n_79_62) );
AOI211_X1 g_57_71 (.ZN (n_57_71), .A (n_61_69), .B (n_67_68), .C1 (n_71_66), .C2 (n_77_63) );
AOI211_X1 g_55_72 (.ZN (n_55_72), .A (n_59_70), .B (n_65_69), .C1 (n_69_67), .C2 (n_75_64) );
AOI211_X1 g_53_73 (.ZN (n_53_73), .A (n_57_71), .B (n_63_70), .C1 (n_67_68), .C2 (n_73_65) );
AOI211_X1 g_51_74 (.ZN (n_51_74), .A (n_55_72), .B (n_61_69), .C1 (n_65_69), .C2 (n_71_66) );
AOI211_X1 g_49_75 (.ZN (n_49_75), .A (n_53_73), .B (n_59_70), .C1 (n_63_70), .C2 (n_69_67) );
AOI211_X1 g_47_76 (.ZN (n_47_76), .A (n_51_74), .B (n_57_71), .C1 (n_61_69), .C2 (n_67_68) );
AOI211_X1 g_45_77 (.ZN (n_45_77), .A (n_49_75), .B (n_55_72), .C1 (n_59_70), .C2 (n_65_69) );
AOI211_X1 g_43_78 (.ZN (n_43_78), .A (n_47_76), .B (n_53_73), .C1 (n_57_71), .C2 (n_63_70) );
AOI211_X1 g_41_79 (.ZN (n_41_79), .A (n_45_77), .B (n_51_74), .C1 (n_55_72), .C2 (n_61_69) );
AOI211_X1 g_39_80 (.ZN (n_39_80), .A (n_43_78), .B (n_49_75), .C1 (n_53_73), .C2 (n_59_70) );
AOI211_X1 g_37_81 (.ZN (n_37_81), .A (n_41_79), .B (n_47_76), .C1 (n_51_74), .C2 (n_57_71) );
AOI211_X1 g_35_82 (.ZN (n_35_82), .A (n_39_80), .B (n_45_77), .C1 (n_49_75), .C2 (n_55_72) );
AOI211_X1 g_36_80 (.ZN (n_36_80), .A (n_37_81), .B (n_43_78), .C1 (n_47_76), .C2 (n_53_73) );
AOI211_X1 g_34_81 (.ZN (n_34_81), .A (n_35_82), .B (n_41_79), .C1 (n_45_77), .C2 (n_51_74) );
AOI211_X1 g_32_82 (.ZN (n_32_82), .A (n_36_80), .B (n_39_80), .C1 (n_43_78), .C2 (n_49_75) );
AOI211_X1 g_30_83 (.ZN (n_30_83), .A (n_34_81), .B (n_37_81), .C1 (n_41_79), .C2 (n_47_76) );
AOI211_X1 g_28_84 (.ZN (n_28_84), .A (n_32_82), .B (n_35_82), .C1 (n_39_80), .C2 (n_45_77) );
AOI211_X1 g_26_85 (.ZN (n_26_85), .A (n_30_83), .B (n_36_80), .C1 (n_37_81), .C2 (n_43_78) );
AOI211_X1 g_24_84 (.ZN (n_24_84), .A (n_28_84), .B (n_34_81), .C1 (n_35_82), .C2 (n_41_79) );
AOI211_X1 g_22_85 (.ZN (n_22_85), .A (n_26_85), .B (n_32_82), .C1 (n_36_80), .C2 (n_39_80) );
AOI211_X1 g_20_86 (.ZN (n_20_86), .A (n_24_84), .B (n_30_83), .C1 (n_34_81), .C2 (n_37_81) );
AOI211_X1 g_18_87 (.ZN (n_18_87), .A (n_22_85), .B (n_28_84), .C1 (n_32_82), .C2 (n_35_82) );
AOI211_X1 g_16_88 (.ZN (n_16_88), .A (n_20_86), .B (n_26_85), .C1 (n_30_83), .C2 (n_36_80) );
AOI211_X1 g_14_89 (.ZN (n_14_89), .A (n_18_87), .B (n_24_84), .C1 (n_28_84), .C2 (n_34_81) );
AOI211_X1 g_12_90 (.ZN (n_12_90), .A (n_16_88), .B (n_22_85), .C1 (n_26_85), .C2 (n_32_82) );
AOI211_X1 g_10_91 (.ZN (n_10_91), .A (n_14_89), .B (n_20_86), .C1 (n_24_84), .C2 (n_30_83) );
AOI211_X1 g_9_93 (.ZN (n_9_93), .A (n_12_90), .B (n_18_87), .C1 (n_22_85), .C2 (n_28_84) );
AOI211_X1 g_11_92 (.ZN (n_11_92), .A (n_10_91), .B (n_16_88), .C1 (n_20_86), .C2 (n_26_85) );
AOI211_X1 g_13_91 (.ZN (n_13_91), .A (n_9_93), .B (n_14_89), .C1 (n_18_87), .C2 (n_24_84) );
AOI211_X1 g_15_90 (.ZN (n_15_90), .A (n_11_92), .B (n_12_90), .C1 (n_16_88), .C2 (n_22_85) );
AOI211_X1 g_17_89 (.ZN (n_17_89), .A (n_13_91), .B (n_10_91), .C1 (n_14_89), .C2 (n_20_86) );
AOI211_X1 g_19_88 (.ZN (n_19_88), .A (n_15_90), .B (n_9_93), .C1 (n_12_90), .C2 (n_18_87) );
AOI211_X1 g_21_87 (.ZN (n_21_87), .A (n_17_89), .B (n_11_92), .C1 (n_10_91), .C2 (n_16_88) );
AOI211_X1 g_23_86 (.ZN (n_23_86), .A (n_19_88), .B (n_13_91), .C1 (n_9_93), .C2 (n_14_89) );
AOI211_X1 g_22_88 (.ZN (n_22_88), .A (n_21_87), .B (n_15_90), .C1 (n_11_92), .C2 (n_12_90) );
AOI211_X1 g_24_87 (.ZN (n_24_87), .A (n_23_86), .B (n_17_89), .C1 (n_13_91), .C2 (n_10_91) );
AOI211_X1 g_26_86 (.ZN (n_26_86), .A (n_22_88), .B (n_19_88), .C1 (n_15_90), .C2 (n_9_93) );
AOI211_X1 g_24_85 (.ZN (n_24_85), .A (n_24_87), .B (n_21_87), .C1 (n_17_89), .C2 (n_11_92) );
AOI211_X1 g_23_87 (.ZN (n_23_87), .A (n_26_86), .B (n_23_86), .C1 (n_19_88), .C2 (n_13_91) );
AOI211_X1 g_25_86 (.ZN (n_25_86), .A (n_24_85), .B (n_22_88), .C1 (n_21_87), .C2 (n_15_90) );
AOI211_X1 g_24_88 (.ZN (n_24_88), .A (n_23_87), .B (n_24_87), .C1 (n_23_86), .C2 (n_17_89) );
AOI211_X1 g_22_87 (.ZN (n_22_87), .A (n_25_86), .B (n_26_86), .C1 (n_22_88), .C2 (n_19_88) );
AOI211_X1 g_24_86 (.ZN (n_24_86), .A (n_24_88), .B (n_24_85), .C1 (n_24_87), .C2 (n_21_87) );
AOI211_X1 g_26_87 (.ZN (n_26_87), .A (n_22_87), .B (n_23_87), .C1 (n_26_86), .C2 (n_23_86) );
AOI211_X1 g_28_86 (.ZN (n_28_86), .A (n_24_86), .B (n_25_86), .C1 (n_24_85), .C2 (n_22_88) );
AOI211_X1 g_29_84 (.ZN (n_29_84), .A (n_26_87), .B (n_24_88), .C1 (n_23_87), .C2 (n_24_87) );
AOI211_X1 g_31_83 (.ZN (n_31_83), .A (n_28_86), .B (n_22_87), .C1 (n_25_86), .C2 (n_26_86) );
AOI211_X1 g_30_85 (.ZN (n_30_85), .A (n_29_84), .B (n_24_86), .C1 (n_24_88), .C2 (n_24_85) );
AOI211_X1 g_32_84 (.ZN (n_32_84), .A (n_31_83), .B (n_26_87), .C1 (n_22_87), .C2 (n_23_87) );
AOI211_X1 g_34_83 (.ZN (n_34_83), .A (n_30_85), .B (n_28_86), .C1 (n_24_86), .C2 (n_25_86) );
AOI211_X1 g_35_81 (.ZN (n_35_81), .A (n_32_84), .B (n_29_84), .C1 (n_26_87), .C2 (n_24_88) );
AOI211_X1 g_37_80 (.ZN (n_37_80), .A (n_34_83), .B (n_31_83), .C1 (n_28_86), .C2 (n_22_87) );
AOI211_X1 g_39_79 (.ZN (n_39_79), .A (n_35_81), .B (n_30_85), .C1 (n_29_84), .C2 (n_24_86) );
AOI211_X1 g_41_78 (.ZN (n_41_78), .A (n_37_80), .B (n_32_84), .C1 (n_31_83), .C2 (n_26_87) );
AOI211_X1 g_43_77 (.ZN (n_43_77), .A (n_39_79), .B (n_34_83), .C1 (n_30_85), .C2 (n_28_86) );
AOI211_X1 g_45_76 (.ZN (n_45_76), .A (n_41_78), .B (n_35_81), .C1 (n_32_84), .C2 (n_29_84) );
AOI211_X1 g_47_75 (.ZN (n_47_75), .A (n_43_77), .B (n_37_80), .C1 (n_34_83), .C2 (n_31_83) );
AOI211_X1 g_49_74 (.ZN (n_49_74), .A (n_45_76), .B (n_39_79), .C1 (n_35_81), .C2 (n_30_85) );
AOI211_X1 g_51_73 (.ZN (n_51_73), .A (n_47_75), .B (n_41_78), .C1 (n_37_80), .C2 (n_32_84) );
AOI211_X1 g_53_72 (.ZN (n_53_72), .A (n_49_74), .B (n_43_77), .C1 (n_39_79), .C2 (n_34_83) );
AOI211_X1 g_55_71 (.ZN (n_55_71), .A (n_51_73), .B (n_45_76), .C1 (n_41_78), .C2 (n_35_81) );
AOI211_X1 g_57_72 (.ZN (n_57_72), .A (n_53_72), .B (n_47_75), .C1 (n_43_77), .C2 (n_37_80) );
AOI211_X1 g_55_73 (.ZN (n_55_73), .A (n_55_71), .B (n_49_74), .C1 (n_45_76), .C2 (n_39_79) );
AOI211_X1 g_53_74 (.ZN (n_53_74), .A (n_57_72), .B (n_51_73), .C1 (n_47_75), .C2 (n_41_78) );
AOI211_X1 g_51_75 (.ZN (n_51_75), .A (n_55_73), .B (n_53_72), .C1 (n_49_74), .C2 (n_43_77) );
AOI211_X1 g_49_76 (.ZN (n_49_76), .A (n_53_74), .B (n_55_71), .C1 (n_51_73), .C2 (n_45_76) );
AOI211_X1 g_50_74 (.ZN (n_50_74), .A (n_51_75), .B (n_57_72), .C1 (n_53_72), .C2 (n_47_75) );
AOI211_X1 g_48_75 (.ZN (n_48_75), .A (n_49_76), .B (n_55_73), .C1 (n_55_71), .C2 (n_49_74) );
AOI211_X1 g_46_76 (.ZN (n_46_76), .A (n_50_74), .B (n_53_74), .C1 (n_57_72), .C2 (n_51_73) );
AOI211_X1 g_44_77 (.ZN (n_44_77), .A (n_48_75), .B (n_51_75), .C1 (n_55_73), .C2 (n_53_72) );
AOI211_X1 g_42_78 (.ZN (n_42_78), .A (n_46_76), .B (n_49_76), .C1 (n_53_74), .C2 (n_55_71) );
AOI211_X1 g_40_79 (.ZN (n_40_79), .A (n_44_77), .B (n_50_74), .C1 (n_51_75), .C2 (n_57_72) );
AOI211_X1 g_38_80 (.ZN (n_38_80), .A (n_42_78), .B (n_48_75), .C1 (n_49_76), .C2 (n_55_73) );
AOI211_X1 g_36_81 (.ZN (n_36_81), .A (n_40_79), .B (n_46_76), .C1 (n_50_74), .C2 (n_53_74) );
AOI211_X1 g_34_82 (.ZN (n_34_82), .A (n_38_80), .B (n_44_77), .C1 (n_48_75), .C2 (n_51_75) );
AOI211_X1 g_32_83 (.ZN (n_32_83), .A (n_36_81), .B (n_42_78), .C1 (n_46_76), .C2 (n_49_76) );
AOI211_X1 g_30_84 (.ZN (n_30_84), .A (n_34_82), .B (n_40_79), .C1 (n_44_77), .C2 (n_50_74) );
AOI211_X1 g_28_85 (.ZN (n_28_85), .A (n_32_83), .B (n_38_80), .C1 (n_42_78), .C2 (n_48_75) );
AOI211_X1 g_27_87 (.ZN (n_27_87), .A (n_30_84), .B (n_36_81), .C1 (n_40_79), .C2 (n_46_76) );
AOI211_X1 g_29_86 (.ZN (n_29_86), .A (n_28_85), .B (n_34_82), .C1 (n_38_80), .C2 (n_44_77) );
AOI211_X1 g_31_85 (.ZN (n_31_85), .A (n_27_87), .B (n_32_83), .C1 (n_36_81), .C2 (n_42_78) );
AOI211_X1 g_33_84 (.ZN (n_33_84), .A (n_29_86), .B (n_30_84), .C1 (n_34_82), .C2 (n_40_79) );
AOI211_X1 g_35_83 (.ZN (n_35_83), .A (n_31_85), .B (n_28_85), .C1 (n_32_83), .C2 (n_38_80) );
AOI211_X1 g_37_82 (.ZN (n_37_82), .A (n_33_84), .B (n_27_87), .C1 (n_30_84), .C2 (n_36_81) );
AOI211_X1 g_39_81 (.ZN (n_39_81), .A (n_35_83), .B (n_29_86), .C1 (n_28_85), .C2 (n_34_82) );
AOI211_X1 g_41_80 (.ZN (n_41_80), .A (n_37_82), .B (n_31_85), .C1 (n_27_87), .C2 (n_32_83) );
AOI211_X1 g_43_79 (.ZN (n_43_79), .A (n_39_81), .B (n_33_84), .C1 (n_29_86), .C2 (n_30_84) );
AOI211_X1 g_45_78 (.ZN (n_45_78), .A (n_41_80), .B (n_35_83), .C1 (n_31_85), .C2 (n_28_85) );
AOI211_X1 g_47_77 (.ZN (n_47_77), .A (n_43_79), .B (n_37_82), .C1 (n_33_84), .C2 (n_27_87) );
AOI211_X1 g_46_79 (.ZN (n_46_79), .A (n_45_78), .B (n_39_81), .C1 (n_35_83), .C2 (n_29_86) );
AOI211_X1 g_44_78 (.ZN (n_44_78), .A (n_47_77), .B (n_41_80), .C1 (n_37_82), .C2 (n_31_85) );
AOI211_X1 g_46_77 (.ZN (n_46_77), .A (n_46_79), .B (n_43_79), .C1 (n_39_81), .C2 (n_33_84) );
AOI211_X1 g_48_76 (.ZN (n_48_76), .A (n_44_78), .B (n_45_78), .C1 (n_41_80), .C2 (n_35_83) );
AOI211_X1 g_50_75 (.ZN (n_50_75), .A (n_46_77), .B (n_47_77), .C1 (n_43_79), .C2 (n_37_82) );
AOI211_X1 g_52_74 (.ZN (n_52_74), .A (n_48_76), .B (n_46_79), .C1 (n_45_78), .C2 (n_39_81) );
AOI211_X1 g_54_73 (.ZN (n_54_73), .A (n_50_75), .B (n_44_78), .C1 (n_47_77), .C2 (n_41_80) );
AOI211_X1 g_56_72 (.ZN (n_56_72), .A (n_52_74), .B (n_46_77), .C1 (n_46_79), .C2 (n_43_79) );
AOI211_X1 g_55_74 (.ZN (n_55_74), .A (n_54_73), .B (n_48_76), .C1 (n_44_78), .C2 (n_45_78) );
AOI211_X1 g_57_73 (.ZN (n_57_73), .A (n_56_72), .B (n_50_75), .C1 (n_46_77), .C2 (n_47_77) );
AOI211_X1 g_59_72 (.ZN (n_59_72), .A (n_55_74), .B (n_52_74), .C1 (n_48_76), .C2 (n_46_79) );
AOI211_X1 g_61_71 (.ZN (n_61_71), .A (n_57_73), .B (n_54_73), .C1 (n_50_75), .C2 (n_44_78) );
AOI211_X1 g_63_72 (.ZN (n_63_72), .A (n_59_72), .B (n_56_72), .C1 (n_52_74), .C2 (n_46_77) );
AOI211_X1 g_62_70 (.ZN (n_62_70), .A (n_61_71), .B (n_55_74), .C1 (n_54_73), .C2 (n_48_76) );
AOI211_X1 g_60_71 (.ZN (n_60_71), .A (n_63_72), .B (n_57_73), .C1 (n_56_72), .C2 (n_50_75) );
AOI211_X1 g_58_72 (.ZN (n_58_72), .A (n_62_70), .B (n_59_72), .C1 (n_55_74), .C2 (n_52_74) );
AOI211_X1 g_56_73 (.ZN (n_56_73), .A (n_60_71), .B (n_61_71), .C1 (n_57_73), .C2 (n_54_73) );
AOI211_X1 g_54_74 (.ZN (n_54_74), .A (n_58_72), .B (n_63_72), .C1 (n_59_72), .C2 (n_56_72) );
AOI211_X1 g_52_75 (.ZN (n_52_75), .A (n_56_73), .B (n_62_70), .C1 (n_61_71), .C2 (n_55_74) );
AOI211_X1 g_50_76 (.ZN (n_50_76), .A (n_54_74), .B (n_60_71), .C1 (n_63_72), .C2 (n_57_73) );
AOI211_X1 g_48_77 (.ZN (n_48_77), .A (n_52_75), .B (n_58_72), .C1 (n_62_70), .C2 (n_59_72) );
AOI211_X1 g_46_78 (.ZN (n_46_78), .A (n_50_76), .B (n_56_73), .C1 (n_60_71), .C2 (n_61_71) );
AOI211_X1 g_44_79 (.ZN (n_44_79), .A (n_48_77), .B (n_54_74), .C1 (n_58_72), .C2 (n_63_72) );
AOI211_X1 g_42_80 (.ZN (n_42_80), .A (n_46_78), .B (n_52_75), .C1 (n_56_73), .C2 (n_62_70) );
AOI211_X1 g_40_81 (.ZN (n_40_81), .A (n_44_79), .B (n_50_76), .C1 (n_54_74), .C2 (n_60_71) );
AOI211_X1 g_38_82 (.ZN (n_38_82), .A (n_42_80), .B (n_48_77), .C1 (n_52_75), .C2 (n_58_72) );
AOI211_X1 g_36_83 (.ZN (n_36_83), .A (n_40_81), .B (n_46_78), .C1 (n_50_76), .C2 (n_56_73) );
AOI211_X1 g_34_84 (.ZN (n_34_84), .A (n_38_82), .B (n_44_79), .C1 (n_48_77), .C2 (n_54_74) );
AOI211_X1 g_32_85 (.ZN (n_32_85), .A (n_36_83), .B (n_42_80), .C1 (n_46_78), .C2 (n_52_75) );
AOI211_X1 g_33_83 (.ZN (n_33_83), .A (n_34_84), .B (n_40_81), .C1 (n_44_79), .C2 (n_50_76) );
AOI211_X1 g_31_84 (.ZN (n_31_84), .A (n_32_85), .B (n_38_82), .C1 (n_42_80), .C2 (n_48_77) );
AOI211_X1 g_29_85 (.ZN (n_29_85), .A (n_33_83), .B (n_36_83), .C1 (n_40_81), .C2 (n_46_78) );
AOI211_X1 g_27_86 (.ZN (n_27_86), .A (n_31_84), .B (n_34_84), .C1 (n_38_82), .C2 (n_44_79) );
AOI211_X1 g_25_87 (.ZN (n_25_87), .A (n_29_85), .B (n_32_85), .C1 (n_36_83), .C2 (n_42_80) );
AOI211_X1 g_23_88 (.ZN (n_23_88), .A (n_27_86), .B (n_33_83), .C1 (n_34_84), .C2 (n_40_81) );
AOI211_X1 g_21_89 (.ZN (n_21_89), .A (n_25_87), .B (n_31_84), .C1 (n_32_85), .C2 (n_38_82) );
AOI211_X1 g_19_90 (.ZN (n_19_90), .A (n_23_88), .B (n_29_85), .C1 (n_33_83), .C2 (n_36_83) );
AOI211_X1 g_20_88 (.ZN (n_20_88), .A (n_21_89), .B (n_27_86), .C1 (n_31_84), .C2 (n_34_84) );
AOI211_X1 g_18_89 (.ZN (n_18_89), .A (n_19_90), .B (n_25_87), .C1 (n_29_85), .C2 (n_32_85) );
AOI211_X1 g_16_90 (.ZN (n_16_90), .A (n_20_88), .B (n_23_88), .C1 (n_27_86), .C2 (n_33_83) );
AOI211_X1 g_14_91 (.ZN (n_14_91), .A (n_18_89), .B (n_21_89), .C1 (n_25_87), .C2 (n_31_84) );
AOI211_X1 g_12_92 (.ZN (n_12_92), .A (n_16_90), .B (n_19_90), .C1 (n_23_88), .C2 (n_29_85) );
AOI211_X1 g_10_93 (.ZN (n_10_93), .A (n_14_91), .B (n_20_88), .C1 (n_21_89), .C2 (n_27_86) );
AOI211_X1 g_8_94 (.ZN (n_8_94), .A (n_12_92), .B (n_18_89), .C1 (n_19_90), .C2 (n_25_87) );
AOI211_X1 g_10_95 (.ZN (n_10_95), .A (n_10_93), .B (n_16_90), .C1 (n_20_88), .C2 (n_23_88) );
AOI211_X1 g_11_93 (.ZN (n_11_93), .A (n_8_94), .B (n_14_91), .C1 (n_18_89), .C2 (n_21_89) );
AOI211_X1 g_13_92 (.ZN (n_13_92), .A (n_10_95), .B (n_12_92), .C1 (n_16_90), .C2 (n_19_90) );
AOI211_X1 g_15_91 (.ZN (n_15_91), .A (n_11_93), .B (n_10_93), .C1 (n_14_91), .C2 (n_20_88) );
AOI211_X1 g_17_90 (.ZN (n_17_90), .A (n_13_92), .B (n_8_94), .C1 (n_12_92), .C2 (n_18_89) );
AOI211_X1 g_19_89 (.ZN (n_19_89), .A (n_15_91), .B (n_10_95), .C1 (n_10_93), .C2 (n_16_90) );
AOI211_X1 g_21_88 (.ZN (n_21_88), .A (n_17_90), .B (n_11_93), .C1 (n_8_94), .C2 (n_14_91) );
AOI211_X1 g_20_90 (.ZN (n_20_90), .A (n_19_89), .B (n_13_92), .C1 (n_10_95), .C2 (n_12_92) );
AOI211_X1 g_22_89 (.ZN (n_22_89), .A (n_21_88), .B (n_15_91), .C1 (n_11_93), .C2 (n_10_93) );
AOI211_X1 g_21_91 (.ZN (n_21_91), .A (n_20_90), .B (n_17_90), .C1 (n_13_92), .C2 (n_8_94) );
AOI211_X1 g_20_89 (.ZN (n_20_89), .A (n_22_89), .B (n_19_89), .C1 (n_15_91), .C2 (n_10_95) );
AOI211_X1 g_18_90 (.ZN (n_18_90), .A (n_21_91), .B (n_21_88), .C1 (n_17_90), .C2 (n_11_93) );
AOI211_X1 g_16_91 (.ZN (n_16_91), .A (n_20_89), .B (n_20_90), .C1 (n_19_89), .C2 (n_13_92) );
AOI211_X1 g_14_92 (.ZN (n_14_92), .A (n_18_90), .B (n_22_89), .C1 (n_21_88), .C2 (n_15_91) );
AOI211_X1 g_12_93 (.ZN (n_12_93), .A (n_16_91), .B (n_21_91), .C1 (n_20_90), .C2 (n_17_90) );
AOI211_X1 g_10_94 (.ZN (n_10_94), .A (n_14_92), .B (n_20_89), .C1 (n_22_89), .C2 (n_19_89) );
AOI211_X1 g_8_93 (.ZN (n_8_93), .A (n_12_93), .B (n_18_90), .C1 (n_21_91), .C2 (n_21_88) );
AOI211_X1 g_6_94 (.ZN (n_6_94), .A (n_10_94), .B (n_16_91), .C1 (n_20_89), .C2 (n_20_90) );
AOI211_X1 g_4_95 (.ZN (n_4_95), .A (n_8_93), .B (n_14_92), .C1 (n_18_90), .C2 (n_22_89) );
AOI211_X1 g_3_97 (.ZN (n_3_97), .A (n_6_94), .B (n_12_93), .C1 (n_16_91), .C2 (n_21_91) );
AOI211_X1 g_5_96 (.ZN (n_5_96), .A (n_4_95), .B (n_10_94), .C1 (n_14_92), .C2 (n_20_89) );
AOI211_X1 g_7_95 (.ZN (n_7_95), .A (n_3_97), .B (n_8_93), .C1 (n_12_93), .C2 (n_18_90) );
AOI211_X1 g_9_94 (.ZN (n_9_94), .A (n_5_96), .B (n_6_94), .C1 (n_10_94), .C2 (n_16_91) );
AOI211_X1 g_8_96 (.ZN (n_8_96), .A (n_7_95), .B (n_4_95), .C1 (n_8_93), .C2 (n_14_92) );
AOI211_X1 g_7_94 (.ZN (n_7_94), .A (n_9_94), .B (n_3_97), .C1 (n_6_94), .C2 (n_12_93) );
AOI211_X1 g_5_95 (.ZN (n_5_95), .A (n_8_96), .B (n_5_96), .C1 (n_4_95), .C2 (n_10_94) );
AOI211_X1 g_3_96 (.ZN (n_3_96), .A (n_7_94), .B (n_7_95), .C1 (n_3_97), .C2 (n_8_93) );
AOI211_X1 g_2_98 (.ZN (n_2_98), .A (n_5_95), .B (n_9_94), .C1 (n_5_96), .C2 (n_6_94) );
AOI211_X1 g_1_100 (.ZN (n_1_100), .A (n_3_96), .B (n_8_96), .C1 (n_7_95), .C2 (n_4_95) );
AOI211_X1 g_3_99 (.ZN (n_3_99), .A (n_2_98), .B (n_7_94), .C1 (n_9_94), .C2 (n_3_97) );
AOI211_X1 g_4_97 (.ZN (n_4_97), .A (n_1_100), .B (n_5_95), .C1 (n_8_96), .C2 (n_5_96) );
AOI211_X1 g_6_96 (.ZN (n_6_96), .A (n_3_99), .B (n_3_96), .C1 (n_7_94), .C2 (n_7_95) );
AOI211_X1 g_8_95 (.ZN (n_8_95), .A (n_4_97), .B (n_2_98), .C1 (n_5_95), .C2 (n_9_94) );
AOI211_X1 g_7_97 (.ZN (n_7_97), .A (n_6_96), .B (n_1_100), .C1 (n_3_96), .C2 (n_8_96) );
AOI211_X1 g_5_98 (.ZN (n_5_98), .A (n_8_95), .B (n_3_99), .C1 (n_2_98), .C2 (n_7_94) );
AOI211_X1 g_6_100 (.ZN (n_6_100), .A (n_7_97), .B (n_4_97), .C1 (n_1_100), .C2 (n_5_95) );
AOI211_X1 g_4_99 (.ZN (n_4_99), .A (n_5_98), .B (n_6_96), .C1 (n_3_99), .C2 (n_3_96) );
AOI211_X1 g_5_97 (.ZN (n_5_97), .A (n_6_100), .B (n_8_95), .C1 (n_4_97), .C2 (n_2_98) );
AOI211_X1 g_7_96 (.ZN (n_7_96), .A (n_4_99), .B (n_7_97), .C1 (n_6_96), .C2 (n_1_100) );
AOI211_X1 g_9_95 (.ZN (n_9_95), .A (n_5_97), .B (n_5_98), .C1 (n_8_95), .C2 (n_3_99) );
AOI211_X1 g_11_94 (.ZN (n_11_94), .A (n_7_96), .B (n_6_100), .C1 (n_7_97), .C2 (n_4_97) );
AOI211_X1 g_13_93 (.ZN (n_13_93), .A (n_9_95), .B (n_4_99), .C1 (n_5_98), .C2 (n_6_96) );
AOI211_X1 g_15_92 (.ZN (n_15_92), .A (n_11_94), .B (n_5_97), .C1 (n_6_100), .C2 (n_8_95) );
AOI211_X1 g_17_91 (.ZN (n_17_91), .A (n_13_93), .B (n_7_96), .C1 (n_4_99), .C2 (n_7_97) );
AOI211_X1 g_19_92 (.ZN (n_19_92), .A (n_15_92), .B (n_9_95), .C1 (n_5_97), .C2 (n_5_98) );
AOI211_X1 g_17_93 (.ZN (n_17_93), .A (n_17_91), .B (n_11_94), .C1 (n_7_96), .C2 (n_6_100) );
AOI211_X1 g_18_91 (.ZN (n_18_91), .A (n_19_92), .B (n_13_93), .C1 (n_9_95), .C2 (n_4_99) );
AOI211_X1 g_16_92 (.ZN (n_16_92), .A (n_17_93), .B (n_15_92), .C1 (n_11_94), .C2 (n_5_97) );
AOI211_X1 g_14_93 (.ZN (n_14_93), .A (n_18_91), .B (n_17_91), .C1 (n_13_93), .C2 (n_7_96) );
AOI211_X1 g_12_94 (.ZN (n_12_94), .A (n_16_92), .B (n_19_92), .C1 (n_15_92), .C2 (n_9_95) );
AOI211_X1 g_11_96 (.ZN (n_11_96), .A (n_14_93), .B (n_17_93), .C1 (n_17_91), .C2 (n_11_94) );
AOI211_X1 g_13_95 (.ZN (n_13_95), .A (n_12_94), .B (n_18_91), .C1 (n_19_92), .C2 (n_13_93) );
AOI211_X1 g_15_94 (.ZN (n_15_94), .A (n_11_96), .B (n_16_92), .C1 (n_17_93), .C2 (n_15_92) );
AOI211_X1 g_14_96 (.ZN (n_14_96), .A (n_13_95), .B (n_14_93), .C1 (n_18_91), .C2 (n_17_91) );
AOI211_X1 g_13_94 (.ZN (n_13_94), .A (n_15_94), .B (n_12_94), .C1 (n_16_92), .C2 (n_19_92) );
AOI211_X1 g_15_93 (.ZN (n_15_93), .A (n_14_96), .B (n_11_96), .C1 (n_14_93), .C2 (n_17_93) );
AOI211_X1 g_17_92 (.ZN (n_17_92), .A (n_13_94), .B (n_13_95), .C1 (n_12_94), .C2 (n_18_91) );
AOI211_X1 g_19_91 (.ZN (n_19_91), .A (n_15_93), .B (n_15_94), .C1 (n_11_96), .C2 (n_16_92) );
AOI211_X1 g_21_90 (.ZN (n_21_90), .A (n_17_92), .B (n_14_96), .C1 (n_13_95), .C2 (n_14_93) );
AOI211_X1 g_23_89 (.ZN (n_23_89), .A (n_19_91), .B (n_13_94), .C1 (n_15_94), .C2 (n_12_94) );
AOI211_X1 g_25_88 (.ZN (n_25_88), .A (n_21_90), .B (n_15_93), .C1 (n_14_96), .C2 (n_11_96) );
AOI211_X1 g_24_90 (.ZN (n_24_90), .A (n_23_89), .B (n_17_92), .C1 (n_13_94), .C2 (n_13_95) );
AOI211_X1 g_26_89 (.ZN (n_26_89), .A (n_25_88), .B (n_19_91), .C1 (n_15_93), .C2 (n_15_94) );
AOI211_X1 g_28_88 (.ZN (n_28_88), .A (n_24_90), .B (n_21_90), .C1 (n_17_92), .C2 (n_14_96) );
AOI211_X1 g_30_87 (.ZN (n_30_87), .A (n_26_89), .B (n_23_89), .C1 (n_19_91), .C2 (n_13_94) );
AOI211_X1 g_32_86 (.ZN (n_32_86), .A (n_28_88), .B (n_25_88), .C1 (n_21_90), .C2 (n_15_93) );
AOI211_X1 g_34_85 (.ZN (n_34_85), .A (n_30_87), .B (n_24_90), .C1 (n_23_89), .C2 (n_17_92) );
AOI211_X1 g_36_84 (.ZN (n_36_84), .A (n_32_86), .B (n_26_89), .C1 (n_25_88), .C2 (n_19_91) );
AOI211_X1 g_38_83 (.ZN (n_38_83), .A (n_34_85), .B (n_28_88), .C1 (n_24_90), .C2 (n_21_90) );
AOI211_X1 g_36_82 (.ZN (n_36_82), .A (n_36_84), .B (n_30_87), .C1 (n_26_89), .C2 (n_23_89) );
AOI211_X1 g_38_81 (.ZN (n_38_81), .A (n_38_83), .B (n_32_86), .C1 (n_28_88), .C2 (n_25_88) );
AOI211_X1 g_40_80 (.ZN (n_40_80), .A (n_36_82), .B (n_34_85), .C1 (n_30_87), .C2 (n_24_90) );
AOI211_X1 g_42_79 (.ZN (n_42_79), .A (n_38_81), .B (n_36_84), .C1 (n_32_86), .C2 (n_26_89) );
AOI211_X1 g_44_80 (.ZN (n_44_80), .A (n_40_80), .B (n_38_83), .C1 (n_34_85), .C2 (n_28_88) );
AOI211_X1 g_42_81 (.ZN (n_42_81), .A (n_42_79), .B (n_36_82), .C1 (n_36_84), .C2 (n_30_87) );
AOI211_X1 g_40_82 (.ZN (n_40_82), .A (n_44_80), .B (n_38_81), .C1 (n_38_83), .C2 (n_32_86) );
AOI211_X1 g_39_84 (.ZN (n_39_84), .A (n_42_81), .B (n_40_80), .C1 (n_36_82), .C2 (n_34_85) );
AOI211_X1 g_37_83 (.ZN (n_37_83), .A (n_40_82), .B (n_42_79), .C1 (n_38_81), .C2 (n_36_84) );
AOI211_X1 g_39_82 (.ZN (n_39_82), .A (n_39_84), .B (n_44_80), .C1 (n_40_80), .C2 (n_38_83) );
AOI211_X1 g_41_81 (.ZN (n_41_81), .A (n_37_83), .B (n_42_81), .C1 (n_42_79), .C2 (n_36_82) );
AOI211_X1 g_43_80 (.ZN (n_43_80), .A (n_39_82), .B (n_40_82), .C1 (n_44_80), .C2 (n_38_81) );
AOI211_X1 g_45_79 (.ZN (n_45_79), .A (n_41_81), .B (n_39_84), .C1 (n_42_81), .C2 (n_40_80) );
AOI211_X1 g_47_78 (.ZN (n_47_78), .A (n_43_80), .B (n_37_83), .C1 (n_40_82), .C2 (n_42_79) );
AOI211_X1 g_49_77 (.ZN (n_49_77), .A (n_45_79), .B (n_39_82), .C1 (n_39_84), .C2 (n_44_80) );
AOI211_X1 g_51_76 (.ZN (n_51_76), .A (n_47_78), .B (n_41_81), .C1 (n_37_83), .C2 (n_42_81) );
AOI211_X1 g_53_75 (.ZN (n_53_75), .A (n_49_77), .B (n_43_80), .C1 (n_39_82), .C2 (n_40_82) );
AOI211_X1 g_52_77 (.ZN (n_52_77), .A (n_51_76), .B (n_45_79), .C1 (n_41_81), .C2 (n_39_84) );
AOI211_X1 g_54_76 (.ZN (n_54_76), .A (n_53_75), .B (n_47_78), .C1 (n_43_80), .C2 (n_37_83) );
AOI211_X1 g_56_75 (.ZN (n_56_75), .A (n_52_77), .B (n_49_77), .C1 (n_45_79), .C2 (n_39_82) );
AOI211_X1 g_58_74 (.ZN (n_58_74), .A (n_54_76), .B (n_51_76), .C1 (n_47_78), .C2 (n_41_81) );
AOI211_X1 g_60_73 (.ZN (n_60_73), .A (n_56_75), .B (n_53_75), .C1 (n_49_77), .C2 (n_43_80) );
AOI211_X1 g_62_72 (.ZN (n_62_72), .A (n_58_74), .B (n_52_77), .C1 (n_51_76), .C2 (n_45_79) );
AOI211_X1 g_64_71 (.ZN (n_64_71), .A (n_60_73), .B (n_54_76), .C1 (n_53_75), .C2 (n_47_78) );
AOI211_X1 g_66_70 (.ZN (n_66_70), .A (n_62_72), .B (n_56_75), .C1 (n_52_77), .C2 (n_49_77) );
AOI211_X1 g_68_69 (.ZN (n_68_69), .A (n_64_71), .B (n_58_74), .C1 (n_54_76), .C2 (n_51_76) );
AOI211_X1 g_70_68 (.ZN (n_70_68), .A (n_66_70), .B (n_60_73), .C1 (n_56_75), .C2 (n_53_75) );
AOI211_X1 g_72_67 (.ZN (n_72_67), .A (n_68_69), .B (n_62_72), .C1 (n_58_74), .C2 (n_52_77) );
AOI211_X1 g_74_66 (.ZN (n_74_66), .A (n_70_68), .B (n_64_71), .C1 (n_60_73), .C2 (n_54_76) );
AOI211_X1 g_76_65 (.ZN (n_76_65), .A (n_72_67), .B (n_66_70), .C1 (n_62_72), .C2 (n_56_75) );
AOI211_X1 g_78_64 (.ZN (n_78_64), .A (n_74_66), .B (n_68_69), .C1 (n_64_71), .C2 (n_58_74) );
AOI211_X1 g_80_63 (.ZN (n_80_63), .A (n_76_65), .B (n_70_68), .C1 (n_66_70), .C2 (n_60_73) );
AOI211_X1 g_82_62 (.ZN (n_82_62), .A (n_78_64), .B (n_72_67), .C1 (n_68_69), .C2 (n_62_72) );
AOI211_X1 g_84_61 (.ZN (n_84_61), .A (n_80_63), .B (n_74_66), .C1 (n_70_68), .C2 (n_64_71) );
AOI211_X1 g_86_60 (.ZN (n_86_60), .A (n_82_62), .B (n_76_65), .C1 (n_72_67), .C2 (n_66_70) );
AOI211_X1 g_88_59 (.ZN (n_88_59), .A (n_84_61), .B (n_78_64), .C1 (n_74_66), .C2 (n_68_69) );
AOI211_X1 g_90_58 (.ZN (n_90_58), .A (n_86_60), .B (n_80_63), .C1 (n_76_65), .C2 (n_70_68) );
AOI211_X1 g_89_60 (.ZN (n_89_60), .A (n_88_59), .B (n_82_62), .C1 (n_78_64), .C2 (n_72_67) );
AOI211_X1 g_91_59 (.ZN (n_91_59), .A (n_90_58), .B (n_84_61), .C1 (n_80_63), .C2 (n_74_66) );
AOI211_X1 g_93_58 (.ZN (n_93_58), .A (n_89_60), .B (n_86_60), .C1 (n_82_62), .C2 (n_76_65) );
AOI211_X1 g_95_57 (.ZN (n_95_57), .A (n_91_59), .B (n_88_59), .C1 (n_84_61), .C2 (n_78_64) );
AOI211_X1 g_97_56 (.ZN (n_97_56), .A (n_93_58), .B (n_90_58), .C1 (n_86_60), .C2 (n_80_63) );
AOI211_X1 g_99_55 (.ZN (n_99_55), .A (n_95_57), .B (n_89_60), .C1 (n_88_59), .C2 (n_82_62) );
AOI211_X1 g_101_54 (.ZN (n_101_54), .A (n_97_56), .B (n_91_59), .C1 (n_90_58), .C2 (n_84_61) );
AOI211_X1 g_103_53 (.ZN (n_103_53), .A (n_99_55), .B (n_93_58), .C1 (n_89_60), .C2 (n_86_60) );
AOI211_X1 g_105_52 (.ZN (n_105_52), .A (n_101_54), .B (n_95_57), .C1 (n_91_59), .C2 (n_88_59) );
AOI211_X1 g_107_51 (.ZN (n_107_51), .A (n_103_53), .B (n_97_56), .C1 (n_93_58), .C2 (n_90_58) );
AOI211_X1 g_109_50 (.ZN (n_109_50), .A (n_105_52), .B (n_99_55), .C1 (n_95_57), .C2 (n_89_60) );
AOI211_X1 g_111_49 (.ZN (n_111_49), .A (n_107_51), .B (n_101_54), .C1 (n_97_56), .C2 (n_91_59) );
AOI211_X1 g_113_48 (.ZN (n_113_48), .A (n_109_50), .B (n_103_53), .C1 (n_99_55), .C2 (n_93_58) );
AOI211_X1 g_115_47 (.ZN (n_115_47), .A (n_111_49), .B (n_105_52), .C1 (n_101_54), .C2 (n_95_57) );
AOI211_X1 g_117_46 (.ZN (n_117_46), .A (n_113_48), .B (n_107_51), .C1 (n_103_53), .C2 (n_97_56) );
AOI211_X1 g_119_45 (.ZN (n_119_45), .A (n_115_47), .B (n_109_50), .C1 (n_105_52), .C2 (n_99_55) );
AOI211_X1 g_121_44 (.ZN (n_121_44), .A (n_117_46), .B (n_111_49), .C1 (n_107_51), .C2 (n_101_54) );
AOI211_X1 g_123_43 (.ZN (n_123_43), .A (n_119_45), .B (n_113_48), .C1 (n_109_50), .C2 (n_103_53) );
AOI211_X1 g_125_42 (.ZN (n_125_42), .A (n_121_44), .B (n_115_47), .C1 (n_111_49), .C2 (n_105_52) );
AOI211_X1 g_127_41 (.ZN (n_127_41), .A (n_123_43), .B (n_117_46), .C1 (n_113_48), .C2 (n_107_51) );
AOI211_X1 g_129_40 (.ZN (n_129_40), .A (n_125_42), .B (n_119_45), .C1 (n_115_47), .C2 (n_109_50) );
AOI211_X1 g_131_39 (.ZN (n_131_39), .A (n_127_41), .B (n_121_44), .C1 (n_117_46), .C2 (n_111_49) );
AOI211_X1 g_133_38 (.ZN (n_133_38), .A (n_129_40), .B (n_123_43), .C1 (n_119_45), .C2 (n_113_48) );
AOI211_X1 g_135_37 (.ZN (n_135_37), .A (n_131_39), .B (n_125_42), .C1 (n_121_44), .C2 (n_115_47) );
AOI211_X1 g_137_36 (.ZN (n_137_36), .A (n_133_38), .B (n_127_41), .C1 (n_123_43), .C2 (n_117_46) );
AOI211_X1 g_139_35 (.ZN (n_139_35), .A (n_135_37), .B (n_129_40), .C1 (n_125_42), .C2 (n_119_45) );
AOI211_X1 g_141_34 (.ZN (n_141_34), .A (n_137_36), .B (n_131_39), .C1 (n_127_41), .C2 (n_121_44) );
AOI211_X1 g_143_33 (.ZN (n_143_33), .A (n_139_35), .B (n_133_38), .C1 (n_129_40), .C2 (n_123_43) );
AOI211_X1 g_145_32 (.ZN (n_145_32), .A (n_141_34), .B (n_135_37), .C1 (n_131_39), .C2 (n_125_42) );
AOI211_X1 g_147_33 (.ZN (n_147_33), .A (n_143_33), .B (n_137_36), .C1 (n_133_38), .C2 (n_127_41) );
AOI211_X1 g_145_34 (.ZN (n_145_34), .A (n_145_32), .B (n_139_35), .C1 (n_135_37), .C2 (n_129_40) );
AOI211_X1 g_143_35 (.ZN (n_143_35), .A (n_147_33), .B (n_141_34), .C1 (n_137_36), .C2 (n_131_39) );
AOI211_X1 g_144_33 (.ZN (n_144_33), .A (n_145_34), .B (n_143_33), .C1 (n_139_35), .C2 (n_133_38) );
AOI211_X1 g_145_35 (.ZN (n_145_35), .A (n_143_35), .B (n_145_32), .C1 (n_141_34), .C2 (n_135_37) );
AOI211_X1 g_147_36 (.ZN (n_147_36), .A (n_144_33), .B (n_147_33), .C1 (n_143_33), .C2 (n_137_36) );
AOI211_X1 g_146_34 (.ZN (n_146_34), .A (n_145_35), .B (n_145_34), .C1 (n_145_32), .C2 (n_139_35) );
AOI211_X1 g_148_35 (.ZN (n_148_35), .A (n_147_36), .B (n_143_35), .C1 (n_147_33), .C2 (n_141_34) );
AOI211_X1 g_149_37 (.ZN (n_149_37), .A (n_146_34), .B (n_144_33), .C1 (n_145_34), .C2 (n_143_33) );
AOI211_X1 g_147_38 (.ZN (n_147_38), .A (n_148_35), .B (n_145_35), .C1 (n_143_35), .C2 (n_145_32) );
AOI211_X1 g_146_36 (.ZN (n_146_36), .A (n_149_37), .B (n_147_36), .C1 (n_144_33), .C2 (n_147_33) );
AOI211_X1 g_144_35 (.ZN (n_144_35), .A (n_147_38), .B (n_146_34), .C1 (n_145_35), .C2 (n_145_34) );
AOI211_X1 g_142_34 (.ZN (n_142_34), .A (n_146_36), .B (n_148_35), .C1 (n_147_36), .C2 (n_143_35) );
AOI211_X1 g_140_35 (.ZN (n_140_35), .A (n_144_35), .B (n_149_37), .C1 (n_146_34), .C2 (n_144_33) );
AOI211_X1 g_138_36 (.ZN (n_138_36), .A (n_142_34), .B (n_147_38), .C1 (n_148_35), .C2 (n_145_35) );
AOI211_X1 g_136_37 (.ZN (n_136_37), .A (n_140_35), .B (n_146_36), .C1 (n_149_37), .C2 (n_147_36) );
AOI211_X1 g_134_38 (.ZN (n_134_38), .A (n_138_36), .B (n_144_35), .C1 (n_147_38), .C2 (n_146_34) );
AOI211_X1 g_132_39 (.ZN (n_132_39), .A (n_136_37), .B (n_142_34), .C1 (n_146_36), .C2 (n_148_35) );
AOI211_X1 g_130_40 (.ZN (n_130_40), .A (n_134_38), .B (n_140_35), .C1 (n_144_35), .C2 (n_149_37) );
AOI211_X1 g_128_41 (.ZN (n_128_41), .A (n_132_39), .B (n_138_36), .C1 (n_142_34), .C2 (n_147_38) );
AOI211_X1 g_126_42 (.ZN (n_126_42), .A (n_130_40), .B (n_136_37), .C1 (n_140_35), .C2 (n_146_36) );
AOI211_X1 g_124_43 (.ZN (n_124_43), .A (n_128_41), .B (n_134_38), .C1 (n_138_36), .C2 (n_144_35) );
AOI211_X1 g_122_44 (.ZN (n_122_44), .A (n_126_42), .B (n_132_39), .C1 (n_136_37), .C2 (n_142_34) );
AOI211_X1 g_120_45 (.ZN (n_120_45), .A (n_124_43), .B (n_130_40), .C1 (n_134_38), .C2 (n_140_35) );
AOI211_X1 g_118_46 (.ZN (n_118_46), .A (n_122_44), .B (n_128_41), .C1 (n_132_39), .C2 (n_138_36) );
AOI211_X1 g_116_47 (.ZN (n_116_47), .A (n_120_45), .B (n_126_42), .C1 (n_130_40), .C2 (n_136_37) );
AOI211_X1 g_114_48 (.ZN (n_114_48), .A (n_118_46), .B (n_124_43), .C1 (n_128_41), .C2 (n_134_38) );
AOI211_X1 g_112_49 (.ZN (n_112_49), .A (n_116_47), .B (n_122_44), .C1 (n_126_42), .C2 (n_132_39) );
AOI211_X1 g_110_50 (.ZN (n_110_50), .A (n_114_48), .B (n_120_45), .C1 (n_124_43), .C2 (n_130_40) );
AOI211_X1 g_111_48 (.ZN (n_111_48), .A (n_112_49), .B (n_118_46), .C1 (n_122_44), .C2 (n_128_41) );
AOI211_X1 g_109_49 (.ZN (n_109_49), .A (n_110_50), .B (n_116_47), .C1 (n_120_45), .C2 (n_126_42) );
AOI211_X1 g_107_50 (.ZN (n_107_50), .A (n_111_48), .B (n_114_48), .C1 (n_118_46), .C2 (n_124_43) );
AOI211_X1 g_105_51 (.ZN (n_105_51), .A (n_109_49), .B (n_112_49), .C1 (n_116_47), .C2 (n_122_44) );
AOI211_X1 g_103_52 (.ZN (n_103_52), .A (n_107_50), .B (n_110_50), .C1 (n_114_48), .C2 (n_120_45) );
AOI211_X1 g_101_53 (.ZN (n_101_53), .A (n_105_51), .B (n_111_48), .C1 (n_112_49), .C2 (n_118_46) );
AOI211_X1 g_99_54 (.ZN (n_99_54), .A (n_103_52), .B (n_109_49), .C1 (n_110_50), .C2 (n_116_47) );
AOI211_X1 g_97_55 (.ZN (n_97_55), .A (n_101_53), .B (n_107_50), .C1 (n_111_48), .C2 (n_114_48) );
AOI211_X1 g_95_56 (.ZN (n_95_56), .A (n_99_54), .B (n_105_51), .C1 (n_109_49), .C2 (n_112_49) );
AOI211_X1 g_93_57 (.ZN (n_93_57), .A (n_97_55), .B (n_103_52), .C1 (n_107_50), .C2 (n_110_50) );
AOI211_X1 g_91_58 (.ZN (n_91_58), .A (n_95_56), .B (n_101_53), .C1 (n_105_51), .C2 (n_111_48) );
AOI211_X1 g_89_59 (.ZN (n_89_59), .A (n_93_57), .B (n_99_54), .C1 (n_103_52), .C2 (n_109_49) );
AOI211_X1 g_87_60 (.ZN (n_87_60), .A (n_91_58), .B (n_97_55), .C1 (n_101_53), .C2 (n_107_50) );
AOI211_X1 g_85_61 (.ZN (n_85_61), .A (n_89_59), .B (n_95_56), .C1 (n_99_54), .C2 (n_105_51) );
AOI211_X1 g_83_62 (.ZN (n_83_62), .A (n_87_60), .B (n_93_57), .C1 (n_97_55), .C2 (n_103_52) );
AOI211_X1 g_81_63 (.ZN (n_81_63), .A (n_85_61), .B (n_91_58), .C1 (n_95_56), .C2 (n_101_53) );
AOI211_X1 g_79_64 (.ZN (n_79_64), .A (n_83_62), .B (n_89_59), .C1 (n_93_57), .C2 (n_99_54) );
AOI211_X1 g_77_65 (.ZN (n_77_65), .A (n_81_63), .B (n_87_60), .C1 (n_91_58), .C2 (n_97_55) );
AOI211_X1 g_75_66 (.ZN (n_75_66), .A (n_79_64), .B (n_85_61), .C1 (n_89_59), .C2 (n_95_56) );
AOI211_X1 g_73_67 (.ZN (n_73_67), .A (n_77_65), .B (n_83_62), .C1 (n_87_60), .C2 (n_93_57) );
AOI211_X1 g_71_68 (.ZN (n_71_68), .A (n_75_66), .B (n_81_63), .C1 (n_85_61), .C2 (n_91_58) );
AOI211_X1 g_69_69 (.ZN (n_69_69), .A (n_73_67), .B (n_79_64), .C1 (n_83_62), .C2 (n_89_59) );
AOI211_X1 g_67_70 (.ZN (n_67_70), .A (n_71_68), .B (n_77_65), .C1 (n_81_63), .C2 (n_87_60) );
AOI211_X1 g_66_72 (.ZN (n_66_72), .A (n_69_69), .B (n_75_66), .C1 (n_79_64), .C2 (n_85_61) );
AOI211_X1 g_65_70 (.ZN (n_65_70), .A (n_67_70), .B (n_73_67), .C1 (n_77_65), .C2 (n_83_62) );
AOI211_X1 g_67_69 (.ZN (n_67_69), .A (n_66_72), .B (n_71_68), .C1 (n_75_66), .C2 (n_81_63) );
AOI211_X1 g_69_68 (.ZN (n_69_68), .A (n_65_70), .B (n_69_69), .C1 (n_73_67), .C2 (n_79_64) );
AOI211_X1 g_71_67 (.ZN (n_71_67), .A (n_67_69), .B (n_67_70), .C1 (n_71_68), .C2 (n_77_65) );
AOI211_X1 g_73_66 (.ZN (n_73_66), .A (n_69_68), .B (n_66_72), .C1 (n_69_69), .C2 (n_75_66) );
AOI211_X1 g_75_65 (.ZN (n_75_65), .A (n_71_67), .B (n_65_70), .C1 (n_67_70), .C2 (n_73_67) );
AOI211_X1 g_77_64 (.ZN (n_77_64), .A (n_73_66), .B (n_67_69), .C1 (n_66_72), .C2 (n_71_68) );
AOI211_X1 g_79_63 (.ZN (n_79_63), .A (n_75_65), .B (n_69_68), .C1 (n_65_70), .C2 (n_69_69) );
AOI211_X1 g_81_62 (.ZN (n_81_62), .A (n_77_64), .B (n_71_67), .C1 (n_67_69), .C2 (n_67_70) );
AOI211_X1 g_83_61 (.ZN (n_83_61), .A (n_79_63), .B (n_73_66), .C1 (n_69_68), .C2 (n_66_72) );
AOI211_X1 g_85_60 (.ZN (n_85_60), .A (n_81_62), .B (n_75_65), .C1 (n_71_67), .C2 (n_65_70) );
AOI211_X1 g_87_61 (.ZN (n_87_61), .A (n_83_61), .B (n_77_64), .C1 (n_73_66), .C2 (n_67_69) );
AOI211_X1 g_85_62 (.ZN (n_85_62), .A (n_85_60), .B (n_79_63), .C1 (n_75_65), .C2 (n_69_68) );
AOI211_X1 g_83_63 (.ZN (n_83_63), .A (n_87_61), .B (n_81_62), .C1 (n_77_64), .C2 (n_71_67) );
AOI211_X1 g_81_64 (.ZN (n_81_64), .A (n_85_62), .B (n_83_61), .C1 (n_79_63), .C2 (n_73_66) );
AOI211_X1 g_79_65 (.ZN (n_79_65), .A (n_83_63), .B (n_85_60), .C1 (n_81_62), .C2 (n_75_65) );
AOI211_X1 g_77_66 (.ZN (n_77_66), .A (n_81_64), .B (n_87_61), .C1 (n_83_61), .C2 (n_77_64) );
AOI211_X1 g_75_67 (.ZN (n_75_67), .A (n_79_65), .B (n_85_62), .C1 (n_85_60), .C2 (n_79_63) );
AOI211_X1 g_73_68 (.ZN (n_73_68), .A (n_77_66), .B (n_83_63), .C1 (n_87_61), .C2 (n_81_62) );
AOI211_X1 g_71_69 (.ZN (n_71_69), .A (n_75_67), .B (n_81_64), .C1 (n_85_62), .C2 (n_83_61) );
AOI211_X1 g_69_70 (.ZN (n_69_70), .A (n_73_68), .B (n_79_65), .C1 (n_83_63), .C2 (n_85_60) );
AOI211_X1 g_67_71 (.ZN (n_67_71), .A (n_71_69), .B (n_77_66), .C1 (n_81_64), .C2 (n_87_61) );
AOI211_X1 g_65_72 (.ZN (n_65_72), .A (n_69_70), .B (n_75_67), .C1 (n_79_65), .C2 (n_85_62) );
AOI211_X1 g_63_71 (.ZN (n_63_71), .A (n_67_71), .B (n_73_68), .C1 (n_77_66), .C2 (n_83_63) );
AOI211_X1 g_61_72 (.ZN (n_61_72), .A (n_65_72), .B (n_71_69), .C1 (n_75_67), .C2 (n_81_64) );
AOI211_X1 g_59_73 (.ZN (n_59_73), .A (n_63_71), .B (n_69_70), .C1 (n_73_68), .C2 (n_79_65) );
AOI211_X1 g_57_74 (.ZN (n_57_74), .A (n_61_72), .B (n_67_71), .C1 (n_71_69), .C2 (n_77_66) );
AOI211_X1 g_55_75 (.ZN (n_55_75), .A (n_59_73), .B (n_65_72), .C1 (n_69_70), .C2 (n_75_67) );
AOI211_X1 g_53_76 (.ZN (n_53_76), .A (n_57_74), .B (n_63_71), .C1 (n_67_71), .C2 (n_73_68) );
AOI211_X1 g_51_77 (.ZN (n_51_77), .A (n_55_75), .B (n_61_72), .C1 (n_65_72), .C2 (n_71_69) );
AOI211_X1 g_49_78 (.ZN (n_49_78), .A (n_53_76), .B (n_59_73), .C1 (n_63_71), .C2 (n_69_70) );
AOI211_X1 g_47_79 (.ZN (n_47_79), .A (n_51_77), .B (n_57_74), .C1 (n_61_72), .C2 (n_67_71) );
AOI211_X1 g_45_80 (.ZN (n_45_80), .A (n_49_78), .B (n_55_75), .C1 (n_59_73), .C2 (n_65_72) );
AOI211_X1 g_43_81 (.ZN (n_43_81), .A (n_47_79), .B (n_53_76), .C1 (n_57_74), .C2 (n_63_71) );
AOI211_X1 g_41_82 (.ZN (n_41_82), .A (n_45_80), .B (n_51_77), .C1 (n_55_75), .C2 (n_61_72) );
AOI211_X1 g_39_83 (.ZN (n_39_83), .A (n_43_81), .B (n_49_78), .C1 (n_53_76), .C2 (n_59_73) );
AOI211_X1 g_37_84 (.ZN (n_37_84), .A (n_41_82), .B (n_47_79), .C1 (n_51_77), .C2 (n_57_74) );
AOI211_X1 g_35_85 (.ZN (n_35_85), .A (n_39_83), .B (n_45_80), .C1 (n_49_78), .C2 (n_55_75) );
AOI211_X1 g_33_86 (.ZN (n_33_86), .A (n_37_84), .B (n_43_81), .C1 (n_47_79), .C2 (n_53_76) );
AOI211_X1 g_31_87 (.ZN (n_31_87), .A (n_35_85), .B (n_41_82), .C1 (n_45_80), .C2 (n_51_77) );
AOI211_X1 g_29_88 (.ZN (n_29_88), .A (n_33_86), .B (n_39_83), .C1 (n_43_81), .C2 (n_49_78) );
AOI211_X1 g_30_86 (.ZN (n_30_86), .A (n_31_87), .B (n_37_84), .C1 (n_41_82), .C2 (n_47_79) );
AOI211_X1 g_28_87 (.ZN (n_28_87), .A (n_29_88), .B (n_35_85), .C1 (n_39_83), .C2 (n_45_80) );
AOI211_X1 g_26_88 (.ZN (n_26_88), .A (n_30_86), .B (n_33_86), .C1 (n_37_84), .C2 (n_43_81) );
AOI211_X1 g_24_89 (.ZN (n_24_89), .A (n_28_87), .B (n_31_87), .C1 (n_35_85), .C2 (n_41_82) );
AOI211_X1 g_22_90 (.ZN (n_22_90), .A (n_26_88), .B (n_29_88), .C1 (n_33_86), .C2 (n_39_83) );
AOI211_X1 g_20_91 (.ZN (n_20_91), .A (n_24_89), .B (n_30_86), .C1 (n_31_87), .C2 (n_37_84) );
AOI211_X1 g_18_92 (.ZN (n_18_92), .A (n_22_90), .B (n_28_87), .C1 (n_29_88), .C2 (n_35_85) );
AOI211_X1 g_16_93 (.ZN (n_16_93), .A (n_20_91), .B (n_26_88), .C1 (n_30_86), .C2 (n_33_86) );
AOI211_X1 g_14_94 (.ZN (n_14_94), .A (n_18_92), .B (n_24_89), .C1 (n_28_87), .C2 (n_31_87) );
AOI211_X1 g_12_95 (.ZN (n_12_95), .A (n_16_93), .B (n_22_90), .C1 (n_26_88), .C2 (n_29_88) );
AOI211_X1 g_10_96 (.ZN (n_10_96), .A (n_14_94), .B (n_20_91), .C1 (n_24_89), .C2 (n_30_86) );
AOI211_X1 g_8_97 (.ZN (n_8_97), .A (n_12_95), .B (n_18_92), .C1 (n_22_90), .C2 (n_28_87) );
AOI211_X1 g_6_98 (.ZN (n_6_98), .A (n_10_96), .B (n_16_93), .C1 (n_20_91), .C2 (n_26_88) );
AOI211_X1 g_8_99 (.ZN (n_8_99), .A (n_8_97), .B (n_14_94), .C1 (n_18_92), .C2 (n_24_89) );
AOI211_X1 g_9_97 (.ZN (n_9_97), .A (n_6_98), .B (n_12_95), .C1 (n_16_93), .C2 (n_22_90) );
AOI211_X1 g_7_98 (.ZN (n_7_98), .A (n_8_99), .B (n_10_96), .C1 (n_14_94), .C2 (n_20_91) );
AOI211_X1 g_5_99 (.ZN (n_5_99), .A (n_9_97), .B (n_8_97), .C1 (n_12_95), .C2 (n_18_92) );
AOI211_X1 g_6_97 (.ZN (n_6_97), .A (n_7_98), .B (n_6_98), .C1 (n_10_96), .C2 (n_16_93) );
AOI211_X1 g_4_98 (.ZN (n_4_98), .A (n_5_99), .B (n_8_99), .C1 (n_8_97), .C2 (n_14_94) );
AOI211_X1 g_3_100 (.ZN (n_3_100), .A (n_6_97), .B (n_9_97), .C1 (n_6_98), .C2 (n_12_95) );
AOI211_X1 g_2_102 (.ZN (n_2_102), .A (n_4_98), .B (n_7_98), .C1 (n_8_99), .C2 (n_10_96) );
AOI211_X1 g_4_101 (.ZN (n_4_101), .A (n_3_100), .B (n_5_99), .C1 (n_9_97), .C2 (n_8_97) );
AOI211_X1 g_3_103 (.ZN (n_3_103), .A (n_2_102), .B (n_6_97), .C1 (n_7_98), .C2 (n_6_98) );
AOI211_X1 g_1_104 (.ZN (n_1_104), .A (n_4_101), .B (n_4_98), .C1 (n_5_99), .C2 (n_8_99) );
AOI211_X1 g_3_105 (.ZN (n_3_105), .A (n_3_103), .B (n_3_100), .C1 (n_6_97), .C2 (n_9_97) );
AOI211_X1 g_4_103 (.ZN (n_4_103), .A (n_1_104), .B (n_2_102), .C1 (n_4_98), .C2 (n_7_98) );
AOI211_X1 g_3_101 (.ZN (n_3_101), .A (n_3_105), .B (n_4_101), .C1 (n_3_100), .C2 (n_5_99) );
AOI211_X1 g_5_102 (.ZN (n_5_102), .A (n_4_103), .B (n_3_103), .C1 (n_2_102), .C2 (n_6_97) );
AOI211_X1 g_7_101 (.ZN (n_7_101), .A (n_3_101), .B (n_1_104), .C1 (n_4_101), .C2 (n_4_98) );
AOI211_X1 g_6_99 (.ZN (n_6_99), .A (n_5_102), .B (n_3_105), .C1 (n_3_103), .C2 (n_3_100) );
AOI211_X1 g_5_101 (.ZN (n_5_101), .A (n_7_101), .B (n_4_103), .C1 (n_1_104), .C2 (n_2_102) );
AOI211_X1 g_7_100 (.ZN (n_7_100), .A (n_6_99), .B (n_3_101), .C1 (n_3_105), .C2 (n_4_101) );
AOI211_X1 g_8_98 (.ZN (n_8_98), .A (n_5_101), .B (n_5_102), .C1 (n_4_103), .C2 (n_3_103) );
AOI211_X1 g_9_96 (.ZN (n_9_96), .A (n_7_100), .B (n_7_101), .C1 (n_3_101), .C2 (n_1_104) );
AOI211_X1 g_11_95 (.ZN (n_11_95), .A (n_8_98), .B (n_6_99), .C1 (n_5_102), .C2 (n_3_105) );
AOI211_X1 g_10_97 (.ZN (n_10_97), .A (n_9_96), .B (n_5_101), .C1 (n_7_101), .C2 (n_4_103) );
AOI211_X1 g_12_96 (.ZN (n_12_96), .A (n_11_95), .B (n_7_100), .C1 (n_6_99), .C2 (n_3_101) );
AOI211_X1 g_14_95 (.ZN (n_14_95), .A (n_10_97), .B (n_8_98), .C1 (n_5_101), .C2 (n_5_102) );
AOI211_X1 g_16_94 (.ZN (n_16_94), .A (n_12_96), .B (n_9_96), .C1 (n_7_100), .C2 (n_7_101) );
AOI211_X1 g_18_93 (.ZN (n_18_93), .A (n_14_95), .B (n_11_95), .C1 (n_8_98), .C2 (n_6_99) );
AOI211_X1 g_20_92 (.ZN (n_20_92), .A (n_16_94), .B (n_10_97), .C1 (n_9_96), .C2 (n_5_101) );
AOI211_X1 g_22_91 (.ZN (n_22_91), .A (n_18_93), .B (n_12_96), .C1 (n_11_95), .C2 (n_7_100) );
AOI211_X1 g_21_93 (.ZN (n_21_93), .A (n_20_92), .B (n_14_95), .C1 (n_10_97), .C2 (n_8_98) );
AOI211_X1 g_23_92 (.ZN (n_23_92), .A (n_22_91), .B (n_16_94), .C1 (n_12_96), .C2 (n_9_96) );
AOI211_X1 g_25_91 (.ZN (n_25_91), .A (n_21_93), .B (n_18_93), .C1 (n_14_95), .C2 (n_11_95) );
AOI211_X1 g_23_90 (.ZN (n_23_90), .A (n_23_92), .B (n_20_92), .C1 (n_16_94), .C2 (n_10_97) );
AOI211_X1 g_25_89 (.ZN (n_25_89), .A (n_25_91), .B (n_22_91), .C1 (n_18_93), .C2 (n_12_96) );
AOI211_X1 g_27_88 (.ZN (n_27_88), .A (n_23_90), .B (n_21_93), .C1 (n_20_92), .C2 (n_14_95) );
AOI211_X1 g_29_87 (.ZN (n_29_87), .A (n_25_89), .B (n_23_92), .C1 (n_22_91), .C2 (n_16_94) );
AOI211_X1 g_31_86 (.ZN (n_31_86), .A (n_27_88), .B (n_25_91), .C1 (n_21_93), .C2 (n_18_93) );
AOI211_X1 g_33_85 (.ZN (n_33_85), .A (n_29_87), .B (n_23_90), .C1 (n_23_92), .C2 (n_20_92) );
AOI211_X1 g_35_84 (.ZN (n_35_84), .A (n_31_86), .B (n_25_89), .C1 (n_25_91), .C2 (n_22_91) );
AOI211_X1 g_37_85 (.ZN (n_37_85), .A (n_33_85), .B (n_27_88), .C1 (n_23_90), .C2 (n_21_93) );
AOI211_X1 g_35_86 (.ZN (n_35_86), .A (n_35_84), .B (n_29_87), .C1 (n_25_89), .C2 (n_23_92) );
AOI211_X1 g_33_87 (.ZN (n_33_87), .A (n_37_85), .B (n_31_86), .C1 (n_27_88), .C2 (n_25_91) );
AOI211_X1 g_31_88 (.ZN (n_31_88), .A (n_35_86), .B (n_33_85), .C1 (n_29_87), .C2 (n_23_90) );
AOI211_X1 g_29_89 (.ZN (n_29_89), .A (n_33_87), .B (n_35_84), .C1 (n_31_86), .C2 (n_25_89) );
AOI211_X1 g_27_90 (.ZN (n_27_90), .A (n_31_88), .B (n_37_85), .C1 (n_33_85), .C2 (n_27_88) );
AOI211_X1 g_26_92 (.ZN (n_26_92), .A (n_29_89), .B (n_35_86), .C1 (n_35_84), .C2 (n_29_87) );
AOI211_X1 g_25_90 (.ZN (n_25_90), .A (n_27_90), .B (n_33_87), .C1 (n_37_85), .C2 (n_31_86) );
AOI211_X1 g_27_89 (.ZN (n_27_89), .A (n_26_92), .B (n_31_88), .C1 (n_35_86), .C2 (n_33_85) );
AOI211_X1 g_26_91 (.ZN (n_26_91), .A (n_25_90), .B (n_29_89), .C1 (n_33_87), .C2 (n_35_84) );
AOI211_X1 g_28_90 (.ZN (n_28_90), .A (n_27_89), .B (n_27_90), .C1 (n_31_88), .C2 (n_37_85) );
AOI211_X1 g_30_89 (.ZN (n_30_89), .A (n_26_91), .B (n_26_92), .C1 (n_29_89), .C2 (n_35_86) );
AOI211_X1 g_32_88 (.ZN (n_32_88), .A (n_28_90), .B (n_25_90), .C1 (n_27_90), .C2 (n_33_87) );
AOI211_X1 g_34_87 (.ZN (n_34_87), .A (n_30_89), .B (n_27_89), .C1 (n_26_92), .C2 (n_31_88) );
AOI211_X1 g_36_86 (.ZN (n_36_86), .A (n_32_88), .B (n_26_91), .C1 (n_25_90), .C2 (n_29_89) );
AOI211_X1 g_38_85 (.ZN (n_38_85), .A (n_34_87), .B (n_28_90), .C1 (n_27_89), .C2 (n_27_90) );
AOI211_X1 g_40_84 (.ZN (n_40_84), .A (n_36_86), .B (n_30_89), .C1 (n_26_91), .C2 (n_26_92) );
AOI211_X1 g_42_83 (.ZN (n_42_83), .A (n_38_85), .B (n_32_88), .C1 (n_28_90), .C2 (n_25_90) );
AOI211_X1 g_44_82 (.ZN (n_44_82), .A (n_40_84), .B (n_34_87), .C1 (n_30_89), .C2 (n_27_89) );
AOI211_X1 g_46_81 (.ZN (n_46_81), .A (n_42_83), .B (n_36_86), .C1 (n_32_88), .C2 (n_26_91) );
AOI211_X1 g_48_80 (.ZN (n_48_80), .A (n_44_82), .B (n_38_85), .C1 (n_34_87), .C2 (n_28_90) );
AOI211_X1 g_50_79 (.ZN (n_50_79), .A (n_46_81), .B (n_40_84), .C1 (n_36_86), .C2 (n_30_89) );
AOI211_X1 g_48_78 (.ZN (n_48_78), .A (n_48_80), .B (n_42_83), .C1 (n_38_85), .C2 (n_32_88) );
AOI211_X1 g_50_77 (.ZN (n_50_77), .A (n_50_79), .B (n_44_82), .C1 (n_40_84), .C2 (n_34_87) );
AOI211_X1 g_52_76 (.ZN (n_52_76), .A (n_48_78), .B (n_46_81), .C1 (n_42_83), .C2 (n_36_86) );
AOI211_X1 g_54_75 (.ZN (n_54_75), .A (n_50_77), .B (n_48_80), .C1 (n_44_82), .C2 (n_38_85) );
AOI211_X1 g_56_74 (.ZN (n_56_74), .A (n_52_76), .B (n_50_79), .C1 (n_46_81), .C2 (n_40_84) );
AOI211_X1 g_58_73 (.ZN (n_58_73), .A (n_54_75), .B (n_48_78), .C1 (n_48_80), .C2 (n_42_83) );
AOI211_X1 g_60_72 (.ZN (n_60_72), .A (n_56_74), .B (n_50_77), .C1 (n_50_79), .C2 (n_44_82) );
AOI211_X1 g_62_71 (.ZN (n_62_71), .A (n_58_73), .B (n_52_76), .C1 (n_48_78), .C2 (n_46_81) );
AOI211_X1 g_61_73 (.ZN (n_61_73), .A (n_60_72), .B (n_54_75), .C1 (n_50_77), .C2 (n_48_80) );
AOI211_X1 g_59_74 (.ZN (n_59_74), .A (n_62_71), .B (n_56_74), .C1 (n_52_76), .C2 (n_50_79) );
AOI211_X1 g_57_75 (.ZN (n_57_75), .A (n_61_73), .B (n_58_73), .C1 (n_54_75), .C2 (n_48_78) );
AOI211_X1 g_55_76 (.ZN (n_55_76), .A (n_59_74), .B (n_60_72), .C1 (n_56_74), .C2 (n_50_77) );
AOI211_X1 g_53_77 (.ZN (n_53_77), .A (n_57_75), .B (n_62_71), .C1 (n_58_73), .C2 (n_52_76) );
AOI211_X1 g_51_78 (.ZN (n_51_78), .A (n_55_76), .B (n_61_73), .C1 (n_60_72), .C2 (n_54_75) );
AOI211_X1 g_49_79 (.ZN (n_49_79), .A (n_53_77), .B (n_59_74), .C1 (n_62_71), .C2 (n_56_74) );
AOI211_X1 g_47_80 (.ZN (n_47_80), .A (n_51_78), .B (n_57_75), .C1 (n_61_73), .C2 (n_58_73) );
AOI211_X1 g_45_81 (.ZN (n_45_81), .A (n_49_79), .B (n_55_76), .C1 (n_59_74), .C2 (n_60_72) );
AOI211_X1 g_43_82 (.ZN (n_43_82), .A (n_47_80), .B (n_53_77), .C1 (n_57_75), .C2 (n_62_71) );
AOI211_X1 g_41_83 (.ZN (n_41_83), .A (n_45_81), .B (n_51_78), .C1 (n_55_76), .C2 (n_61_73) );
AOI211_X1 g_40_85 (.ZN (n_40_85), .A (n_43_82), .B (n_49_79), .C1 (n_53_77), .C2 (n_59_74) );
AOI211_X1 g_38_84 (.ZN (n_38_84), .A (n_41_83), .B (n_47_80), .C1 (n_51_78), .C2 (n_57_75) );
AOI211_X1 g_40_83 (.ZN (n_40_83), .A (n_40_85), .B (n_45_81), .C1 (n_49_79), .C2 (n_55_76) );
AOI211_X1 g_42_82 (.ZN (n_42_82), .A (n_38_84), .B (n_43_82), .C1 (n_47_80), .C2 (n_53_77) );
AOI211_X1 g_44_81 (.ZN (n_44_81), .A (n_40_83), .B (n_41_83), .C1 (n_45_81), .C2 (n_51_78) );
AOI211_X1 g_46_80 (.ZN (n_46_80), .A (n_42_82), .B (n_40_85), .C1 (n_43_82), .C2 (n_49_79) );
AOI211_X1 g_48_79 (.ZN (n_48_79), .A (n_44_81), .B (n_38_84), .C1 (n_41_83), .C2 (n_47_80) );
AOI211_X1 g_50_78 (.ZN (n_50_78), .A (n_46_80), .B (n_40_83), .C1 (n_40_85), .C2 (n_45_81) );
AOI211_X1 g_49_80 (.ZN (n_49_80), .A (n_48_79), .B (n_42_82), .C1 (n_38_84), .C2 (n_43_82) );
AOI211_X1 g_51_79 (.ZN (n_51_79), .A (n_50_78), .B (n_44_81), .C1 (n_40_83), .C2 (n_41_83) );
AOI211_X1 g_53_78 (.ZN (n_53_78), .A (n_49_80), .B (n_46_80), .C1 (n_42_82), .C2 (n_40_85) );
AOI211_X1 g_55_77 (.ZN (n_55_77), .A (n_51_79), .B (n_48_79), .C1 (n_44_81), .C2 (n_38_84) );
AOI211_X1 g_57_76 (.ZN (n_57_76), .A (n_53_78), .B (n_50_78), .C1 (n_46_80), .C2 (n_40_83) );
AOI211_X1 g_59_75 (.ZN (n_59_75), .A (n_55_77), .B (n_49_80), .C1 (n_48_79), .C2 (n_42_82) );
AOI211_X1 g_61_74 (.ZN (n_61_74), .A (n_57_76), .B (n_51_79), .C1 (n_50_78), .C2 (n_44_81) );
AOI211_X1 g_63_73 (.ZN (n_63_73), .A (n_59_75), .B (n_53_78), .C1 (n_49_80), .C2 (n_46_80) );
AOI211_X1 g_62_75 (.ZN (n_62_75), .A (n_61_74), .B (n_55_77), .C1 (n_51_79), .C2 (n_48_79) );
AOI211_X1 g_60_74 (.ZN (n_60_74), .A (n_63_73), .B (n_57_76), .C1 (n_53_78), .C2 (n_50_78) );
AOI211_X1 g_62_73 (.ZN (n_62_73), .A (n_62_75), .B (n_59_75), .C1 (n_55_77), .C2 (n_49_80) );
AOI211_X1 g_64_72 (.ZN (n_64_72), .A (n_60_74), .B (n_61_74), .C1 (n_57_76), .C2 (n_51_79) );
AOI211_X1 g_66_71 (.ZN (n_66_71), .A (n_62_73), .B (n_63_73), .C1 (n_59_75), .C2 (n_53_78) );
AOI211_X1 g_68_70 (.ZN (n_68_70), .A (n_64_72), .B (n_62_75), .C1 (n_61_74), .C2 (n_55_77) );
AOI211_X1 g_70_69 (.ZN (n_70_69), .A (n_66_71), .B (n_60_74), .C1 (n_63_73), .C2 (n_57_76) );
AOI211_X1 g_72_68 (.ZN (n_72_68), .A (n_68_70), .B (n_62_73), .C1 (n_62_75), .C2 (n_59_75) );
AOI211_X1 g_74_67 (.ZN (n_74_67), .A (n_70_69), .B (n_64_72), .C1 (n_60_74), .C2 (n_61_74) );
AOI211_X1 g_76_66 (.ZN (n_76_66), .A (n_72_68), .B (n_66_71), .C1 (n_62_73), .C2 (n_63_73) );
AOI211_X1 g_78_65 (.ZN (n_78_65), .A (n_74_67), .B (n_68_70), .C1 (n_64_72), .C2 (n_62_75) );
AOI211_X1 g_80_64 (.ZN (n_80_64), .A (n_76_66), .B (n_70_69), .C1 (n_66_71), .C2 (n_60_74) );
AOI211_X1 g_82_63 (.ZN (n_82_63), .A (n_78_65), .B (n_72_68), .C1 (n_68_70), .C2 (n_62_73) );
AOI211_X1 g_84_62 (.ZN (n_84_62), .A (n_80_64), .B (n_74_67), .C1 (n_70_69), .C2 (n_64_72) );
AOI211_X1 g_86_61 (.ZN (n_86_61), .A (n_82_63), .B (n_76_66), .C1 (n_72_68), .C2 (n_66_71) );
AOI211_X1 g_88_60 (.ZN (n_88_60), .A (n_84_62), .B (n_78_65), .C1 (n_74_67), .C2 (n_68_70) );
AOI211_X1 g_90_59 (.ZN (n_90_59), .A (n_86_61), .B (n_80_64), .C1 (n_76_66), .C2 (n_70_69) );
AOI211_X1 g_92_58 (.ZN (n_92_58), .A (n_88_60), .B (n_82_63), .C1 (n_78_65), .C2 (n_72_68) );
AOI211_X1 g_94_57 (.ZN (n_94_57), .A (n_90_59), .B (n_84_62), .C1 (n_80_64), .C2 (n_74_67) );
AOI211_X1 g_96_56 (.ZN (n_96_56), .A (n_92_58), .B (n_86_61), .C1 (n_82_63), .C2 (n_76_66) );
AOI211_X1 g_98_55 (.ZN (n_98_55), .A (n_94_57), .B (n_88_60), .C1 (n_84_62), .C2 (n_78_65) );
AOI211_X1 g_100_54 (.ZN (n_100_54), .A (n_96_56), .B (n_90_59), .C1 (n_86_61), .C2 (n_80_64) );
AOI211_X1 g_102_53 (.ZN (n_102_53), .A (n_98_55), .B (n_92_58), .C1 (n_88_60), .C2 (n_82_63) );
AOI211_X1 g_104_52 (.ZN (n_104_52), .A (n_100_54), .B (n_94_57), .C1 (n_90_59), .C2 (n_84_62) );
AOI211_X1 g_106_51 (.ZN (n_106_51), .A (n_102_53), .B (n_96_56), .C1 (n_92_58), .C2 (n_86_61) );
AOI211_X1 g_108_50 (.ZN (n_108_50), .A (n_104_52), .B (n_98_55), .C1 (n_94_57), .C2 (n_88_60) );
AOI211_X1 g_110_49 (.ZN (n_110_49), .A (n_106_51), .B (n_100_54), .C1 (n_96_56), .C2 (n_90_59) );
AOI211_X1 g_112_48 (.ZN (n_112_48), .A (n_108_50), .B (n_102_53), .C1 (n_98_55), .C2 (n_92_58) );
AOI211_X1 g_111_50 (.ZN (n_111_50), .A (n_110_49), .B (n_104_52), .C1 (n_100_54), .C2 (n_94_57) );
AOI211_X1 g_113_49 (.ZN (n_113_49), .A (n_112_48), .B (n_106_51), .C1 (n_102_53), .C2 (n_96_56) );
AOI211_X1 g_115_48 (.ZN (n_115_48), .A (n_111_50), .B (n_108_50), .C1 (n_104_52), .C2 (n_98_55) );
AOI211_X1 g_117_47 (.ZN (n_117_47), .A (n_113_49), .B (n_110_49), .C1 (n_106_51), .C2 (n_100_54) );
AOI211_X1 g_119_46 (.ZN (n_119_46), .A (n_115_48), .B (n_112_48), .C1 (n_108_50), .C2 (n_102_53) );
AOI211_X1 g_120_44 (.ZN (n_120_44), .A (n_117_47), .B (n_111_50), .C1 (n_110_49), .C2 (n_104_52) );
AOI211_X1 g_122_43 (.ZN (n_122_43), .A (n_119_46), .B (n_113_49), .C1 (n_112_48), .C2 (n_106_51) );
AOI211_X1 g_121_45 (.ZN (n_121_45), .A (n_120_44), .B (n_115_48), .C1 (n_111_50), .C2 (n_108_50) );
AOI211_X1 g_120_47 (.ZN (n_120_47), .A (n_122_43), .B (n_117_47), .C1 (n_113_49), .C2 (n_110_49) );
AOI211_X1 g_122_46 (.ZN (n_122_46), .A (n_121_45), .B (n_119_46), .C1 (n_115_48), .C2 (n_112_48) );
AOI211_X1 g_124_45 (.ZN (n_124_45), .A (n_120_47), .B (n_120_44), .C1 (n_117_47), .C2 (n_111_50) );
AOI211_X1 g_126_44 (.ZN (n_126_44), .A (n_122_46), .B (n_122_43), .C1 (n_119_46), .C2 (n_113_49) );
AOI211_X1 g_128_43 (.ZN (n_128_43), .A (n_124_45), .B (n_121_45), .C1 (n_120_44), .C2 (n_115_48) );
AOI211_X1 g_130_42 (.ZN (n_130_42), .A (n_126_44), .B (n_120_47), .C1 (n_122_43), .C2 (n_117_47) );
AOI211_X1 g_132_41 (.ZN (n_132_41), .A (n_128_43), .B (n_122_46), .C1 (n_121_45), .C2 (n_119_46) );
AOI211_X1 g_134_40 (.ZN (n_134_40), .A (n_130_42), .B (n_124_45), .C1 (n_120_47), .C2 (n_120_44) );
AOI211_X1 g_136_39 (.ZN (n_136_39), .A (n_132_41), .B (n_126_44), .C1 (n_122_46), .C2 (n_122_43) );
AOI211_X1 g_138_38 (.ZN (n_138_38), .A (n_134_40), .B (n_128_43), .C1 (n_124_45), .C2 (n_121_45) );
AOI211_X1 g_140_37 (.ZN (n_140_37), .A (n_136_39), .B (n_130_42), .C1 (n_126_44), .C2 (n_120_47) );
AOI211_X1 g_142_36 (.ZN (n_142_36), .A (n_138_38), .B (n_132_41), .C1 (n_128_43), .C2 (n_122_46) );
AOI211_X1 g_144_37 (.ZN (n_144_37), .A (n_140_37), .B (n_134_40), .C1 (n_130_42), .C2 (n_124_45) );
AOI211_X1 g_145_39 (.ZN (n_145_39), .A (n_142_36), .B (n_136_39), .C1 (n_132_41), .C2 (n_126_44) );
AOI211_X1 g_147_40 (.ZN (n_147_40), .A (n_144_37), .B (n_138_38), .C1 (n_134_40), .C2 (n_128_43) );
AOI211_X1 g_149_41 (.ZN (n_149_41), .A (n_145_39), .B (n_140_37), .C1 (n_136_39), .C2 (n_130_42) );
AOI211_X1 g_148_39 (.ZN (n_148_39), .A (n_147_40), .B (n_142_36), .C1 (n_138_38), .C2 (n_132_41) );
AOI211_X1 g_146_38 (.ZN (n_146_38), .A (n_149_41), .B (n_144_37), .C1 (n_140_37), .C2 (n_134_40) );
AOI211_X1 g_145_36 (.ZN (n_145_36), .A (n_148_39), .B (n_145_39), .C1 (n_142_36), .C2 (n_136_39) );
AOI211_X1 g_144_34 (.ZN (n_144_34), .A (n_146_38), .B (n_147_40), .C1 (n_144_37), .C2 (n_138_38) );
AOI211_X1 g_146_35 (.ZN (n_146_35), .A (n_145_36), .B (n_149_41), .C1 (n_145_39), .C2 (n_140_37) );
AOI211_X1 g_147_37 (.ZN (n_147_37), .A (n_144_34), .B (n_148_39), .C1 (n_147_40), .C2 (n_142_36) );
AOI211_X1 g_145_38 (.ZN (n_145_38), .A (n_146_35), .B (n_146_38), .C1 (n_149_41), .C2 (n_144_37) );
AOI211_X1 g_144_36 (.ZN (n_144_36), .A (n_147_37), .B (n_145_36), .C1 (n_148_39), .C2 (n_145_39) );
AOI211_X1 g_142_35 (.ZN (n_142_35), .A (n_145_38), .B (n_144_34), .C1 (n_146_38), .C2 (n_147_40) );
AOI211_X1 g_140_36 (.ZN (n_140_36), .A (n_144_36), .B (n_146_35), .C1 (n_145_36), .C2 (n_149_41) );
AOI211_X1 g_138_37 (.ZN (n_138_37), .A (n_142_35), .B (n_147_37), .C1 (n_144_34), .C2 (n_148_39) );
AOI211_X1 g_136_38 (.ZN (n_136_38), .A (n_140_36), .B (n_145_38), .C1 (n_146_35), .C2 (n_146_38) );
AOI211_X1 g_134_39 (.ZN (n_134_39), .A (n_138_37), .B (n_144_36), .C1 (n_147_37), .C2 (n_145_36) );
AOI211_X1 g_132_40 (.ZN (n_132_40), .A (n_136_38), .B (n_142_35), .C1 (n_145_38), .C2 (n_144_34) );
AOI211_X1 g_130_41 (.ZN (n_130_41), .A (n_134_39), .B (n_140_36), .C1 (n_144_36), .C2 (n_146_35) );
AOI211_X1 g_128_42 (.ZN (n_128_42), .A (n_132_40), .B (n_138_37), .C1 (n_142_35), .C2 (n_147_37) );
AOI211_X1 g_126_43 (.ZN (n_126_43), .A (n_130_41), .B (n_136_38), .C1 (n_140_36), .C2 (n_145_38) );
AOI211_X1 g_124_44 (.ZN (n_124_44), .A (n_128_42), .B (n_134_39), .C1 (n_138_37), .C2 (n_144_36) );
AOI211_X1 g_122_45 (.ZN (n_122_45), .A (n_126_43), .B (n_132_40), .C1 (n_136_38), .C2 (n_142_35) );
AOI211_X1 g_120_46 (.ZN (n_120_46), .A (n_124_44), .B (n_130_41), .C1 (n_134_39), .C2 (n_140_36) );
AOI211_X1 g_118_47 (.ZN (n_118_47), .A (n_122_45), .B (n_128_42), .C1 (n_132_40), .C2 (n_138_37) );
AOI211_X1 g_116_48 (.ZN (n_116_48), .A (n_120_46), .B (n_126_43), .C1 (n_130_41), .C2 (n_136_38) );
AOI211_X1 g_114_49 (.ZN (n_114_49), .A (n_118_47), .B (n_124_44), .C1 (n_128_42), .C2 (n_134_39) );
AOI211_X1 g_112_50 (.ZN (n_112_50), .A (n_116_48), .B (n_122_45), .C1 (n_126_43), .C2 (n_132_40) );
AOI211_X1 g_110_51 (.ZN (n_110_51), .A (n_114_49), .B (n_120_46), .C1 (n_124_44), .C2 (n_130_41) );
AOI211_X1 g_108_52 (.ZN (n_108_52), .A (n_112_50), .B (n_118_47), .C1 (n_122_45), .C2 (n_128_42) );
AOI211_X1 g_106_53 (.ZN (n_106_53), .A (n_110_51), .B (n_116_48), .C1 (n_120_46), .C2 (n_126_43) );
AOI211_X1 g_104_54 (.ZN (n_104_54), .A (n_108_52), .B (n_114_49), .C1 (n_118_47), .C2 (n_124_44) );
AOI211_X1 g_102_55 (.ZN (n_102_55), .A (n_106_53), .B (n_112_50), .C1 (n_116_48), .C2 (n_122_45) );
AOI211_X1 g_100_56 (.ZN (n_100_56), .A (n_104_54), .B (n_110_51), .C1 (n_114_49), .C2 (n_120_46) );
AOI211_X1 g_98_57 (.ZN (n_98_57), .A (n_102_55), .B (n_108_52), .C1 (n_112_50), .C2 (n_118_47) );
AOI211_X1 g_96_58 (.ZN (n_96_58), .A (n_100_56), .B (n_106_53), .C1 (n_110_51), .C2 (n_116_48) );
AOI211_X1 g_94_59 (.ZN (n_94_59), .A (n_98_57), .B (n_104_54), .C1 (n_108_52), .C2 (n_114_49) );
AOI211_X1 g_92_60 (.ZN (n_92_60), .A (n_96_58), .B (n_102_55), .C1 (n_106_53), .C2 (n_112_50) );
AOI211_X1 g_90_61 (.ZN (n_90_61), .A (n_94_59), .B (n_100_56), .C1 (n_104_54), .C2 (n_110_51) );
AOI211_X1 g_88_62 (.ZN (n_88_62), .A (n_92_60), .B (n_98_57), .C1 (n_102_55), .C2 (n_108_52) );
AOI211_X1 g_86_63 (.ZN (n_86_63), .A (n_90_61), .B (n_96_58), .C1 (n_100_56), .C2 (n_106_53) );
AOI211_X1 g_84_64 (.ZN (n_84_64), .A (n_88_62), .B (n_94_59), .C1 (n_98_57), .C2 (n_104_54) );
AOI211_X1 g_82_65 (.ZN (n_82_65), .A (n_86_63), .B (n_92_60), .C1 (n_96_58), .C2 (n_102_55) );
AOI211_X1 g_80_66 (.ZN (n_80_66), .A (n_84_64), .B (n_90_61), .C1 (n_94_59), .C2 (n_100_56) );
AOI211_X1 g_78_67 (.ZN (n_78_67), .A (n_82_65), .B (n_88_62), .C1 (n_92_60), .C2 (n_98_57) );
AOI211_X1 g_76_68 (.ZN (n_76_68), .A (n_80_66), .B (n_86_63), .C1 (n_90_61), .C2 (n_96_58) );
AOI211_X1 g_74_69 (.ZN (n_74_69), .A (n_78_67), .B (n_84_64), .C1 (n_88_62), .C2 (n_94_59) );
AOI211_X1 g_72_70 (.ZN (n_72_70), .A (n_76_68), .B (n_82_65), .C1 (n_86_63), .C2 (n_92_60) );
AOI211_X1 g_70_71 (.ZN (n_70_71), .A (n_74_69), .B (n_80_66), .C1 (n_84_64), .C2 (n_90_61) );
AOI211_X1 g_68_72 (.ZN (n_68_72), .A (n_72_70), .B (n_78_67), .C1 (n_82_65), .C2 (n_88_62) );
AOI211_X1 g_66_73 (.ZN (n_66_73), .A (n_70_71), .B (n_76_68), .C1 (n_80_66), .C2 (n_86_63) );
AOI211_X1 g_64_74 (.ZN (n_64_74), .A (n_68_72), .B (n_74_69), .C1 (n_78_67), .C2 (n_84_64) );
AOI211_X1 g_63_76 (.ZN (n_63_76), .A (n_66_73), .B (n_72_70), .C1 (n_76_68), .C2 (n_82_65) );
AOI211_X1 g_62_74 (.ZN (n_62_74), .A (n_64_74), .B (n_70_71), .C1 (n_74_69), .C2 (n_80_66) );
AOI211_X1 g_64_73 (.ZN (n_64_73), .A (n_63_76), .B (n_68_72), .C1 (n_72_70), .C2 (n_78_67) );
AOI211_X1 g_63_75 (.ZN (n_63_75), .A (n_62_74), .B (n_66_73), .C1 (n_70_71), .C2 (n_76_68) );
AOI211_X1 g_65_74 (.ZN (n_65_74), .A (n_64_73), .B (n_64_74), .C1 (n_68_72), .C2 (n_74_69) );
AOI211_X1 g_67_73 (.ZN (n_67_73), .A (n_63_75), .B (n_63_76), .C1 (n_66_73), .C2 (n_72_70) );
AOI211_X1 g_68_71 (.ZN (n_68_71), .A (n_65_74), .B (n_62_74), .C1 (n_64_74), .C2 (n_70_71) );
AOI211_X1 g_70_70 (.ZN (n_70_70), .A (n_67_73), .B (n_64_73), .C1 (n_63_76), .C2 (n_68_72) );
AOI211_X1 g_72_69 (.ZN (n_72_69), .A (n_68_71), .B (n_63_75), .C1 (n_62_74), .C2 (n_66_73) );
AOI211_X1 g_74_68 (.ZN (n_74_68), .A (n_70_70), .B (n_65_74), .C1 (n_64_73), .C2 (n_64_74) );
AOI211_X1 g_76_67 (.ZN (n_76_67), .A (n_72_69), .B (n_67_73), .C1 (n_63_75), .C2 (n_63_76) );
AOI211_X1 g_78_66 (.ZN (n_78_66), .A (n_74_68), .B (n_68_71), .C1 (n_65_74), .C2 (n_62_74) );
AOI211_X1 g_80_65 (.ZN (n_80_65), .A (n_76_67), .B (n_70_70), .C1 (n_67_73), .C2 (n_64_73) );
AOI211_X1 g_82_64 (.ZN (n_82_64), .A (n_78_66), .B (n_72_69), .C1 (n_68_71), .C2 (n_63_75) );
AOI211_X1 g_84_63 (.ZN (n_84_63), .A (n_80_65), .B (n_74_68), .C1 (n_70_70), .C2 (n_65_74) );
AOI211_X1 g_86_62 (.ZN (n_86_62), .A (n_82_64), .B (n_76_67), .C1 (n_72_69), .C2 (n_67_73) );
AOI211_X1 g_88_61 (.ZN (n_88_61), .A (n_84_63), .B (n_78_66), .C1 (n_74_68), .C2 (n_68_71) );
AOI211_X1 g_90_60 (.ZN (n_90_60), .A (n_86_62), .B (n_80_65), .C1 (n_76_67), .C2 (n_70_70) );
AOI211_X1 g_92_59 (.ZN (n_92_59), .A (n_88_61), .B (n_82_64), .C1 (n_78_66), .C2 (n_72_69) );
AOI211_X1 g_94_58 (.ZN (n_94_58), .A (n_90_60), .B (n_84_63), .C1 (n_80_65), .C2 (n_74_68) );
AOI211_X1 g_96_57 (.ZN (n_96_57), .A (n_92_59), .B (n_86_62), .C1 (n_82_64), .C2 (n_76_67) );
AOI211_X1 g_98_56 (.ZN (n_98_56), .A (n_94_58), .B (n_88_61), .C1 (n_84_63), .C2 (n_78_66) );
AOI211_X1 g_100_55 (.ZN (n_100_55), .A (n_96_57), .B (n_90_60), .C1 (n_86_62), .C2 (n_80_65) );
AOI211_X1 g_102_54 (.ZN (n_102_54), .A (n_98_56), .B (n_92_59), .C1 (n_88_61), .C2 (n_82_64) );
AOI211_X1 g_104_53 (.ZN (n_104_53), .A (n_100_55), .B (n_94_58), .C1 (n_90_60), .C2 (n_84_63) );
AOI211_X1 g_106_52 (.ZN (n_106_52), .A (n_102_54), .B (n_96_57), .C1 (n_92_59), .C2 (n_86_62) );
AOI211_X1 g_108_51 (.ZN (n_108_51), .A (n_104_53), .B (n_98_56), .C1 (n_94_58), .C2 (n_88_61) );
AOI211_X1 g_107_53 (.ZN (n_107_53), .A (n_106_52), .B (n_100_55), .C1 (n_96_57), .C2 (n_90_60) );
AOI211_X1 g_109_52 (.ZN (n_109_52), .A (n_108_51), .B (n_102_54), .C1 (n_98_56), .C2 (n_92_59) );
AOI211_X1 g_111_51 (.ZN (n_111_51), .A (n_107_53), .B (n_104_53), .C1 (n_100_55), .C2 (n_94_58) );
AOI211_X1 g_113_50 (.ZN (n_113_50), .A (n_109_52), .B (n_106_52), .C1 (n_102_54), .C2 (n_96_57) );
AOI211_X1 g_115_49 (.ZN (n_115_49), .A (n_111_51), .B (n_108_51), .C1 (n_104_53), .C2 (n_98_56) );
AOI211_X1 g_117_48 (.ZN (n_117_48), .A (n_113_50), .B (n_107_53), .C1 (n_106_52), .C2 (n_100_55) );
AOI211_X1 g_119_47 (.ZN (n_119_47), .A (n_115_49), .B (n_109_52), .C1 (n_108_51), .C2 (n_102_54) );
AOI211_X1 g_121_46 (.ZN (n_121_46), .A (n_117_48), .B (n_111_51), .C1 (n_107_53), .C2 (n_104_53) );
AOI211_X1 g_123_45 (.ZN (n_123_45), .A (n_119_47), .B (n_113_50), .C1 (n_109_52), .C2 (n_106_52) );
AOI211_X1 g_125_44 (.ZN (n_125_44), .A (n_121_46), .B (n_115_49), .C1 (n_111_51), .C2 (n_108_51) );
AOI211_X1 g_127_43 (.ZN (n_127_43), .A (n_123_45), .B (n_117_48), .C1 (n_113_50), .C2 (n_107_53) );
AOI211_X1 g_129_42 (.ZN (n_129_42), .A (n_125_44), .B (n_119_47), .C1 (n_115_49), .C2 (n_109_52) );
AOI211_X1 g_131_41 (.ZN (n_131_41), .A (n_127_43), .B (n_121_46), .C1 (n_117_48), .C2 (n_111_51) );
AOI211_X1 g_133_40 (.ZN (n_133_40), .A (n_129_42), .B (n_123_45), .C1 (n_119_47), .C2 (n_113_50) );
AOI211_X1 g_135_39 (.ZN (n_135_39), .A (n_131_41), .B (n_125_44), .C1 (n_121_46), .C2 (n_115_49) );
AOI211_X1 g_137_38 (.ZN (n_137_38), .A (n_133_40), .B (n_127_43), .C1 (n_123_45), .C2 (n_117_48) );
AOI211_X1 g_139_37 (.ZN (n_139_37), .A (n_135_39), .B (n_129_42), .C1 (n_125_44), .C2 (n_119_47) );
AOI211_X1 g_141_36 (.ZN (n_141_36), .A (n_137_38), .B (n_131_41), .C1 (n_127_43), .C2 (n_121_46) );
AOI211_X1 g_143_37 (.ZN (n_143_37), .A (n_139_37), .B (n_133_40), .C1 (n_129_42), .C2 (n_123_45) );
AOI211_X1 g_141_38 (.ZN (n_141_38), .A (n_141_36), .B (n_135_39), .C1 (n_131_41), .C2 (n_125_44) );
AOI211_X1 g_139_39 (.ZN (n_139_39), .A (n_143_37), .B (n_137_38), .C1 (n_133_40), .C2 (n_127_43) );
AOI211_X1 g_137_40 (.ZN (n_137_40), .A (n_141_38), .B (n_139_37), .C1 (n_135_39), .C2 (n_129_42) );
AOI211_X1 g_135_41 (.ZN (n_135_41), .A (n_139_39), .B (n_141_36), .C1 (n_137_38), .C2 (n_131_41) );
AOI211_X1 g_133_42 (.ZN (n_133_42), .A (n_137_40), .B (n_143_37), .C1 (n_139_37), .C2 (n_133_40) );
AOI211_X1 g_131_43 (.ZN (n_131_43), .A (n_135_41), .B (n_141_38), .C1 (n_141_36), .C2 (n_135_39) );
AOI211_X1 g_129_44 (.ZN (n_129_44), .A (n_133_42), .B (n_139_39), .C1 (n_143_37), .C2 (n_137_38) );
AOI211_X1 g_127_45 (.ZN (n_127_45), .A (n_131_43), .B (n_137_40), .C1 (n_141_38), .C2 (n_139_37) );
AOI211_X1 g_125_46 (.ZN (n_125_46), .A (n_129_44), .B (n_135_41), .C1 (n_139_39), .C2 (n_141_36) );
AOI211_X1 g_123_47 (.ZN (n_123_47), .A (n_127_45), .B (n_133_42), .C1 (n_137_40), .C2 (n_143_37) );
AOI211_X1 g_121_48 (.ZN (n_121_48), .A (n_125_46), .B (n_131_43), .C1 (n_135_41), .C2 (n_141_38) );
AOI211_X1 g_119_49 (.ZN (n_119_49), .A (n_123_47), .B (n_129_44), .C1 (n_133_42), .C2 (n_139_39) );
AOI211_X1 g_117_50 (.ZN (n_117_50), .A (n_121_48), .B (n_127_45), .C1 (n_131_43), .C2 (n_137_40) );
AOI211_X1 g_118_48 (.ZN (n_118_48), .A (n_119_49), .B (n_125_46), .C1 (n_129_44), .C2 (n_135_41) );
AOI211_X1 g_116_49 (.ZN (n_116_49), .A (n_117_50), .B (n_123_47), .C1 (n_127_45), .C2 (n_133_42) );
AOI211_X1 g_114_50 (.ZN (n_114_50), .A (n_118_48), .B (n_121_48), .C1 (n_125_46), .C2 (n_131_43) );
AOI211_X1 g_112_51 (.ZN (n_112_51), .A (n_116_49), .B (n_119_49), .C1 (n_123_47), .C2 (n_129_44) );
AOI211_X1 g_110_52 (.ZN (n_110_52), .A (n_114_50), .B (n_117_50), .C1 (n_121_48), .C2 (n_127_45) );
AOI211_X1 g_108_53 (.ZN (n_108_53), .A (n_112_51), .B (n_118_48), .C1 (n_119_49), .C2 (n_125_46) );
AOI211_X1 g_109_51 (.ZN (n_109_51), .A (n_110_52), .B (n_116_49), .C1 (n_117_50), .C2 (n_123_47) );
AOI211_X1 g_107_52 (.ZN (n_107_52), .A (n_108_53), .B (n_114_50), .C1 (n_118_48), .C2 (n_121_48) );
AOI211_X1 g_105_53 (.ZN (n_105_53), .A (n_109_51), .B (n_112_51), .C1 (n_116_49), .C2 (n_119_49) );
AOI211_X1 g_103_54 (.ZN (n_103_54), .A (n_107_52), .B (n_110_52), .C1 (n_114_50), .C2 (n_117_50) );
AOI211_X1 g_101_55 (.ZN (n_101_55), .A (n_105_53), .B (n_108_53), .C1 (n_112_51), .C2 (n_118_48) );
AOI211_X1 g_99_56 (.ZN (n_99_56), .A (n_103_54), .B (n_109_51), .C1 (n_110_52), .C2 (n_116_49) );
AOI211_X1 g_97_57 (.ZN (n_97_57), .A (n_101_55), .B (n_107_52), .C1 (n_108_53), .C2 (n_114_50) );
AOI211_X1 g_95_58 (.ZN (n_95_58), .A (n_99_56), .B (n_105_53), .C1 (n_109_51), .C2 (n_112_51) );
AOI211_X1 g_93_59 (.ZN (n_93_59), .A (n_97_57), .B (n_103_54), .C1 (n_107_52), .C2 (n_110_52) );
AOI211_X1 g_91_60 (.ZN (n_91_60), .A (n_95_58), .B (n_101_55), .C1 (n_105_53), .C2 (n_108_53) );
AOI211_X1 g_89_61 (.ZN (n_89_61), .A (n_93_59), .B (n_99_56), .C1 (n_103_54), .C2 (n_109_51) );
AOI211_X1 g_87_62 (.ZN (n_87_62), .A (n_91_60), .B (n_97_57), .C1 (n_101_55), .C2 (n_107_52) );
AOI211_X1 g_85_63 (.ZN (n_85_63), .A (n_89_61), .B (n_95_58), .C1 (n_99_56), .C2 (n_105_53) );
AOI211_X1 g_83_64 (.ZN (n_83_64), .A (n_87_62), .B (n_93_59), .C1 (n_97_57), .C2 (n_103_54) );
AOI211_X1 g_81_65 (.ZN (n_81_65), .A (n_85_63), .B (n_91_60), .C1 (n_95_58), .C2 (n_101_55) );
AOI211_X1 g_79_66 (.ZN (n_79_66), .A (n_83_64), .B (n_89_61), .C1 (n_93_59), .C2 (n_99_56) );
AOI211_X1 g_77_67 (.ZN (n_77_67), .A (n_81_65), .B (n_87_62), .C1 (n_91_60), .C2 (n_97_57) );
AOI211_X1 g_75_68 (.ZN (n_75_68), .A (n_79_66), .B (n_85_63), .C1 (n_89_61), .C2 (n_95_58) );
AOI211_X1 g_73_69 (.ZN (n_73_69), .A (n_77_67), .B (n_83_64), .C1 (n_87_62), .C2 (n_93_59) );
AOI211_X1 g_71_70 (.ZN (n_71_70), .A (n_75_68), .B (n_81_65), .C1 (n_85_63), .C2 (n_91_60) );
AOI211_X1 g_69_71 (.ZN (n_69_71), .A (n_73_69), .B (n_79_66), .C1 (n_83_64), .C2 (n_89_61) );
AOI211_X1 g_67_72 (.ZN (n_67_72), .A (n_71_70), .B (n_77_67), .C1 (n_81_65), .C2 (n_87_62) );
AOI211_X1 g_65_73 (.ZN (n_65_73), .A (n_69_71), .B (n_75_68), .C1 (n_79_66), .C2 (n_85_63) );
AOI211_X1 g_63_74 (.ZN (n_63_74), .A (n_67_72), .B (n_73_69), .C1 (n_77_67), .C2 (n_83_64) );
AOI211_X1 g_61_75 (.ZN (n_61_75), .A (n_65_73), .B (n_71_70), .C1 (n_75_68), .C2 (n_81_65) );
AOI211_X1 g_59_76 (.ZN (n_59_76), .A (n_63_74), .B (n_69_71), .C1 (n_73_69), .C2 (n_79_66) );
AOI211_X1 g_57_77 (.ZN (n_57_77), .A (n_61_75), .B (n_67_72), .C1 (n_71_70), .C2 (n_77_67) );
AOI211_X1 g_58_75 (.ZN (n_58_75), .A (n_59_76), .B (n_65_73), .C1 (n_69_71), .C2 (n_75_68) );
AOI211_X1 g_56_76 (.ZN (n_56_76), .A (n_57_77), .B (n_63_74), .C1 (n_67_72), .C2 (n_73_69) );
AOI211_X1 g_54_77 (.ZN (n_54_77), .A (n_58_75), .B (n_61_75), .C1 (n_65_73), .C2 (n_71_70) );
AOI211_X1 g_52_78 (.ZN (n_52_78), .A (n_56_76), .B (n_59_76), .C1 (n_63_74), .C2 (n_69_71) );
AOI211_X1 g_51_80 (.ZN (n_51_80), .A (n_54_77), .B (n_57_77), .C1 (n_61_75), .C2 (n_67_72) );
AOI211_X1 g_53_79 (.ZN (n_53_79), .A (n_52_78), .B (n_58_75), .C1 (n_59_76), .C2 (n_65_73) );
AOI211_X1 g_55_78 (.ZN (n_55_78), .A (n_51_80), .B (n_56_76), .C1 (n_57_77), .C2 (n_63_74) );
AOI211_X1 g_54_80 (.ZN (n_54_80), .A (n_53_79), .B (n_54_77), .C1 (n_58_75), .C2 (n_61_75) );
AOI211_X1 g_52_79 (.ZN (n_52_79), .A (n_55_78), .B (n_52_78), .C1 (n_56_76), .C2 (n_59_76) );
AOI211_X1 g_54_78 (.ZN (n_54_78), .A (n_54_80), .B (n_51_80), .C1 (n_54_77), .C2 (n_57_77) );
AOI211_X1 g_56_77 (.ZN (n_56_77), .A (n_52_79), .B (n_53_79), .C1 (n_52_78), .C2 (n_58_75) );
AOI211_X1 g_58_76 (.ZN (n_58_76), .A (n_54_78), .B (n_55_78), .C1 (n_51_80), .C2 (n_56_76) );
AOI211_X1 g_60_75 (.ZN (n_60_75), .A (n_56_77), .B (n_54_80), .C1 (n_53_79), .C2 (n_54_77) );
AOI211_X1 g_61_77 (.ZN (n_61_77), .A (n_58_76), .B (n_52_79), .C1 (n_55_78), .C2 (n_52_78) );
AOI211_X1 g_59_78 (.ZN (n_59_78), .A (n_60_75), .B (n_54_78), .C1 (n_54_80), .C2 (n_51_80) );
AOI211_X1 g_60_76 (.ZN (n_60_76), .A (n_61_77), .B (n_56_77), .C1 (n_52_79), .C2 (n_53_79) );
AOI211_X1 g_58_77 (.ZN (n_58_77), .A (n_59_78), .B (n_58_76), .C1 (n_54_78), .C2 (n_55_78) );
AOI211_X1 g_56_78 (.ZN (n_56_78), .A (n_60_76), .B (n_60_75), .C1 (n_56_77), .C2 (n_54_80) );
AOI211_X1 g_54_79 (.ZN (n_54_79), .A (n_58_77), .B (n_61_77), .C1 (n_58_76), .C2 (n_52_79) );
AOI211_X1 g_52_80 (.ZN (n_52_80), .A (n_56_78), .B (n_59_78), .C1 (n_60_75), .C2 (n_54_78) );
AOI211_X1 g_50_81 (.ZN (n_50_81), .A (n_54_79), .B (n_60_76), .C1 (n_61_77), .C2 (n_56_77) );
AOI211_X1 g_48_82 (.ZN (n_48_82), .A (n_52_80), .B (n_58_77), .C1 (n_59_78), .C2 (n_58_76) );
AOI211_X1 g_46_83 (.ZN (n_46_83), .A (n_50_81), .B (n_56_78), .C1 (n_60_76), .C2 (n_60_75) );
AOI211_X1 g_47_81 (.ZN (n_47_81), .A (n_48_82), .B (n_54_79), .C1 (n_58_77), .C2 (n_61_77) );
AOI211_X1 g_45_82 (.ZN (n_45_82), .A (n_46_83), .B (n_52_80), .C1 (n_56_78), .C2 (n_59_78) );
AOI211_X1 g_43_83 (.ZN (n_43_83), .A (n_47_81), .B (n_50_81), .C1 (n_54_79), .C2 (n_60_76) );
AOI211_X1 g_41_84 (.ZN (n_41_84), .A (n_45_82), .B (n_48_82), .C1 (n_52_80), .C2 (n_58_77) );
AOI211_X1 g_39_85 (.ZN (n_39_85), .A (n_43_83), .B (n_46_83), .C1 (n_50_81), .C2 (n_56_78) );
AOI211_X1 g_37_86 (.ZN (n_37_86), .A (n_41_84), .B (n_47_81), .C1 (n_48_82), .C2 (n_54_79) );
AOI211_X1 g_35_87 (.ZN (n_35_87), .A (n_39_85), .B (n_45_82), .C1 (n_46_83), .C2 (n_52_80) );
AOI211_X1 g_36_85 (.ZN (n_36_85), .A (n_37_86), .B (n_43_83), .C1 (n_47_81), .C2 (n_50_81) );
AOI211_X1 g_34_86 (.ZN (n_34_86), .A (n_35_87), .B (n_41_84), .C1 (n_45_82), .C2 (n_48_82) );
AOI211_X1 g_32_87 (.ZN (n_32_87), .A (n_36_85), .B (n_39_85), .C1 (n_43_83), .C2 (n_46_83) );
AOI211_X1 g_30_88 (.ZN (n_30_88), .A (n_34_86), .B (n_37_86), .C1 (n_41_84), .C2 (n_47_81) );
AOI211_X1 g_28_89 (.ZN (n_28_89), .A (n_32_87), .B (n_35_87), .C1 (n_39_85), .C2 (n_45_82) );
AOI211_X1 g_26_90 (.ZN (n_26_90), .A (n_30_88), .B (n_36_85), .C1 (n_37_86), .C2 (n_43_83) );
AOI211_X1 g_24_91 (.ZN (n_24_91), .A (n_28_89), .B (n_34_86), .C1 (n_35_87), .C2 (n_41_84) );
AOI211_X1 g_22_92 (.ZN (n_22_92), .A (n_26_90), .B (n_32_87), .C1 (n_36_85), .C2 (n_39_85) );
AOI211_X1 g_20_93 (.ZN (n_20_93), .A (n_24_91), .B (n_30_88), .C1 (n_34_86), .C2 (n_37_86) );
AOI211_X1 g_18_94 (.ZN (n_18_94), .A (n_22_92), .B (n_28_89), .C1 (n_32_87), .C2 (n_35_87) );
AOI211_X1 g_16_95 (.ZN (n_16_95), .A (n_20_93), .B (n_26_90), .C1 (n_30_88), .C2 (n_36_85) );
AOI211_X1 g_15_97 (.ZN (n_15_97), .A (n_18_94), .B (n_24_91), .C1 (n_28_89), .C2 (n_34_86) );
AOI211_X1 g_13_96 (.ZN (n_13_96), .A (n_16_95), .B (n_22_92), .C1 (n_26_90), .C2 (n_32_87) );
AOI211_X1 g_15_95 (.ZN (n_15_95), .A (n_15_97), .B (n_20_93), .C1 (n_24_91), .C2 (n_30_88) );
AOI211_X1 g_17_94 (.ZN (n_17_94), .A (n_13_96), .B (n_18_94), .C1 (n_22_92), .C2 (n_28_89) );
AOI211_X1 g_19_93 (.ZN (n_19_93), .A (n_15_95), .B (n_16_95), .C1 (n_20_93), .C2 (n_26_90) );
AOI211_X1 g_21_92 (.ZN (n_21_92), .A (n_17_94), .B (n_15_97), .C1 (n_18_94), .C2 (n_24_91) );
AOI211_X1 g_23_91 (.ZN (n_23_91), .A (n_19_93), .B (n_13_96), .C1 (n_16_95), .C2 (n_22_92) );
AOI211_X1 g_24_93 (.ZN (n_24_93), .A (n_21_92), .B (n_15_95), .C1 (n_15_97), .C2 (n_20_93) );
AOI211_X1 g_22_94 (.ZN (n_22_94), .A (n_23_91), .B (n_17_94), .C1 (n_13_96), .C2 (n_18_94) );
AOI211_X1 g_20_95 (.ZN (n_20_95), .A (n_24_93), .B (n_19_93), .C1 (n_15_95), .C2 (n_16_95) );
AOI211_X1 g_18_96 (.ZN (n_18_96), .A (n_22_94), .B (n_21_92), .C1 (n_17_94), .C2 (n_15_97) );
AOI211_X1 g_19_94 (.ZN (n_19_94), .A (n_20_95), .B (n_23_91), .C1 (n_19_93), .C2 (n_13_96) );
AOI211_X1 g_17_95 (.ZN (n_17_95), .A (n_18_96), .B (n_24_93), .C1 (n_21_92), .C2 (n_15_95) );
AOI211_X1 g_15_96 (.ZN (n_15_96), .A (n_19_94), .B (n_22_94), .C1 (n_23_91), .C2 (n_17_94) );
AOI211_X1 g_13_97 (.ZN (n_13_97), .A (n_17_95), .B (n_20_95), .C1 (n_24_93), .C2 (n_19_93) );
AOI211_X1 g_11_98 (.ZN (n_11_98), .A (n_15_96), .B (n_18_96), .C1 (n_22_94), .C2 (n_21_92) );
AOI211_X1 g_9_99 (.ZN (n_9_99), .A (n_13_97), .B (n_19_94), .C1 (n_20_95), .C2 (n_23_91) );
AOI211_X1 g_8_101 (.ZN (n_8_101), .A (n_11_98), .B (n_17_95), .C1 (n_18_96), .C2 (n_24_93) );
AOI211_X1 g_7_99 (.ZN (n_7_99), .A (n_9_99), .B (n_15_96), .C1 (n_19_94), .C2 (n_22_94) );
AOI211_X1 g_5_100 (.ZN (n_5_100), .A (n_8_101), .B (n_13_97), .C1 (n_17_95), .C2 (n_20_95) );
AOI211_X1 g_6_102 (.ZN (n_6_102), .A (n_7_99), .B (n_11_98), .C1 (n_15_96), .C2 (n_18_96) );
AOI211_X1 g_5_104 (.ZN (n_5_104), .A (n_5_100), .B (n_9_99), .C1 (n_13_97), .C2 (n_19_94) );
AOI211_X1 g_4_102 (.ZN (n_4_102), .A (n_6_102), .B (n_8_101), .C1 (n_11_98), .C2 (n_17_95) );
AOI211_X1 g_6_101 (.ZN (n_6_101), .A (n_5_104), .B (n_7_99), .C1 (n_9_99), .C2 (n_15_96) );
AOI211_X1 g_7_103 (.ZN (n_7_103), .A (n_4_102), .B (n_5_100), .C1 (n_8_101), .C2 (n_13_97) );
AOI211_X1 g_9_102 (.ZN (n_9_102), .A (n_6_101), .B (n_6_102), .C1 (n_7_99), .C2 (n_11_98) );
AOI211_X1 g_10_100 (.ZN (n_10_100), .A (n_7_103), .B (n_5_104), .C1 (n_5_100), .C2 (n_9_99) );
AOI211_X1 g_9_98 (.ZN (n_9_98), .A (n_9_102), .B (n_4_102), .C1 (n_6_102), .C2 (n_8_101) );
AOI211_X1 g_11_97 (.ZN (n_11_97), .A (n_10_100), .B (n_6_101), .C1 (n_5_104), .C2 (n_7_99) );
AOI211_X1 g_13_98 (.ZN (n_13_98), .A (n_9_98), .B (n_7_103), .C1 (n_4_102), .C2 (n_5_100) );
AOI211_X1 g_11_99 (.ZN (n_11_99), .A (n_11_97), .B (n_9_102), .C1 (n_6_101), .C2 (n_6_102) );
AOI211_X1 g_12_97 (.ZN (n_12_97), .A (n_13_98), .B (n_10_100), .C1 (n_7_103), .C2 (n_5_104) );
AOI211_X1 g_10_98 (.ZN (n_10_98), .A (n_11_99), .B (n_9_98), .C1 (n_9_102), .C2 (n_4_102) );
AOI211_X1 g_9_100 (.ZN (n_9_100), .A (n_12_97), .B (n_11_97), .C1 (n_10_100), .C2 (n_6_101) );
AOI211_X1 g_8_102 (.ZN (n_8_102), .A (n_10_98), .B (n_13_98), .C1 (n_9_98), .C2 (n_7_103) );
AOI211_X1 g_6_103 (.ZN (n_6_103), .A (n_9_100), .B (n_11_99), .C1 (n_11_97), .C2 (n_9_102) );
AOI211_X1 g_5_105 (.ZN (n_5_105), .A (n_8_102), .B (n_12_97), .C1 (n_13_98), .C2 (n_10_100) );
AOI211_X1 g_3_104 (.ZN (n_3_104), .A (n_6_103), .B (n_10_98), .C1 (n_11_99), .C2 (n_9_98) );
AOI211_X1 g_5_103 (.ZN (n_5_103), .A (n_5_105), .B (n_9_100), .C1 (n_12_97), .C2 (n_11_97) );
AOI211_X1 g_7_104 (.ZN (n_7_104), .A (n_3_104), .B (n_8_102), .C1 (n_10_98), .C2 (n_13_98) );
AOI211_X1 g_9_103 (.ZN (n_9_103), .A (n_5_103), .B (n_6_103), .C1 (n_9_100), .C2 (n_11_99) );
AOI211_X1 g_10_101 (.ZN (n_10_101), .A (n_7_104), .B (n_5_105), .C1 (n_8_102), .C2 (n_12_97) );
AOI211_X1 g_8_100 (.ZN (n_8_100), .A (n_9_103), .B (n_3_104), .C1 (n_6_103), .C2 (n_10_98) );
AOI211_X1 g_7_102 (.ZN (n_7_102), .A (n_10_101), .B (n_5_103), .C1 (n_5_105), .C2 (n_9_100) );
AOI211_X1 g_9_101 (.ZN (n_9_101), .A (n_8_100), .B (n_7_104), .C1 (n_3_104), .C2 (n_8_102) );
AOI211_X1 g_10_99 (.ZN (n_10_99), .A (n_7_102), .B (n_9_103), .C1 (n_5_103), .C2 (n_6_103) );
AOI211_X1 g_12_98 (.ZN (n_12_98), .A (n_9_101), .B (n_10_101), .C1 (n_7_104), .C2 (n_5_105) );
AOI211_X1 g_14_97 (.ZN (n_14_97), .A (n_10_99), .B (n_8_100), .C1 (n_9_103), .C2 (n_3_104) );
AOI211_X1 g_16_96 (.ZN (n_16_96), .A (n_12_98), .B (n_7_102), .C1 (n_10_101), .C2 (n_5_103) );
AOI211_X1 g_18_95 (.ZN (n_18_95), .A (n_14_97), .B (n_9_101), .C1 (n_8_100), .C2 (n_7_104) );
AOI211_X1 g_20_94 (.ZN (n_20_94), .A (n_16_96), .B (n_10_99), .C1 (n_7_102), .C2 (n_9_103) );
AOI211_X1 g_22_93 (.ZN (n_22_93), .A (n_18_95), .B (n_12_98), .C1 (n_9_101), .C2 (n_10_101) );
AOI211_X1 g_24_92 (.ZN (n_24_92), .A (n_20_94), .B (n_14_97), .C1 (n_10_99), .C2 (n_8_100) );
AOI211_X1 g_23_94 (.ZN (n_23_94), .A (n_22_93), .B (n_16_96), .C1 (n_12_98), .C2 (n_7_102) );
AOI211_X1 g_25_93 (.ZN (n_25_93), .A (n_24_92), .B (n_18_95), .C1 (n_14_97), .C2 (n_9_101) );
AOI211_X1 g_27_92 (.ZN (n_27_92), .A (n_23_94), .B (n_20_94), .C1 (n_16_96), .C2 (n_10_99) );
AOI211_X1 g_29_91 (.ZN (n_29_91), .A (n_25_93), .B (n_22_93), .C1 (n_18_95), .C2 (n_12_98) );
AOI211_X1 g_31_90 (.ZN (n_31_90), .A (n_27_92), .B (n_24_92), .C1 (n_20_94), .C2 (n_14_97) );
AOI211_X1 g_33_89 (.ZN (n_33_89), .A (n_29_91), .B (n_23_94), .C1 (n_22_93), .C2 (n_16_96) );
AOI211_X1 g_35_88 (.ZN (n_35_88), .A (n_31_90), .B (n_25_93), .C1 (n_24_92), .C2 (n_18_95) );
AOI211_X1 g_37_87 (.ZN (n_37_87), .A (n_33_89), .B (n_27_92), .C1 (n_23_94), .C2 (n_20_94) );
AOI211_X1 g_39_86 (.ZN (n_39_86), .A (n_35_88), .B (n_29_91), .C1 (n_25_93), .C2 (n_22_93) );
AOI211_X1 g_41_85 (.ZN (n_41_85), .A (n_37_87), .B (n_31_90), .C1 (n_27_92), .C2 (n_24_92) );
AOI211_X1 g_43_84 (.ZN (n_43_84), .A (n_39_86), .B (n_33_89), .C1 (n_29_91), .C2 (n_23_94) );
AOI211_X1 g_45_83 (.ZN (n_45_83), .A (n_41_85), .B (n_35_88), .C1 (n_31_90), .C2 (n_25_93) );
AOI211_X1 g_47_82 (.ZN (n_47_82), .A (n_43_84), .B (n_37_87), .C1 (n_33_89), .C2 (n_27_92) );
AOI211_X1 g_49_81 (.ZN (n_49_81), .A (n_45_83), .B (n_39_86), .C1 (n_35_88), .C2 (n_29_91) );
AOI211_X1 g_48_83 (.ZN (n_48_83), .A (n_47_82), .B (n_41_85), .C1 (n_37_87), .C2 (n_31_90) );
AOI211_X1 g_46_82 (.ZN (n_46_82), .A (n_49_81), .B (n_43_84), .C1 (n_39_86), .C2 (n_33_89) );
AOI211_X1 g_48_81 (.ZN (n_48_81), .A (n_48_83), .B (n_45_83), .C1 (n_41_85), .C2 (n_35_88) );
AOI211_X1 g_50_80 (.ZN (n_50_80), .A (n_46_82), .B (n_47_82), .C1 (n_43_84), .C2 (n_37_87) );
AOI211_X1 g_52_81 (.ZN (n_52_81), .A (n_48_81), .B (n_49_81), .C1 (n_45_83), .C2 (n_39_86) );
AOI211_X1 g_50_82 (.ZN (n_50_82), .A (n_50_80), .B (n_48_83), .C1 (n_47_82), .C2 (n_41_85) );
AOI211_X1 g_49_84 (.ZN (n_49_84), .A (n_52_81), .B (n_46_82), .C1 (n_49_81), .C2 (n_43_84) );
AOI211_X1 g_47_83 (.ZN (n_47_83), .A (n_50_82), .B (n_48_81), .C1 (n_48_83), .C2 (n_45_83) );
AOI211_X1 g_49_82 (.ZN (n_49_82), .A (n_49_84), .B (n_50_80), .C1 (n_46_82), .C2 (n_47_82) );
AOI211_X1 g_51_81 (.ZN (n_51_81), .A (n_47_83), .B (n_52_81), .C1 (n_48_81), .C2 (n_49_81) );
AOI211_X1 g_53_80 (.ZN (n_53_80), .A (n_49_82), .B (n_50_82), .C1 (n_50_80), .C2 (n_48_83) );
AOI211_X1 g_55_79 (.ZN (n_55_79), .A (n_51_81), .B (n_49_84), .C1 (n_52_81), .C2 (n_46_82) );
AOI211_X1 g_57_78 (.ZN (n_57_78), .A (n_53_80), .B (n_47_83), .C1 (n_50_82), .C2 (n_48_81) );
AOI211_X1 g_59_77 (.ZN (n_59_77), .A (n_55_79), .B (n_49_82), .C1 (n_49_84), .C2 (n_50_80) );
AOI211_X1 g_61_76 (.ZN (n_61_76), .A (n_57_78), .B (n_51_81), .C1 (n_47_83), .C2 (n_52_81) );
AOI211_X1 g_60_78 (.ZN (n_60_78), .A (n_59_77), .B (n_53_80), .C1 (n_49_82), .C2 (n_50_82) );
AOI211_X1 g_62_77 (.ZN (n_62_77), .A (n_61_76), .B (n_55_79), .C1 (n_51_81), .C2 (n_49_84) );
AOI211_X1 g_64_76 (.ZN (n_64_76), .A (n_60_78), .B (n_57_78), .C1 (n_53_80), .C2 (n_47_83) );
AOI211_X1 g_66_75 (.ZN (n_66_75), .A (n_62_77), .B (n_59_77), .C1 (n_55_79), .C2 (n_49_82) );
AOI211_X1 g_68_74 (.ZN (n_68_74), .A (n_64_76), .B (n_61_76), .C1 (n_57_78), .C2 (n_51_81) );
AOI211_X1 g_69_72 (.ZN (n_69_72), .A (n_66_75), .B (n_60_78), .C1 (n_59_77), .C2 (n_53_80) );
AOI211_X1 g_71_71 (.ZN (n_71_71), .A (n_68_74), .B (n_62_77), .C1 (n_61_76), .C2 (n_55_79) );
AOI211_X1 g_73_70 (.ZN (n_73_70), .A (n_69_72), .B (n_64_76), .C1 (n_60_78), .C2 (n_57_78) );
AOI211_X1 g_75_69 (.ZN (n_75_69), .A (n_71_71), .B (n_66_75), .C1 (n_62_77), .C2 (n_59_77) );
AOI211_X1 g_77_68 (.ZN (n_77_68), .A (n_73_70), .B (n_68_74), .C1 (n_64_76), .C2 (n_61_76) );
AOI211_X1 g_79_67 (.ZN (n_79_67), .A (n_75_69), .B (n_69_72), .C1 (n_66_75), .C2 (n_60_78) );
AOI211_X1 g_81_66 (.ZN (n_81_66), .A (n_77_68), .B (n_71_71), .C1 (n_68_74), .C2 (n_62_77) );
AOI211_X1 g_83_65 (.ZN (n_83_65), .A (n_79_67), .B (n_73_70), .C1 (n_69_72), .C2 (n_64_76) );
AOI211_X1 g_85_64 (.ZN (n_85_64), .A (n_81_66), .B (n_75_69), .C1 (n_71_71), .C2 (n_66_75) );
AOI211_X1 g_87_63 (.ZN (n_87_63), .A (n_83_65), .B (n_77_68), .C1 (n_73_70), .C2 (n_68_74) );
AOI211_X1 g_89_62 (.ZN (n_89_62), .A (n_85_64), .B (n_79_67), .C1 (n_75_69), .C2 (n_69_72) );
AOI211_X1 g_91_61 (.ZN (n_91_61), .A (n_87_63), .B (n_81_66), .C1 (n_77_68), .C2 (n_71_71) );
AOI211_X1 g_93_60 (.ZN (n_93_60), .A (n_89_62), .B (n_83_65), .C1 (n_79_67), .C2 (n_73_70) );
AOI211_X1 g_95_59 (.ZN (n_95_59), .A (n_91_61), .B (n_85_64), .C1 (n_81_66), .C2 (n_75_69) );
AOI211_X1 g_97_58 (.ZN (n_97_58), .A (n_93_60), .B (n_87_63), .C1 (n_83_65), .C2 (n_77_68) );
AOI211_X1 g_99_57 (.ZN (n_99_57), .A (n_95_59), .B (n_89_62), .C1 (n_85_64), .C2 (n_79_67) );
AOI211_X1 g_101_56 (.ZN (n_101_56), .A (n_97_58), .B (n_91_61), .C1 (n_87_63), .C2 (n_81_66) );
AOI211_X1 g_103_55 (.ZN (n_103_55), .A (n_99_57), .B (n_93_60), .C1 (n_89_62), .C2 (n_83_65) );
AOI211_X1 g_105_54 (.ZN (n_105_54), .A (n_101_56), .B (n_95_59), .C1 (n_91_61), .C2 (n_85_64) );
AOI211_X1 g_104_56 (.ZN (n_104_56), .A (n_103_55), .B (n_97_58), .C1 (n_93_60), .C2 (n_87_63) );
AOI211_X1 g_106_55 (.ZN (n_106_55), .A (n_105_54), .B (n_99_57), .C1 (n_95_59), .C2 (n_89_62) );
AOI211_X1 g_108_54 (.ZN (n_108_54), .A (n_104_56), .B (n_101_56), .C1 (n_97_58), .C2 (n_91_61) );
AOI211_X1 g_110_53 (.ZN (n_110_53), .A (n_106_55), .B (n_103_55), .C1 (n_99_57), .C2 (n_93_60) );
AOI211_X1 g_112_52 (.ZN (n_112_52), .A (n_108_54), .B (n_105_54), .C1 (n_101_56), .C2 (n_95_59) );
AOI211_X1 g_114_51 (.ZN (n_114_51), .A (n_110_53), .B (n_104_56), .C1 (n_103_55), .C2 (n_97_58) );
AOI211_X1 g_116_50 (.ZN (n_116_50), .A (n_112_52), .B (n_106_55), .C1 (n_105_54), .C2 (n_99_57) );
AOI211_X1 g_118_49 (.ZN (n_118_49), .A (n_114_51), .B (n_108_54), .C1 (n_104_56), .C2 (n_101_56) );
AOI211_X1 g_120_48 (.ZN (n_120_48), .A (n_116_50), .B (n_110_53), .C1 (n_106_55), .C2 (n_103_55) );
AOI211_X1 g_122_47 (.ZN (n_122_47), .A (n_118_49), .B (n_112_52), .C1 (n_108_54), .C2 (n_105_54) );
AOI211_X1 g_124_46 (.ZN (n_124_46), .A (n_120_48), .B (n_114_51), .C1 (n_110_53), .C2 (n_104_56) );
AOI211_X1 g_126_45 (.ZN (n_126_45), .A (n_122_47), .B (n_116_50), .C1 (n_112_52), .C2 (n_106_55) );
AOI211_X1 g_128_44 (.ZN (n_128_44), .A (n_124_46), .B (n_118_49), .C1 (n_114_51), .C2 (n_108_54) );
AOI211_X1 g_130_43 (.ZN (n_130_43), .A (n_126_45), .B (n_120_48), .C1 (n_116_50), .C2 (n_110_53) );
AOI211_X1 g_132_42 (.ZN (n_132_42), .A (n_128_44), .B (n_122_47), .C1 (n_118_49), .C2 (n_112_52) );
AOI211_X1 g_134_41 (.ZN (n_134_41), .A (n_130_43), .B (n_124_46), .C1 (n_120_48), .C2 (n_114_51) );
AOI211_X1 g_136_40 (.ZN (n_136_40), .A (n_132_42), .B (n_126_45), .C1 (n_122_47), .C2 (n_116_50) );
AOI211_X1 g_138_39 (.ZN (n_138_39), .A (n_134_41), .B (n_128_44), .C1 (n_124_46), .C2 (n_118_49) );
AOI211_X1 g_140_38 (.ZN (n_140_38), .A (n_136_40), .B (n_130_43), .C1 (n_126_45), .C2 (n_120_48) );
AOI211_X1 g_142_37 (.ZN (n_142_37), .A (n_138_39), .B (n_132_42), .C1 (n_128_44), .C2 (n_122_47) );
AOI211_X1 g_143_39 (.ZN (n_143_39), .A (n_140_38), .B (n_134_41), .C1 (n_130_43), .C2 (n_124_46) );
AOI211_X1 g_141_40 (.ZN (n_141_40), .A (n_142_37), .B (n_136_40), .C1 (n_132_42), .C2 (n_126_45) );
AOI211_X1 g_142_38 (.ZN (n_142_38), .A (n_143_39), .B (n_138_39), .C1 (n_134_41), .C2 (n_128_44) );
AOI211_X1 g_143_36 (.ZN (n_143_36), .A (n_141_40), .B (n_140_38), .C1 (n_136_40), .C2 (n_130_43) );
AOI211_X1 g_145_37 (.ZN (n_145_37), .A (n_142_38), .B (n_142_37), .C1 (n_138_39), .C2 (n_132_42) );
AOI211_X1 g_143_38 (.ZN (n_143_38), .A (n_143_36), .B (n_143_39), .C1 (n_140_38), .C2 (n_134_41) );
AOI211_X1 g_141_37 (.ZN (n_141_37), .A (n_145_37), .B (n_141_40), .C1 (n_142_37), .C2 (n_136_40) );
AOI211_X1 g_139_38 (.ZN (n_139_38), .A (n_143_38), .B (n_142_38), .C1 (n_143_39), .C2 (n_138_39) );
AOI211_X1 g_137_39 (.ZN (n_137_39), .A (n_141_37), .B (n_143_36), .C1 (n_141_40), .C2 (n_140_38) );
AOI211_X1 g_135_40 (.ZN (n_135_40), .A (n_139_38), .B (n_145_37), .C1 (n_142_38), .C2 (n_142_37) );
AOI211_X1 g_133_41 (.ZN (n_133_41), .A (n_137_39), .B (n_143_38), .C1 (n_143_36), .C2 (n_143_39) );
AOI211_X1 g_131_42 (.ZN (n_131_42), .A (n_135_40), .B (n_141_37), .C1 (n_145_37), .C2 (n_141_40) );
AOI211_X1 g_129_43 (.ZN (n_129_43), .A (n_133_41), .B (n_139_38), .C1 (n_143_38), .C2 (n_142_38) );
AOI211_X1 g_127_44 (.ZN (n_127_44), .A (n_131_42), .B (n_137_39), .C1 (n_141_37), .C2 (n_143_36) );
AOI211_X1 g_125_45 (.ZN (n_125_45), .A (n_129_43), .B (n_135_40), .C1 (n_139_38), .C2 (n_145_37) );
AOI211_X1 g_123_46 (.ZN (n_123_46), .A (n_127_44), .B (n_133_41), .C1 (n_137_39), .C2 (n_143_38) );
AOI211_X1 g_121_47 (.ZN (n_121_47), .A (n_125_45), .B (n_131_42), .C1 (n_135_40), .C2 (n_141_37) );
AOI211_X1 g_119_48 (.ZN (n_119_48), .A (n_123_46), .B (n_129_43), .C1 (n_133_41), .C2 (n_139_38) );
AOI211_X1 g_117_49 (.ZN (n_117_49), .A (n_121_47), .B (n_127_44), .C1 (n_131_42), .C2 (n_137_39) );
AOI211_X1 g_115_50 (.ZN (n_115_50), .A (n_119_48), .B (n_125_45), .C1 (n_129_43), .C2 (n_135_40) );
AOI211_X1 g_113_51 (.ZN (n_113_51), .A (n_117_49), .B (n_123_46), .C1 (n_127_44), .C2 (n_133_41) );
AOI211_X1 g_111_52 (.ZN (n_111_52), .A (n_115_50), .B (n_121_47), .C1 (n_125_45), .C2 (n_131_42) );
AOI211_X1 g_109_53 (.ZN (n_109_53), .A (n_113_51), .B (n_119_48), .C1 (n_123_46), .C2 (n_129_43) );
AOI211_X1 g_107_54 (.ZN (n_107_54), .A (n_111_52), .B (n_117_49), .C1 (n_121_47), .C2 (n_127_44) );
AOI211_X1 g_105_55 (.ZN (n_105_55), .A (n_109_53), .B (n_115_50), .C1 (n_119_48), .C2 (n_125_45) );
AOI211_X1 g_103_56 (.ZN (n_103_56), .A (n_107_54), .B (n_113_51), .C1 (n_117_49), .C2 (n_123_46) );
AOI211_X1 g_101_57 (.ZN (n_101_57), .A (n_105_55), .B (n_111_52), .C1 (n_115_50), .C2 (n_121_47) );
AOI211_X1 g_99_58 (.ZN (n_99_58), .A (n_103_56), .B (n_109_53), .C1 (n_113_51), .C2 (n_119_48) );
AOI211_X1 g_97_59 (.ZN (n_97_59), .A (n_101_57), .B (n_107_54), .C1 (n_111_52), .C2 (n_117_49) );
AOI211_X1 g_95_60 (.ZN (n_95_60), .A (n_99_58), .B (n_105_55), .C1 (n_109_53), .C2 (n_115_50) );
AOI211_X1 g_93_61 (.ZN (n_93_61), .A (n_97_59), .B (n_103_56), .C1 (n_107_54), .C2 (n_113_51) );
AOI211_X1 g_91_62 (.ZN (n_91_62), .A (n_95_60), .B (n_101_57), .C1 (n_105_55), .C2 (n_111_52) );
AOI211_X1 g_89_63 (.ZN (n_89_63), .A (n_93_61), .B (n_99_58), .C1 (n_103_56), .C2 (n_109_53) );
AOI211_X1 g_87_64 (.ZN (n_87_64), .A (n_91_62), .B (n_97_59), .C1 (n_101_57), .C2 (n_107_54) );
AOI211_X1 g_85_65 (.ZN (n_85_65), .A (n_89_63), .B (n_95_60), .C1 (n_99_58), .C2 (n_105_55) );
AOI211_X1 g_83_66 (.ZN (n_83_66), .A (n_87_64), .B (n_93_61), .C1 (n_97_59), .C2 (n_103_56) );
AOI211_X1 g_81_67 (.ZN (n_81_67), .A (n_85_65), .B (n_91_62), .C1 (n_95_60), .C2 (n_101_57) );
AOI211_X1 g_79_68 (.ZN (n_79_68), .A (n_83_66), .B (n_89_63), .C1 (n_93_61), .C2 (n_99_58) );
AOI211_X1 g_77_69 (.ZN (n_77_69), .A (n_81_67), .B (n_87_64), .C1 (n_91_62), .C2 (n_97_59) );
AOI211_X1 g_75_70 (.ZN (n_75_70), .A (n_79_68), .B (n_85_65), .C1 (n_89_63), .C2 (n_95_60) );
AOI211_X1 g_73_71 (.ZN (n_73_71), .A (n_77_69), .B (n_83_66), .C1 (n_87_64), .C2 (n_93_61) );
AOI211_X1 g_71_72 (.ZN (n_71_72), .A (n_75_70), .B (n_81_67), .C1 (n_85_65), .C2 (n_91_62) );
AOI211_X1 g_69_73 (.ZN (n_69_73), .A (n_73_71), .B (n_79_68), .C1 (n_83_66), .C2 (n_89_63) );
AOI211_X1 g_67_74 (.ZN (n_67_74), .A (n_71_72), .B (n_77_69), .C1 (n_81_67), .C2 (n_87_64) );
AOI211_X1 g_65_75 (.ZN (n_65_75), .A (n_69_73), .B (n_75_70), .C1 (n_79_68), .C2 (n_85_65) );
AOI211_X1 g_64_77 (.ZN (n_64_77), .A (n_67_74), .B (n_73_71), .C1 (n_77_69), .C2 (n_83_66) );
AOI211_X1 g_62_76 (.ZN (n_62_76), .A (n_65_75), .B (n_71_72), .C1 (n_75_70), .C2 (n_81_67) );
AOI211_X1 g_64_75 (.ZN (n_64_75), .A (n_64_77), .B (n_69_73), .C1 (n_73_71), .C2 (n_79_68) );
AOI211_X1 g_66_74 (.ZN (n_66_74), .A (n_62_76), .B (n_67_74), .C1 (n_71_72), .C2 (n_77_69) );
AOI211_X1 g_68_73 (.ZN (n_68_73), .A (n_64_75), .B (n_65_75), .C1 (n_69_73), .C2 (n_75_70) );
AOI211_X1 g_70_72 (.ZN (n_70_72), .A (n_66_74), .B (n_64_77), .C1 (n_67_74), .C2 (n_73_71) );
AOI211_X1 g_72_71 (.ZN (n_72_71), .A (n_68_73), .B (n_62_76), .C1 (n_65_75), .C2 (n_71_72) );
AOI211_X1 g_74_70 (.ZN (n_74_70), .A (n_70_72), .B (n_64_75), .C1 (n_64_77), .C2 (n_69_73) );
AOI211_X1 g_76_69 (.ZN (n_76_69), .A (n_72_71), .B (n_66_74), .C1 (n_62_76), .C2 (n_67_74) );
AOI211_X1 g_78_68 (.ZN (n_78_68), .A (n_74_70), .B (n_68_73), .C1 (n_64_75), .C2 (n_65_75) );
AOI211_X1 g_80_67 (.ZN (n_80_67), .A (n_76_69), .B (n_70_72), .C1 (n_66_74), .C2 (n_64_77) );
AOI211_X1 g_82_66 (.ZN (n_82_66), .A (n_78_68), .B (n_72_71), .C1 (n_68_73), .C2 (n_62_76) );
AOI211_X1 g_84_65 (.ZN (n_84_65), .A (n_80_67), .B (n_74_70), .C1 (n_70_72), .C2 (n_64_75) );
AOI211_X1 g_86_64 (.ZN (n_86_64), .A (n_82_66), .B (n_76_69), .C1 (n_72_71), .C2 (n_66_74) );
AOI211_X1 g_88_63 (.ZN (n_88_63), .A (n_84_65), .B (n_78_68), .C1 (n_74_70), .C2 (n_68_73) );
AOI211_X1 g_90_62 (.ZN (n_90_62), .A (n_86_64), .B (n_80_67), .C1 (n_76_69), .C2 (n_70_72) );
AOI211_X1 g_92_61 (.ZN (n_92_61), .A (n_88_63), .B (n_82_66), .C1 (n_78_68), .C2 (n_72_71) );
AOI211_X1 g_94_60 (.ZN (n_94_60), .A (n_90_62), .B (n_84_65), .C1 (n_80_67), .C2 (n_74_70) );
AOI211_X1 g_96_59 (.ZN (n_96_59), .A (n_92_61), .B (n_86_64), .C1 (n_82_66), .C2 (n_76_69) );
AOI211_X1 g_98_58 (.ZN (n_98_58), .A (n_94_60), .B (n_88_63), .C1 (n_84_65), .C2 (n_78_68) );
AOI211_X1 g_100_57 (.ZN (n_100_57), .A (n_96_59), .B (n_90_62), .C1 (n_86_64), .C2 (n_80_67) );
AOI211_X1 g_102_56 (.ZN (n_102_56), .A (n_98_58), .B (n_92_61), .C1 (n_88_63), .C2 (n_82_66) );
AOI211_X1 g_104_55 (.ZN (n_104_55), .A (n_100_57), .B (n_94_60), .C1 (n_90_62), .C2 (n_84_65) );
AOI211_X1 g_106_54 (.ZN (n_106_54), .A (n_102_56), .B (n_96_59), .C1 (n_92_61), .C2 (n_86_64) );
AOI211_X1 g_105_56 (.ZN (n_105_56), .A (n_104_55), .B (n_98_58), .C1 (n_94_60), .C2 (n_88_63) );
AOI211_X1 g_107_55 (.ZN (n_107_55), .A (n_106_54), .B (n_100_57), .C1 (n_96_59), .C2 (n_90_62) );
AOI211_X1 g_109_54 (.ZN (n_109_54), .A (n_105_56), .B (n_102_56), .C1 (n_98_58), .C2 (n_92_61) );
AOI211_X1 g_111_53 (.ZN (n_111_53), .A (n_107_55), .B (n_104_55), .C1 (n_100_57), .C2 (n_94_60) );
AOI211_X1 g_113_52 (.ZN (n_113_52), .A (n_109_54), .B (n_106_54), .C1 (n_102_56), .C2 (n_96_59) );
AOI211_X1 g_115_51 (.ZN (n_115_51), .A (n_111_53), .B (n_105_56), .C1 (n_104_55), .C2 (n_98_58) );
AOI211_X1 g_114_53 (.ZN (n_114_53), .A (n_113_52), .B (n_107_55), .C1 (n_106_54), .C2 (n_100_57) );
AOI211_X1 g_116_52 (.ZN (n_116_52), .A (n_115_51), .B (n_109_54), .C1 (n_105_56), .C2 (n_102_56) );
AOI211_X1 g_118_51 (.ZN (n_118_51), .A (n_114_53), .B (n_111_53), .C1 (n_107_55), .C2 (n_104_55) );
AOI211_X1 g_120_50 (.ZN (n_120_50), .A (n_116_52), .B (n_113_52), .C1 (n_109_54), .C2 (n_106_54) );
AOI211_X1 g_122_49 (.ZN (n_122_49), .A (n_118_51), .B (n_115_51), .C1 (n_111_53), .C2 (n_105_56) );
AOI211_X1 g_124_48 (.ZN (n_124_48), .A (n_120_50), .B (n_114_53), .C1 (n_113_52), .C2 (n_107_55) );
AOI211_X1 g_126_47 (.ZN (n_126_47), .A (n_122_49), .B (n_116_52), .C1 (n_115_51), .C2 (n_109_54) );
AOI211_X1 g_128_46 (.ZN (n_128_46), .A (n_124_48), .B (n_118_51), .C1 (n_114_53), .C2 (n_111_53) );
AOI211_X1 g_130_45 (.ZN (n_130_45), .A (n_126_47), .B (n_120_50), .C1 (n_116_52), .C2 (n_113_52) );
AOI211_X1 g_132_44 (.ZN (n_132_44), .A (n_128_46), .B (n_122_49), .C1 (n_118_51), .C2 (n_115_51) );
AOI211_X1 g_134_43 (.ZN (n_134_43), .A (n_130_45), .B (n_124_48), .C1 (n_120_50), .C2 (n_114_53) );
AOI211_X1 g_136_42 (.ZN (n_136_42), .A (n_132_44), .B (n_126_47), .C1 (n_122_49), .C2 (n_116_52) );
AOI211_X1 g_138_41 (.ZN (n_138_41), .A (n_134_43), .B (n_128_46), .C1 (n_124_48), .C2 (n_118_51) );
AOI211_X1 g_140_40 (.ZN (n_140_40), .A (n_136_42), .B (n_130_45), .C1 (n_126_47), .C2 (n_120_50) );
AOI211_X1 g_142_39 (.ZN (n_142_39), .A (n_138_41), .B (n_132_44), .C1 (n_128_46), .C2 (n_122_49) );
AOI211_X1 g_144_38 (.ZN (n_144_38), .A (n_140_40), .B (n_134_43), .C1 (n_130_45), .C2 (n_124_48) );
AOI211_X1 g_146_39 (.ZN (n_146_39), .A (n_142_39), .B (n_136_42), .C1 (n_132_44), .C2 (n_126_47) );
AOI211_X1 g_144_40 (.ZN (n_144_40), .A (n_144_38), .B (n_138_41), .C1 (n_134_43), .C2 (n_128_46) );
AOI211_X1 g_142_41 (.ZN (n_142_41), .A (n_146_39), .B (n_140_40), .C1 (n_136_42), .C2 (n_130_45) );
AOI211_X1 g_141_39 (.ZN (n_141_39), .A (n_144_40), .B (n_142_39), .C1 (n_138_41), .C2 (n_132_44) );
AOI211_X1 g_139_40 (.ZN (n_139_40), .A (n_142_41), .B (n_144_38), .C1 (n_140_40), .C2 (n_134_43) );
AOI211_X1 g_137_41 (.ZN (n_137_41), .A (n_141_39), .B (n_146_39), .C1 (n_142_39), .C2 (n_136_42) );
AOI211_X1 g_135_42 (.ZN (n_135_42), .A (n_139_40), .B (n_144_40), .C1 (n_144_38), .C2 (n_138_41) );
AOI211_X1 g_133_43 (.ZN (n_133_43), .A (n_137_41), .B (n_142_41), .C1 (n_146_39), .C2 (n_140_40) );
AOI211_X1 g_131_44 (.ZN (n_131_44), .A (n_135_42), .B (n_141_39), .C1 (n_144_40), .C2 (n_142_39) );
AOI211_X1 g_129_45 (.ZN (n_129_45), .A (n_133_43), .B (n_139_40), .C1 (n_142_41), .C2 (n_144_38) );
AOI211_X1 g_127_46 (.ZN (n_127_46), .A (n_131_44), .B (n_137_41), .C1 (n_141_39), .C2 (n_146_39) );
AOI211_X1 g_125_47 (.ZN (n_125_47), .A (n_129_45), .B (n_135_42), .C1 (n_139_40), .C2 (n_144_40) );
AOI211_X1 g_123_48 (.ZN (n_123_48), .A (n_127_46), .B (n_133_43), .C1 (n_137_41), .C2 (n_142_41) );
AOI211_X1 g_121_49 (.ZN (n_121_49), .A (n_125_47), .B (n_131_44), .C1 (n_135_42), .C2 (n_141_39) );
AOI211_X1 g_119_50 (.ZN (n_119_50), .A (n_123_48), .B (n_129_45), .C1 (n_133_43), .C2 (n_139_40) );
AOI211_X1 g_117_51 (.ZN (n_117_51), .A (n_121_49), .B (n_127_46), .C1 (n_131_44), .C2 (n_137_41) );
AOI211_X1 g_115_52 (.ZN (n_115_52), .A (n_119_50), .B (n_125_47), .C1 (n_129_45), .C2 (n_135_42) );
AOI211_X1 g_113_53 (.ZN (n_113_53), .A (n_117_51), .B (n_123_48), .C1 (n_127_46), .C2 (n_133_43) );
AOI211_X1 g_111_54 (.ZN (n_111_54), .A (n_115_52), .B (n_121_49), .C1 (n_125_47), .C2 (n_131_44) );
AOI211_X1 g_109_55 (.ZN (n_109_55), .A (n_113_53), .B (n_119_50), .C1 (n_123_48), .C2 (n_129_45) );
AOI211_X1 g_107_56 (.ZN (n_107_56), .A (n_111_54), .B (n_117_51), .C1 (n_121_49), .C2 (n_127_46) );
AOI211_X1 g_105_57 (.ZN (n_105_57), .A (n_109_55), .B (n_115_52), .C1 (n_119_50), .C2 (n_125_47) );
AOI211_X1 g_103_58 (.ZN (n_103_58), .A (n_107_56), .B (n_113_53), .C1 (n_117_51), .C2 (n_123_48) );
AOI211_X1 g_101_59 (.ZN (n_101_59), .A (n_105_57), .B (n_111_54), .C1 (n_115_52), .C2 (n_121_49) );
AOI211_X1 g_102_57 (.ZN (n_102_57), .A (n_103_58), .B (n_109_55), .C1 (n_113_53), .C2 (n_119_50) );
AOI211_X1 g_100_58 (.ZN (n_100_58), .A (n_101_59), .B (n_107_56), .C1 (n_111_54), .C2 (n_117_51) );
AOI211_X1 g_98_59 (.ZN (n_98_59), .A (n_102_57), .B (n_105_57), .C1 (n_109_55), .C2 (n_115_52) );
AOI211_X1 g_96_60 (.ZN (n_96_60), .A (n_100_58), .B (n_103_58), .C1 (n_107_56), .C2 (n_113_53) );
AOI211_X1 g_94_61 (.ZN (n_94_61), .A (n_98_59), .B (n_101_59), .C1 (n_105_57), .C2 (n_111_54) );
AOI211_X1 g_92_62 (.ZN (n_92_62), .A (n_96_60), .B (n_102_57), .C1 (n_103_58), .C2 (n_109_55) );
AOI211_X1 g_90_63 (.ZN (n_90_63), .A (n_94_61), .B (n_100_58), .C1 (n_101_59), .C2 (n_107_56) );
AOI211_X1 g_88_64 (.ZN (n_88_64), .A (n_92_62), .B (n_98_59), .C1 (n_102_57), .C2 (n_105_57) );
AOI211_X1 g_86_65 (.ZN (n_86_65), .A (n_90_63), .B (n_96_60), .C1 (n_100_58), .C2 (n_103_58) );
AOI211_X1 g_84_66 (.ZN (n_84_66), .A (n_88_64), .B (n_94_61), .C1 (n_98_59), .C2 (n_101_59) );
AOI211_X1 g_82_67 (.ZN (n_82_67), .A (n_86_65), .B (n_92_62), .C1 (n_96_60), .C2 (n_102_57) );
AOI211_X1 g_80_68 (.ZN (n_80_68), .A (n_84_66), .B (n_90_63), .C1 (n_94_61), .C2 (n_100_58) );
AOI211_X1 g_78_69 (.ZN (n_78_69), .A (n_82_67), .B (n_88_64), .C1 (n_92_62), .C2 (n_98_59) );
AOI211_X1 g_76_70 (.ZN (n_76_70), .A (n_80_68), .B (n_86_65), .C1 (n_90_63), .C2 (n_96_60) );
AOI211_X1 g_74_71 (.ZN (n_74_71), .A (n_78_69), .B (n_84_66), .C1 (n_88_64), .C2 (n_94_61) );
AOI211_X1 g_72_72 (.ZN (n_72_72), .A (n_76_70), .B (n_82_67), .C1 (n_86_65), .C2 (n_92_62) );
AOI211_X1 g_70_73 (.ZN (n_70_73), .A (n_74_71), .B (n_80_68), .C1 (n_84_66), .C2 (n_90_63) );
AOI211_X1 g_69_75 (.ZN (n_69_75), .A (n_72_72), .B (n_78_69), .C1 (n_82_67), .C2 (n_88_64) );
AOI211_X1 g_71_74 (.ZN (n_71_74), .A (n_70_73), .B (n_76_70), .C1 (n_80_68), .C2 (n_86_65) );
AOI211_X1 g_73_73 (.ZN (n_73_73), .A (n_69_75), .B (n_74_71), .C1 (n_78_69), .C2 (n_84_66) );
AOI211_X1 g_75_72 (.ZN (n_75_72), .A (n_71_74), .B (n_72_72), .C1 (n_76_70), .C2 (n_82_67) );
AOI211_X1 g_77_71 (.ZN (n_77_71), .A (n_73_73), .B (n_70_73), .C1 (n_74_71), .C2 (n_80_68) );
AOI211_X1 g_79_70 (.ZN (n_79_70), .A (n_75_72), .B (n_69_75), .C1 (n_72_72), .C2 (n_78_69) );
AOI211_X1 g_81_69 (.ZN (n_81_69), .A (n_77_71), .B (n_71_74), .C1 (n_70_73), .C2 (n_76_70) );
AOI211_X1 g_83_68 (.ZN (n_83_68), .A (n_79_70), .B (n_73_73), .C1 (n_69_75), .C2 (n_74_71) );
AOI211_X1 g_85_67 (.ZN (n_85_67), .A (n_81_69), .B (n_75_72), .C1 (n_71_74), .C2 (n_72_72) );
AOI211_X1 g_87_66 (.ZN (n_87_66), .A (n_83_68), .B (n_77_71), .C1 (n_73_73), .C2 (n_70_73) );
AOI211_X1 g_89_65 (.ZN (n_89_65), .A (n_85_67), .B (n_79_70), .C1 (n_75_72), .C2 (n_69_75) );
AOI211_X1 g_91_64 (.ZN (n_91_64), .A (n_87_66), .B (n_81_69), .C1 (n_77_71), .C2 (n_71_74) );
AOI211_X1 g_93_63 (.ZN (n_93_63), .A (n_89_65), .B (n_83_68), .C1 (n_79_70), .C2 (n_73_73) );
AOI211_X1 g_95_62 (.ZN (n_95_62), .A (n_91_64), .B (n_85_67), .C1 (n_81_69), .C2 (n_75_72) );
AOI211_X1 g_97_61 (.ZN (n_97_61), .A (n_93_63), .B (n_87_66), .C1 (n_83_68), .C2 (n_77_71) );
AOI211_X1 g_99_60 (.ZN (n_99_60), .A (n_95_62), .B (n_89_65), .C1 (n_85_67), .C2 (n_79_70) );
AOI211_X1 g_98_62 (.ZN (n_98_62), .A (n_97_61), .B (n_91_64), .C1 (n_87_66), .C2 (n_81_69) );
AOI211_X1 g_97_60 (.ZN (n_97_60), .A (n_99_60), .B (n_93_63), .C1 (n_89_65), .C2 (n_83_68) );
AOI211_X1 g_99_59 (.ZN (n_99_59), .A (n_98_62), .B (n_95_62), .C1 (n_91_64), .C2 (n_85_67) );
AOI211_X1 g_101_58 (.ZN (n_101_58), .A (n_97_60), .B (n_97_61), .C1 (n_93_63), .C2 (n_87_66) );
AOI211_X1 g_103_57 (.ZN (n_103_57), .A (n_99_59), .B (n_99_60), .C1 (n_95_62), .C2 (n_89_65) );
AOI211_X1 g_102_59 (.ZN (n_102_59), .A (n_101_58), .B (n_98_62), .C1 (n_97_61), .C2 (n_91_64) );
AOI211_X1 g_104_58 (.ZN (n_104_58), .A (n_103_57), .B (n_97_60), .C1 (n_99_60), .C2 (n_93_63) );
AOI211_X1 g_106_57 (.ZN (n_106_57), .A (n_102_59), .B (n_99_59), .C1 (n_98_62), .C2 (n_95_62) );
AOI211_X1 g_108_56 (.ZN (n_108_56), .A (n_104_58), .B (n_101_58), .C1 (n_97_60), .C2 (n_97_61) );
AOI211_X1 g_110_55 (.ZN (n_110_55), .A (n_106_57), .B (n_103_57), .C1 (n_99_59), .C2 (n_99_60) );
AOI211_X1 g_112_54 (.ZN (n_112_54), .A (n_108_56), .B (n_102_59), .C1 (n_101_58), .C2 (n_98_62) );
AOI211_X1 g_111_56 (.ZN (n_111_56), .A (n_110_55), .B (n_104_58), .C1 (n_103_57), .C2 (n_97_60) );
AOI211_X1 g_110_54 (.ZN (n_110_54), .A (n_112_54), .B (n_106_57), .C1 (n_102_59), .C2 (n_99_59) );
AOI211_X1 g_112_53 (.ZN (n_112_53), .A (n_111_56), .B (n_108_56), .C1 (n_104_58), .C2 (n_101_58) );
AOI211_X1 g_114_52 (.ZN (n_114_52), .A (n_110_54), .B (n_110_55), .C1 (n_106_57), .C2 (n_103_57) );
AOI211_X1 g_116_51 (.ZN (n_116_51), .A (n_112_53), .B (n_112_54), .C1 (n_108_56), .C2 (n_102_59) );
AOI211_X1 g_118_50 (.ZN (n_118_50), .A (n_114_52), .B (n_111_56), .C1 (n_110_55), .C2 (n_104_58) );
AOI211_X1 g_120_49 (.ZN (n_120_49), .A (n_116_51), .B (n_110_54), .C1 (n_112_54), .C2 (n_106_57) );
AOI211_X1 g_122_48 (.ZN (n_122_48), .A (n_118_50), .B (n_112_53), .C1 (n_111_56), .C2 (n_108_56) );
AOI211_X1 g_124_47 (.ZN (n_124_47), .A (n_120_49), .B (n_114_52), .C1 (n_110_54), .C2 (n_110_55) );
AOI211_X1 g_126_46 (.ZN (n_126_46), .A (n_122_48), .B (n_116_51), .C1 (n_112_53), .C2 (n_112_54) );
AOI211_X1 g_128_45 (.ZN (n_128_45), .A (n_124_47), .B (n_118_50), .C1 (n_114_52), .C2 (n_111_56) );
AOI211_X1 g_130_44 (.ZN (n_130_44), .A (n_126_46), .B (n_120_49), .C1 (n_116_51), .C2 (n_110_54) );
AOI211_X1 g_132_43 (.ZN (n_132_43), .A (n_128_45), .B (n_122_48), .C1 (n_118_50), .C2 (n_112_53) );
AOI211_X1 g_134_42 (.ZN (n_134_42), .A (n_130_44), .B (n_124_47), .C1 (n_120_49), .C2 (n_114_52) );
AOI211_X1 g_136_41 (.ZN (n_136_41), .A (n_132_43), .B (n_126_46), .C1 (n_122_48), .C2 (n_116_51) );
AOI211_X1 g_138_40 (.ZN (n_138_40), .A (n_134_42), .B (n_128_45), .C1 (n_124_47), .C2 (n_118_50) );
AOI211_X1 g_140_39 (.ZN (n_140_39), .A (n_136_41), .B (n_130_44), .C1 (n_126_46), .C2 (n_120_49) );
AOI211_X1 g_139_41 (.ZN (n_139_41), .A (n_138_40), .B (n_132_43), .C1 (n_128_45), .C2 (n_122_48) );
AOI211_X1 g_137_42 (.ZN (n_137_42), .A (n_140_39), .B (n_134_42), .C1 (n_130_44), .C2 (n_124_47) );
AOI211_X1 g_135_43 (.ZN (n_135_43), .A (n_139_41), .B (n_136_41), .C1 (n_132_43), .C2 (n_126_46) );
AOI211_X1 g_133_44 (.ZN (n_133_44), .A (n_137_42), .B (n_138_40), .C1 (n_134_42), .C2 (n_128_45) );
AOI211_X1 g_131_45 (.ZN (n_131_45), .A (n_135_43), .B (n_140_39), .C1 (n_136_41), .C2 (n_130_44) );
AOI211_X1 g_129_46 (.ZN (n_129_46), .A (n_133_44), .B (n_139_41), .C1 (n_138_40), .C2 (n_132_43) );
AOI211_X1 g_127_47 (.ZN (n_127_47), .A (n_131_45), .B (n_137_42), .C1 (n_140_39), .C2 (n_134_42) );
AOI211_X1 g_125_48 (.ZN (n_125_48), .A (n_129_46), .B (n_135_43), .C1 (n_139_41), .C2 (n_136_41) );
AOI211_X1 g_123_49 (.ZN (n_123_49), .A (n_127_47), .B (n_133_44), .C1 (n_137_42), .C2 (n_138_40) );
AOI211_X1 g_121_50 (.ZN (n_121_50), .A (n_125_48), .B (n_131_45), .C1 (n_135_43), .C2 (n_140_39) );
AOI211_X1 g_119_51 (.ZN (n_119_51), .A (n_123_49), .B (n_129_46), .C1 (n_133_44), .C2 (n_139_41) );
AOI211_X1 g_117_52 (.ZN (n_117_52), .A (n_121_50), .B (n_127_47), .C1 (n_131_45), .C2 (n_137_42) );
AOI211_X1 g_115_53 (.ZN (n_115_53), .A (n_119_51), .B (n_125_48), .C1 (n_129_46), .C2 (n_135_43) );
AOI211_X1 g_113_54 (.ZN (n_113_54), .A (n_117_52), .B (n_123_49), .C1 (n_127_47), .C2 (n_133_44) );
AOI211_X1 g_111_55 (.ZN (n_111_55), .A (n_115_53), .B (n_121_50), .C1 (n_125_48), .C2 (n_131_45) );
AOI211_X1 g_109_56 (.ZN (n_109_56), .A (n_113_54), .B (n_119_51), .C1 (n_123_49), .C2 (n_129_46) );
AOI211_X1 g_107_57 (.ZN (n_107_57), .A (n_111_55), .B (n_117_52), .C1 (n_121_50), .C2 (n_127_47) );
AOI211_X1 g_108_55 (.ZN (n_108_55), .A (n_109_56), .B (n_115_53), .C1 (n_119_51), .C2 (n_125_48) );
AOI211_X1 g_106_56 (.ZN (n_106_56), .A (n_107_57), .B (n_113_54), .C1 (n_117_52), .C2 (n_123_49) );
AOI211_X1 g_104_57 (.ZN (n_104_57), .A (n_108_55), .B (n_111_55), .C1 (n_115_53), .C2 (n_121_50) );
AOI211_X1 g_102_58 (.ZN (n_102_58), .A (n_106_56), .B (n_109_56), .C1 (n_113_54), .C2 (n_119_51) );
AOI211_X1 g_100_59 (.ZN (n_100_59), .A (n_104_57), .B (n_107_57), .C1 (n_111_55), .C2 (n_117_52) );
AOI211_X1 g_98_60 (.ZN (n_98_60), .A (n_102_58), .B (n_108_55), .C1 (n_109_56), .C2 (n_115_53) );
AOI211_X1 g_96_61 (.ZN (n_96_61), .A (n_100_59), .B (n_106_56), .C1 (n_107_57), .C2 (n_113_54) );
AOI211_X1 g_94_62 (.ZN (n_94_62), .A (n_98_60), .B (n_104_57), .C1 (n_108_55), .C2 (n_111_55) );
AOI211_X1 g_92_63 (.ZN (n_92_63), .A (n_96_61), .B (n_102_58), .C1 (n_106_56), .C2 (n_109_56) );
AOI211_X1 g_90_64 (.ZN (n_90_64), .A (n_94_62), .B (n_100_59), .C1 (n_104_57), .C2 (n_107_57) );
AOI211_X1 g_88_65 (.ZN (n_88_65), .A (n_92_63), .B (n_98_60), .C1 (n_102_58), .C2 (n_108_55) );
AOI211_X1 g_86_66 (.ZN (n_86_66), .A (n_90_64), .B (n_96_61), .C1 (n_100_59), .C2 (n_106_56) );
AOI211_X1 g_84_67 (.ZN (n_84_67), .A (n_88_65), .B (n_94_62), .C1 (n_98_60), .C2 (n_104_57) );
AOI211_X1 g_82_68 (.ZN (n_82_68), .A (n_86_66), .B (n_92_63), .C1 (n_96_61), .C2 (n_102_58) );
AOI211_X1 g_80_69 (.ZN (n_80_69), .A (n_84_67), .B (n_90_64), .C1 (n_94_62), .C2 (n_100_59) );
AOI211_X1 g_78_70 (.ZN (n_78_70), .A (n_82_68), .B (n_88_65), .C1 (n_92_63), .C2 (n_98_60) );
AOI211_X1 g_76_71 (.ZN (n_76_71), .A (n_80_69), .B (n_86_66), .C1 (n_90_64), .C2 (n_96_61) );
AOI211_X1 g_74_72 (.ZN (n_74_72), .A (n_78_70), .B (n_84_67), .C1 (n_88_65), .C2 (n_94_62) );
AOI211_X1 g_72_73 (.ZN (n_72_73), .A (n_76_71), .B (n_82_68), .C1 (n_86_66), .C2 (n_92_63) );
AOI211_X1 g_70_74 (.ZN (n_70_74), .A (n_74_72), .B (n_80_69), .C1 (n_84_67), .C2 (n_90_64) );
AOI211_X1 g_68_75 (.ZN (n_68_75), .A (n_72_73), .B (n_78_70), .C1 (n_82_68), .C2 (n_88_65) );
AOI211_X1 g_66_76 (.ZN (n_66_76), .A (n_70_74), .B (n_76_71), .C1 (n_80_69), .C2 (n_86_66) );
AOI211_X1 g_65_78 (.ZN (n_65_78), .A (n_68_75), .B (n_74_72), .C1 (n_78_70), .C2 (n_84_67) );
AOI211_X1 g_63_77 (.ZN (n_63_77), .A (n_66_76), .B (n_72_73), .C1 (n_76_71), .C2 (n_82_68) );
AOI211_X1 g_65_76 (.ZN (n_65_76), .A (n_65_78), .B (n_70_74), .C1 (n_74_72), .C2 (n_80_69) );
AOI211_X1 g_67_75 (.ZN (n_67_75), .A (n_63_77), .B (n_68_75), .C1 (n_72_73), .C2 (n_78_70) );
AOI211_X1 g_69_74 (.ZN (n_69_74), .A (n_65_76), .B (n_66_76), .C1 (n_70_74), .C2 (n_76_71) );
AOI211_X1 g_71_73 (.ZN (n_71_73), .A (n_67_75), .B (n_65_78), .C1 (n_68_75), .C2 (n_74_72) );
AOI211_X1 g_73_72 (.ZN (n_73_72), .A (n_69_74), .B (n_63_77), .C1 (n_66_76), .C2 (n_72_73) );
AOI211_X1 g_75_71 (.ZN (n_75_71), .A (n_71_73), .B (n_65_76), .C1 (n_65_78), .C2 (n_70_74) );
AOI211_X1 g_77_70 (.ZN (n_77_70), .A (n_73_72), .B (n_67_75), .C1 (n_63_77), .C2 (n_68_75) );
AOI211_X1 g_79_69 (.ZN (n_79_69), .A (n_75_71), .B (n_69_74), .C1 (n_65_76), .C2 (n_66_76) );
AOI211_X1 g_81_68 (.ZN (n_81_68), .A (n_77_70), .B (n_71_73), .C1 (n_67_75), .C2 (n_65_78) );
AOI211_X1 g_83_67 (.ZN (n_83_67), .A (n_79_69), .B (n_73_72), .C1 (n_69_74), .C2 (n_63_77) );
AOI211_X1 g_85_66 (.ZN (n_85_66), .A (n_81_68), .B (n_75_71), .C1 (n_71_73), .C2 (n_65_76) );
AOI211_X1 g_87_65 (.ZN (n_87_65), .A (n_83_67), .B (n_77_70), .C1 (n_73_72), .C2 (n_67_75) );
AOI211_X1 g_89_64 (.ZN (n_89_64), .A (n_85_66), .B (n_79_69), .C1 (n_75_71), .C2 (n_69_74) );
AOI211_X1 g_91_63 (.ZN (n_91_63), .A (n_87_65), .B (n_81_68), .C1 (n_77_70), .C2 (n_71_73) );
AOI211_X1 g_93_62 (.ZN (n_93_62), .A (n_89_64), .B (n_83_67), .C1 (n_79_69), .C2 (n_73_72) );
AOI211_X1 g_95_61 (.ZN (n_95_61), .A (n_91_63), .B (n_85_66), .C1 (n_81_68), .C2 (n_75_71) );
AOI211_X1 g_96_63 (.ZN (n_96_63), .A (n_93_62), .B (n_87_65), .C1 (n_83_67), .C2 (n_77_70) );
AOI211_X1 g_94_64 (.ZN (n_94_64), .A (n_95_61), .B (n_89_64), .C1 (n_85_66), .C2 (n_79_69) );
AOI211_X1 g_92_65 (.ZN (n_92_65), .A (n_96_63), .B (n_91_63), .C1 (n_87_65), .C2 (n_81_68) );
AOI211_X1 g_90_66 (.ZN (n_90_66), .A (n_94_64), .B (n_93_62), .C1 (n_89_64), .C2 (n_83_67) );
AOI211_X1 g_88_67 (.ZN (n_88_67), .A (n_92_65), .B (n_95_61), .C1 (n_91_63), .C2 (n_85_66) );
AOI211_X1 g_86_68 (.ZN (n_86_68), .A (n_90_66), .B (n_96_63), .C1 (n_93_62), .C2 (n_87_65) );
AOI211_X1 g_84_69 (.ZN (n_84_69), .A (n_88_67), .B (n_94_64), .C1 (n_95_61), .C2 (n_89_64) );
AOI211_X1 g_82_70 (.ZN (n_82_70), .A (n_86_68), .B (n_92_65), .C1 (n_96_63), .C2 (n_91_63) );
AOI211_X1 g_80_71 (.ZN (n_80_71), .A (n_84_69), .B (n_90_66), .C1 (n_94_64), .C2 (n_93_62) );
AOI211_X1 g_78_72 (.ZN (n_78_72), .A (n_82_70), .B (n_88_67), .C1 (n_92_65), .C2 (n_95_61) );
AOI211_X1 g_76_73 (.ZN (n_76_73), .A (n_80_71), .B (n_86_68), .C1 (n_90_66), .C2 (n_96_63) );
AOI211_X1 g_74_74 (.ZN (n_74_74), .A (n_78_72), .B (n_84_69), .C1 (n_88_67), .C2 (n_94_64) );
AOI211_X1 g_72_75 (.ZN (n_72_75), .A (n_76_73), .B (n_82_70), .C1 (n_86_68), .C2 (n_92_65) );
AOI211_X1 g_70_76 (.ZN (n_70_76), .A (n_74_74), .B (n_80_71), .C1 (n_84_69), .C2 (n_90_66) );
AOI211_X1 g_68_77 (.ZN (n_68_77), .A (n_72_75), .B (n_78_72), .C1 (n_82_70), .C2 (n_88_67) );
AOI211_X1 g_66_78 (.ZN (n_66_78), .A (n_70_76), .B (n_76_73), .C1 (n_80_71), .C2 (n_86_68) );
AOI211_X1 g_67_76 (.ZN (n_67_76), .A (n_68_77), .B (n_74_74), .C1 (n_78_72), .C2 (n_84_69) );
AOI211_X1 g_65_77 (.ZN (n_65_77), .A (n_66_78), .B (n_72_75), .C1 (n_76_73), .C2 (n_82_70) );
AOI211_X1 g_63_78 (.ZN (n_63_78), .A (n_67_76), .B (n_70_76), .C1 (n_74_74), .C2 (n_80_71) );
AOI211_X1 g_61_79 (.ZN (n_61_79), .A (n_65_77), .B (n_68_77), .C1 (n_72_75), .C2 (n_78_72) );
AOI211_X1 g_60_77 (.ZN (n_60_77), .A (n_63_78), .B (n_66_78), .C1 (n_70_76), .C2 (n_76_73) );
AOI211_X1 g_58_78 (.ZN (n_58_78), .A (n_61_79), .B (n_67_76), .C1 (n_68_77), .C2 (n_74_74) );
AOI211_X1 g_56_79 (.ZN (n_56_79), .A (n_60_77), .B (n_65_77), .C1 (n_66_78), .C2 (n_72_75) );
AOI211_X1 g_55_81 (.ZN (n_55_81), .A (n_58_78), .B (n_63_78), .C1 (n_67_76), .C2 (n_70_76) );
AOI211_X1 g_57_80 (.ZN (n_57_80), .A (n_56_79), .B (n_61_79), .C1 (n_65_77), .C2 (n_68_77) );
AOI211_X1 g_59_79 (.ZN (n_59_79), .A (n_55_81), .B (n_60_77), .C1 (n_63_78), .C2 (n_66_78) );
AOI211_X1 g_61_78 (.ZN (n_61_78), .A (n_57_80), .B (n_58_78), .C1 (n_61_79), .C2 (n_67_76) );
AOI211_X1 g_63_79 (.ZN (n_63_79), .A (n_59_79), .B (n_56_79), .C1 (n_60_77), .C2 (n_65_77) );
AOI211_X1 g_61_80 (.ZN (n_61_80), .A (n_61_78), .B (n_55_81), .C1 (n_58_78), .C2 (n_63_78) );
AOI211_X1 g_62_78 (.ZN (n_62_78), .A (n_63_79), .B (n_57_80), .C1 (n_56_79), .C2 (n_61_79) );
AOI211_X1 g_60_79 (.ZN (n_60_79), .A (n_61_80), .B (n_59_79), .C1 (n_55_81), .C2 (n_60_77) );
AOI211_X1 g_58_80 (.ZN (n_58_80), .A (n_62_78), .B (n_61_78), .C1 (n_57_80), .C2 (n_58_78) );
AOI211_X1 g_56_81 (.ZN (n_56_81), .A (n_60_79), .B (n_63_79), .C1 (n_59_79), .C2 (n_56_79) );
AOI211_X1 g_57_79 (.ZN (n_57_79), .A (n_58_80), .B (n_61_80), .C1 (n_61_78), .C2 (n_55_81) );
AOI211_X1 g_55_80 (.ZN (n_55_80), .A (n_56_81), .B (n_62_78), .C1 (n_63_79), .C2 (n_57_80) );
AOI211_X1 g_53_81 (.ZN (n_53_81), .A (n_57_79), .B (n_60_79), .C1 (n_61_80), .C2 (n_59_79) );
AOI211_X1 g_51_82 (.ZN (n_51_82), .A (n_55_80), .B (n_58_80), .C1 (n_62_78), .C2 (n_61_78) );
AOI211_X1 g_49_83 (.ZN (n_49_83), .A (n_53_81), .B (n_56_81), .C1 (n_60_79), .C2 (n_63_79) );
AOI211_X1 g_47_84 (.ZN (n_47_84), .A (n_51_82), .B (n_57_79), .C1 (n_58_80), .C2 (n_61_80) );
AOI211_X1 g_45_85 (.ZN (n_45_85), .A (n_49_83), .B (n_55_80), .C1 (n_56_81), .C2 (n_62_78) );
AOI211_X1 g_44_83 (.ZN (n_44_83), .A (n_47_84), .B (n_53_81), .C1 (n_57_79), .C2 (n_60_79) );
AOI211_X1 g_42_84 (.ZN (n_42_84), .A (n_45_85), .B (n_51_82), .C1 (n_55_80), .C2 (n_58_80) );
AOI211_X1 g_41_86 (.ZN (n_41_86), .A (n_44_83), .B (n_49_83), .C1 (n_53_81), .C2 (n_56_81) );
AOI211_X1 g_43_85 (.ZN (n_43_85), .A (n_42_84), .B (n_47_84), .C1 (n_51_82), .C2 (n_57_79) );
AOI211_X1 g_45_84 (.ZN (n_45_84), .A (n_41_86), .B (n_45_85), .C1 (n_49_83), .C2 (n_55_80) );
AOI211_X1 g_47_85 (.ZN (n_47_85), .A (n_43_85), .B (n_44_83), .C1 (n_47_84), .C2 (n_53_81) );
AOI211_X1 g_45_86 (.ZN (n_45_86), .A (n_45_84), .B (n_42_84), .C1 (n_45_85), .C2 (n_51_82) );
AOI211_X1 g_46_84 (.ZN (n_46_84), .A (n_47_85), .B (n_41_86), .C1 (n_44_83), .C2 (n_49_83) );
AOI211_X1 g_44_85 (.ZN (n_44_85), .A (n_45_86), .B (n_43_85), .C1 (n_42_84), .C2 (n_47_84) );
AOI211_X1 g_42_86 (.ZN (n_42_86), .A (n_46_84), .B (n_45_84), .C1 (n_41_86), .C2 (n_45_85) );
AOI211_X1 g_40_87 (.ZN (n_40_87), .A (n_44_85), .B (n_47_85), .C1 (n_43_85), .C2 (n_44_83) );
AOI211_X1 g_38_86 (.ZN (n_38_86), .A (n_42_86), .B (n_45_86), .C1 (n_45_84), .C2 (n_42_84) );
AOI211_X1 g_36_87 (.ZN (n_36_87), .A (n_40_87), .B (n_46_84), .C1 (n_47_85), .C2 (n_41_86) );
AOI211_X1 g_34_88 (.ZN (n_34_88), .A (n_38_86), .B (n_44_85), .C1 (n_45_86), .C2 (n_43_85) );
AOI211_X1 g_32_89 (.ZN (n_32_89), .A (n_36_87), .B (n_42_86), .C1 (n_46_84), .C2 (n_45_84) );
AOI211_X1 g_30_90 (.ZN (n_30_90), .A (n_34_88), .B (n_40_87), .C1 (n_44_85), .C2 (n_47_85) );
AOI211_X1 g_28_91 (.ZN (n_28_91), .A (n_32_89), .B (n_38_86), .C1 (n_42_86), .C2 (n_45_86) );
AOI211_X1 g_27_93 (.ZN (n_27_93), .A (n_30_90), .B (n_36_87), .C1 (n_40_87), .C2 (n_46_84) );
AOI211_X1 g_25_92 (.ZN (n_25_92), .A (n_28_91), .B (n_34_88), .C1 (n_38_86), .C2 (n_44_85) );
AOI211_X1 g_27_91 (.ZN (n_27_91), .A (n_27_93), .B (n_32_89), .C1 (n_36_87), .C2 (n_42_86) );
AOI211_X1 g_29_90 (.ZN (n_29_90), .A (n_25_92), .B (n_30_90), .C1 (n_34_88), .C2 (n_40_87) );
AOI211_X1 g_31_89 (.ZN (n_31_89), .A (n_27_91), .B (n_28_91), .C1 (n_32_89), .C2 (n_38_86) );
AOI211_X1 g_33_88 (.ZN (n_33_88), .A (n_29_90), .B (n_27_93), .C1 (n_30_90), .C2 (n_36_87) );
AOI211_X1 g_32_90 (.ZN (n_32_90), .A (n_31_89), .B (n_25_92), .C1 (n_28_91), .C2 (n_34_88) );
AOI211_X1 g_34_89 (.ZN (n_34_89), .A (n_33_88), .B (n_27_91), .C1 (n_27_93), .C2 (n_32_89) );
AOI211_X1 g_36_88 (.ZN (n_36_88), .A (n_32_90), .B (n_29_90), .C1 (n_25_92), .C2 (n_30_90) );
AOI211_X1 g_38_87 (.ZN (n_38_87), .A (n_34_89), .B (n_31_89), .C1 (n_27_91), .C2 (n_28_91) );
AOI211_X1 g_40_86 (.ZN (n_40_86), .A (n_36_88), .B (n_33_88), .C1 (n_29_90), .C2 (n_27_93) );
AOI211_X1 g_42_85 (.ZN (n_42_85), .A (n_38_87), .B (n_32_90), .C1 (n_31_89), .C2 (n_25_92) );
AOI211_X1 g_44_84 (.ZN (n_44_84), .A (n_40_86), .B (n_34_89), .C1 (n_33_88), .C2 (n_27_91) );
AOI211_X1 g_43_86 (.ZN (n_43_86), .A (n_42_85), .B (n_36_88), .C1 (n_32_90), .C2 (n_29_90) );
AOI211_X1 g_41_87 (.ZN (n_41_87), .A (n_44_84), .B (n_38_87), .C1 (n_34_89), .C2 (n_31_89) );
AOI211_X1 g_39_88 (.ZN (n_39_88), .A (n_43_86), .B (n_40_86), .C1 (n_36_88), .C2 (n_33_88) );
AOI211_X1 g_37_89 (.ZN (n_37_89), .A (n_41_87), .B (n_42_85), .C1 (n_38_87), .C2 (n_32_90) );
AOI211_X1 g_35_90 (.ZN (n_35_90), .A (n_39_88), .B (n_44_84), .C1 (n_40_86), .C2 (n_34_89) );
AOI211_X1 g_33_91 (.ZN (n_33_91), .A (n_37_89), .B (n_43_86), .C1 (n_42_85), .C2 (n_36_88) );
AOI211_X1 g_31_92 (.ZN (n_31_92), .A (n_35_90), .B (n_41_87), .C1 (n_44_84), .C2 (n_38_87) );
AOI211_X1 g_29_93 (.ZN (n_29_93), .A (n_33_91), .B (n_39_88), .C1 (n_43_86), .C2 (n_40_86) );
AOI211_X1 g_30_91 (.ZN (n_30_91), .A (n_31_92), .B (n_37_89), .C1 (n_41_87), .C2 (n_42_85) );
AOI211_X1 g_28_92 (.ZN (n_28_92), .A (n_29_93), .B (n_35_90), .C1 (n_39_88), .C2 (n_44_84) );
AOI211_X1 g_26_93 (.ZN (n_26_93), .A (n_30_91), .B (n_33_91), .C1 (n_37_89), .C2 (n_43_86) );
AOI211_X1 g_24_94 (.ZN (n_24_94), .A (n_28_92), .B (n_31_92), .C1 (n_35_90), .C2 (n_41_87) );
AOI211_X1 g_22_95 (.ZN (n_22_95), .A (n_26_93), .B (n_29_93), .C1 (n_33_91), .C2 (n_39_88) );
AOI211_X1 g_23_93 (.ZN (n_23_93), .A (n_24_94), .B (n_30_91), .C1 (n_31_92), .C2 (n_37_89) );
AOI211_X1 g_21_94 (.ZN (n_21_94), .A (n_22_95), .B (n_28_92), .C1 (n_29_93), .C2 (n_35_90) );
AOI211_X1 g_19_95 (.ZN (n_19_95), .A (n_23_93), .B (n_26_93), .C1 (n_30_91), .C2 (n_33_91) );
AOI211_X1 g_17_96 (.ZN (n_17_96), .A (n_21_94), .B (n_24_94), .C1 (n_28_92), .C2 (n_31_92) );
AOI211_X1 g_16_98 (.ZN (n_16_98), .A (n_19_95), .B (n_22_95), .C1 (n_26_93), .C2 (n_29_93) );
AOI211_X1 g_18_97 (.ZN (n_18_97), .A (n_17_96), .B (n_23_93), .C1 (n_24_94), .C2 (n_30_91) );
AOI211_X1 g_20_96 (.ZN (n_20_96), .A (n_16_98), .B (n_21_94), .C1 (n_22_95), .C2 (n_28_92) );
AOI211_X1 g_19_98 (.ZN (n_19_98), .A (n_18_97), .B (n_19_95), .C1 (n_23_93), .C2 (n_26_93) );
AOI211_X1 g_17_97 (.ZN (n_17_97), .A (n_20_96), .B (n_17_96), .C1 (n_21_94), .C2 (n_24_94) );
AOI211_X1 g_19_96 (.ZN (n_19_96), .A (n_19_98), .B (n_16_98), .C1 (n_19_95), .C2 (n_22_95) );
AOI211_X1 g_21_95 (.ZN (n_21_95), .A (n_17_97), .B (n_18_97), .C1 (n_17_96), .C2 (n_23_93) );
AOI211_X1 g_20_97 (.ZN (n_20_97), .A (n_19_96), .B (n_20_96), .C1 (n_16_98), .C2 (n_21_94) );
AOI211_X1 g_22_96 (.ZN (n_22_96), .A (n_21_95), .B (n_19_98), .C1 (n_18_97), .C2 (n_19_95) );
AOI211_X1 g_24_95 (.ZN (n_24_95), .A (n_20_97), .B (n_17_97), .C1 (n_20_96), .C2 (n_17_96) );
AOI211_X1 g_26_94 (.ZN (n_26_94), .A (n_22_96), .B (n_19_96), .C1 (n_19_98), .C2 (n_16_98) );
AOI211_X1 g_28_93 (.ZN (n_28_93), .A (n_24_95), .B (n_21_95), .C1 (n_17_97), .C2 (n_18_97) );
AOI211_X1 g_30_92 (.ZN (n_30_92), .A (n_26_94), .B (n_20_97), .C1 (n_19_96), .C2 (n_20_96) );
AOI211_X1 g_32_91 (.ZN (n_32_91), .A (n_28_93), .B (n_22_96), .C1 (n_21_95), .C2 (n_19_98) );
AOI211_X1 g_34_90 (.ZN (n_34_90), .A (n_30_92), .B (n_24_95), .C1 (n_20_97), .C2 (n_17_97) );
AOI211_X1 g_36_89 (.ZN (n_36_89), .A (n_32_91), .B (n_26_94), .C1 (n_22_96), .C2 (n_19_96) );
AOI211_X1 g_38_88 (.ZN (n_38_88), .A (n_34_90), .B (n_28_93), .C1 (n_24_95), .C2 (n_21_95) );
AOI211_X1 g_37_90 (.ZN (n_37_90), .A (n_36_89), .B (n_30_92), .C1 (n_26_94), .C2 (n_20_97) );
AOI211_X1 g_35_89 (.ZN (n_35_89), .A (n_38_88), .B (n_32_91), .C1 (n_28_93), .C2 (n_22_96) );
AOI211_X1 g_37_88 (.ZN (n_37_88), .A (n_37_90), .B (n_34_90), .C1 (n_30_92), .C2 (n_24_95) );
AOI211_X1 g_39_87 (.ZN (n_39_87), .A (n_35_89), .B (n_36_89), .C1 (n_32_91), .C2 (n_26_94) );
AOI211_X1 g_38_89 (.ZN (n_38_89), .A (n_37_88), .B (n_38_88), .C1 (n_34_90), .C2 (n_28_93) );
AOI211_X1 g_40_88 (.ZN (n_40_88), .A (n_39_87), .B (n_37_90), .C1 (n_36_89), .C2 (n_30_92) );
AOI211_X1 g_42_87 (.ZN (n_42_87), .A (n_38_89), .B (n_35_89), .C1 (n_38_88), .C2 (n_32_91) );
AOI211_X1 g_44_86 (.ZN (n_44_86), .A (n_40_88), .B (n_37_88), .C1 (n_37_90), .C2 (n_34_90) );
AOI211_X1 g_46_85 (.ZN (n_46_85), .A (n_42_87), .B (n_39_87), .C1 (n_35_89), .C2 (n_36_89) );
AOI211_X1 g_48_84 (.ZN (n_48_84), .A (n_44_86), .B (n_38_89), .C1 (n_37_88), .C2 (n_38_88) );
AOI211_X1 g_50_83 (.ZN (n_50_83), .A (n_46_85), .B (n_40_88), .C1 (n_39_87), .C2 (n_37_90) );
AOI211_X1 g_52_82 (.ZN (n_52_82), .A (n_48_84), .B (n_42_87), .C1 (n_38_89), .C2 (n_35_89) );
AOI211_X1 g_54_81 (.ZN (n_54_81), .A (n_50_83), .B (n_44_86), .C1 (n_40_88), .C2 (n_37_88) );
AOI211_X1 g_56_80 (.ZN (n_56_80), .A (n_52_82), .B (n_46_85), .C1 (n_42_87), .C2 (n_39_87) );
AOI211_X1 g_58_79 (.ZN (n_58_79), .A (n_54_81), .B (n_48_84), .C1 (n_44_86), .C2 (n_38_89) );
AOI211_X1 g_59_81 (.ZN (n_59_81), .A (n_56_80), .B (n_50_83), .C1 (n_46_85), .C2 (n_40_88) );
AOI211_X1 g_57_82 (.ZN (n_57_82), .A (n_58_79), .B (n_52_82), .C1 (n_48_84), .C2 (n_42_87) );
AOI211_X1 g_55_83 (.ZN (n_55_83), .A (n_59_81), .B (n_54_81), .C1 (n_50_83), .C2 (n_44_86) );
AOI211_X1 g_53_82 (.ZN (n_53_82), .A (n_57_82), .B (n_56_80), .C1 (n_52_82), .C2 (n_46_85) );
AOI211_X1 g_51_83 (.ZN (n_51_83), .A (n_55_83), .B (n_58_79), .C1 (n_54_81), .C2 (n_48_84) );
AOI211_X1 g_50_85 (.ZN (n_50_85), .A (n_53_82), .B (n_59_81), .C1 (n_56_80), .C2 (n_50_83) );
AOI211_X1 g_52_84 (.ZN (n_52_84), .A (n_51_83), .B (n_57_82), .C1 (n_58_79), .C2 (n_52_82) );
AOI211_X1 g_54_83 (.ZN (n_54_83), .A (n_50_85), .B (n_55_83), .C1 (n_59_81), .C2 (n_54_81) );
AOI211_X1 g_56_82 (.ZN (n_56_82), .A (n_52_84), .B (n_53_82), .C1 (n_57_82), .C2 (n_56_80) );
AOI211_X1 g_58_81 (.ZN (n_58_81), .A (n_54_83), .B (n_51_83), .C1 (n_55_83), .C2 (n_58_79) );
AOI211_X1 g_60_80 (.ZN (n_60_80), .A (n_56_82), .B (n_50_85), .C1 (n_53_82), .C2 (n_59_81) );
AOI211_X1 g_62_79 (.ZN (n_62_79), .A (n_58_81), .B (n_52_84), .C1 (n_51_83), .C2 (n_57_82) );
AOI211_X1 g_64_78 (.ZN (n_64_78), .A (n_60_80), .B (n_54_83), .C1 (n_50_85), .C2 (n_55_83) );
AOI211_X1 g_66_77 (.ZN (n_66_77), .A (n_62_79), .B (n_56_82), .C1 (n_52_84), .C2 (n_53_82) );
AOI211_X1 g_68_76 (.ZN (n_68_76), .A (n_64_78), .B (n_58_81), .C1 (n_54_83), .C2 (n_51_83) );
AOI211_X1 g_70_75 (.ZN (n_70_75), .A (n_66_77), .B (n_60_80), .C1 (n_56_82), .C2 (n_50_85) );
AOI211_X1 g_72_74 (.ZN (n_72_74), .A (n_68_76), .B (n_62_79), .C1 (n_58_81), .C2 (n_52_84) );
AOI211_X1 g_74_73 (.ZN (n_74_73), .A (n_70_75), .B (n_64_78), .C1 (n_60_80), .C2 (n_54_83) );
AOI211_X1 g_76_72 (.ZN (n_76_72), .A (n_72_74), .B (n_66_77), .C1 (n_62_79), .C2 (n_56_82) );
AOI211_X1 g_78_71 (.ZN (n_78_71), .A (n_74_73), .B (n_68_76), .C1 (n_64_78), .C2 (n_58_81) );
AOI211_X1 g_80_70 (.ZN (n_80_70), .A (n_76_72), .B (n_70_75), .C1 (n_66_77), .C2 (n_60_80) );
AOI211_X1 g_82_69 (.ZN (n_82_69), .A (n_78_71), .B (n_72_74), .C1 (n_68_76), .C2 (n_62_79) );
AOI211_X1 g_84_68 (.ZN (n_84_68), .A (n_80_70), .B (n_74_73), .C1 (n_70_75), .C2 (n_64_78) );
AOI211_X1 g_86_67 (.ZN (n_86_67), .A (n_82_69), .B (n_76_72), .C1 (n_72_74), .C2 (n_66_77) );
AOI211_X1 g_88_66 (.ZN (n_88_66), .A (n_84_68), .B (n_78_71), .C1 (n_74_73), .C2 (n_68_76) );
AOI211_X1 g_90_65 (.ZN (n_90_65), .A (n_86_67), .B (n_80_70), .C1 (n_76_72), .C2 (n_70_75) );
AOI211_X1 g_92_64 (.ZN (n_92_64), .A (n_88_66), .B (n_82_69), .C1 (n_78_71), .C2 (n_72_74) );
AOI211_X1 g_94_63 (.ZN (n_94_63), .A (n_90_65), .B (n_84_68), .C1 (n_80_70), .C2 (n_74_73) );
AOI211_X1 g_96_62 (.ZN (n_96_62), .A (n_92_64), .B (n_86_67), .C1 (n_82_69), .C2 (n_76_72) );
AOI211_X1 g_98_61 (.ZN (n_98_61), .A (n_94_63), .B (n_88_66), .C1 (n_84_68), .C2 (n_78_71) );
AOI211_X1 g_100_60 (.ZN (n_100_60), .A (n_96_62), .B (n_90_65), .C1 (n_86_67), .C2 (n_80_70) );
AOI211_X1 g_99_62 (.ZN (n_99_62), .A (n_98_61), .B (n_92_64), .C1 (n_88_66), .C2 (n_82_69) );
AOI211_X1 g_101_61 (.ZN (n_101_61), .A (n_100_60), .B (n_94_63), .C1 (n_90_65), .C2 (n_84_68) );
AOI211_X1 g_103_60 (.ZN (n_103_60), .A (n_99_62), .B (n_96_62), .C1 (n_92_64), .C2 (n_86_67) );
AOI211_X1 g_105_59 (.ZN (n_105_59), .A (n_101_61), .B (n_98_61), .C1 (n_94_63), .C2 (n_88_66) );
AOI211_X1 g_107_58 (.ZN (n_107_58), .A (n_103_60), .B (n_100_60), .C1 (n_96_62), .C2 (n_90_65) );
AOI211_X1 g_109_57 (.ZN (n_109_57), .A (n_105_59), .B (n_99_62), .C1 (n_98_61), .C2 (n_92_64) );
AOI211_X1 g_108_59 (.ZN (n_108_59), .A (n_107_58), .B (n_101_61), .C1 (n_100_60), .C2 (n_94_63) );
AOI211_X1 g_106_58 (.ZN (n_106_58), .A (n_109_57), .B (n_103_60), .C1 (n_99_62), .C2 (n_96_62) );
AOI211_X1 g_108_57 (.ZN (n_108_57), .A (n_108_59), .B (n_105_59), .C1 (n_101_61), .C2 (n_98_61) );
AOI211_X1 g_110_56 (.ZN (n_110_56), .A (n_106_58), .B (n_107_58), .C1 (n_103_60), .C2 (n_100_60) );
AOI211_X1 g_112_55 (.ZN (n_112_55), .A (n_108_57), .B (n_109_57), .C1 (n_105_59), .C2 (n_99_62) );
AOI211_X1 g_114_54 (.ZN (n_114_54), .A (n_110_56), .B (n_108_59), .C1 (n_107_58), .C2 (n_101_61) );
AOI211_X1 g_116_53 (.ZN (n_116_53), .A (n_112_55), .B (n_106_58), .C1 (n_109_57), .C2 (n_103_60) );
AOI211_X1 g_118_52 (.ZN (n_118_52), .A (n_114_54), .B (n_108_57), .C1 (n_108_59), .C2 (n_105_59) );
AOI211_X1 g_120_51 (.ZN (n_120_51), .A (n_116_53), .B (n_110_56), .C1 (n_106_58), .C2 (n_107_58) );
AOI211_X1 g_122_50 (.ZN (n_122_50), .A (n_118_52), .B (n_112_55), .C1 (n_108_57), .C2 (n_109_57) );
AOI211_X1 g_124_49 (.ZN (n_124_49), .A (n_120_51), .B (n_114_54), .C1 (n_110_56), .C2 (n_108_59) );
AOI211_X1 g_126_48 (.ZN (n_126_48), .A (n_122_50), .B (n_116_53), .C1 (n_112_55), .C2 (n_106_58) );
AOI211_X1 g_128_47 (.ZN (n_128_47), .A (n_124_49), .B (n_118_52), .C1 (n_114_54), .C2 (n_108_57) );
AOI211_X1 g_130_46 (.ZN (n_130_46), .A (n_126_48), .B (n_120_51), .C1 (n_116_53), .C2 (n_110_56) );
AOI211_X1 g_132_45 (.ZN (n_132_45), .A (n_128_47), .B (n_122_50), .C1 (n_118_52), .C2 (n_112_55) );
AOI211_X1 g_134_44 (.ZN (n_134_44), .A (n_130_46), .B (n_124_49), .C1 (n_120_51), .C2 (n_114_54) );
AOI211_X1 g_136_43 (.ZN (n_136_43), .A (n_132_45), .B (n_126_48), .C1 (n_122_50), .C2 (n_116_53) );
AOI211_X1 g_138_42 (.ZN (n_138_42), .A (n_134_44), .B (n_128_47), .C1 (n_124_49), .C2 (n_118_52) );
AOI211_X1 g_140_41 (.ZN (n_140_41), .A (n_136_43), .B (n_130_46), .C1 (n_126_48), .C2 (n_120_51) );
AOI211_X1 g_142_40 (.ZN (n_142_40), .A (n_138_42), .B (n_132_45), .C1 (n_128_47), .C2 (n_122_50) );
AOI211_X1 g_144_39 (.ZN (n_144_39), .A (n_140_41), .B (n_134_44), .C1 (n_130_46), .C2 (n_124_49) );
AOI211_X1 g_146_40 (.ZN (n_146_40), .A (n_142_40), .B (n_136_43), .C1 (n_132_45), .C2 (n_126_48) );
AOI211_X1 g_147_42 (.ZN (n_147_42), .A (n_144_39), .B (n_138_42), .C1 (n_134_44), .C2 (n_128_47) );
AOI211_X1 g_145_41 (.ZN (n_145_41), .A (n_146_40), .B (n_140_41), .C1 (n_136_43), .C2 (n_130_46) );
AOI211_X1 g_143_40 (.ZN (n_143_40), .A (n_147_42), .B (n_142_40), .C1 (n_138_42), .C2 (n_132_45) );
AOI211_X1 g_141_41 (.ZN (n_141_41), .A (n_145_41), .B (n_144_39), .C1 (n_140_41), .C2 (n_134_44) );
AOI211_X1 g_139_42 (.ZN (n_139_42), .A (n_143_40), .B (n_146_40), .C1 (n_142_40), .C2 (n_136_43) );
AOI211_X1 g_137_43 (.ZN (n_137_43), .A (n_141_41), .B (n_147_42), .C1 (n_144_39), .C2 (n_138_42) );
AOI211_X1 g_135_44 (.ZN (n_135_44), .A (n_139_42), .B (n_145_41), .C1 (n_146_40), .C2 (n_140_41) );
AOI211_X1 g_133_45 (.ZN (n_133_45), .A (n_137_43), .B (n_143_40), .C1 (n_147_42), .C2 (n_142_40) );
AOI211_X1 g_131_46 (.ZN (n_131_46), .A (n_135_44), .B (n_141_41), .C1 (n_145_41), .C2 (n_144_39) );
AOI211_X1 g_129_47 (.ZN (n_129_47), .A (n_133_45), .B (n_139_42), .C1 (n_143_40), .C2 (n_146_40) );
AOI211_X1 g_127_48 (.ZN (n_127_48), .A (n_131_46), .B (n_137_43), .C1 (n_141_41), .C2 (n_147_42) );
AOI211_X1 g_125_49 (.ZN (n_125_49), .A (n_129_47), .B (n_135_44), .C1 (n_139_42), .C2 (n_145_41) );
AOI211_X1 g_123_50 (.ZN (n_123_50), .A (n_127_48), .B (n_133_45), .C1 (n_137_43), .C2 (n_143_40) );
AOI211_X1 g_121_51 (.ZN (n_121_51), .A (n_125_49), .B (n_131_46), .C1 (n_135_44), .C2 (n_141_41) );
AOI211_X1 g_119_52 (.ZN (n_119_52), .A (n_123_50), .B (n_129_47), .C1 (n_133_45), .C2 (n_139_42) );
AOI211_X1 g_117_53 (.ZN (n_117_53), .A (n_121_51), .B (n_127_48), .C1 (n_131_46), .C2 (n_137_43) );
AOI211_X1 g_115_54 (.ZN (n_115_54), .A (n_119_52), .B (n_125_49), .C1 (n_129_47), .C2 (n_135_44) );
AOI211_X1 g_113_55 (.ZN (n_113_55), .A (n_117_53), .B (n_123_50), .C1 (n_127_48), .C2 (n_133_45) );
AOI211_X1 g_112_57 (.ZN (n_112_57), .A (n_115_54), .B (n_121_51), .C1 (n_125_49), .C2 (n_131_46) );
AOI211_X1 g_110_58 (.ZN (n_110_58), .A (n_113_55), .B (n_119_52), .C1 (n_123_50), .C2 (n_129_47) );
AOI211_X1 g_109_60 (.ZN (n_109_60), .A (n_112_57), .B (n_117_53), .C1 (n_121_51), .C2 (n_127_48) );
AOI211_X1 g_108_58 (.ZN (n_108_58), .A (n_110_58), .B (n_115_54), .C1 (n_119_52), .C2 (n_125_49) );
AOI211_X1 g_110_57 (.ZN (n_110_57), .A (n_109_60), .B (n_113_55), .C1 (n_117_53), .C2 (n_123_50) );
AOI211_X1 g_112_56 (.ZN (n_112_56), .A (n_108_58), .B (n_112_57), .C1 (n_115_54), .C2 (n_121_51) );
AOI211_X1 g_114_55 (.ZN (n_114_55), .A (n_110_57), .B (n_110_58), .C1 (n_113_55), .C2 (n_119_52) );
AOI211_X1 g_116_54 (.ZN (n_116_54), .A (n_112_56), .B (n_109_60), .C1 (n_112_57), .C2 (n_117_53) );
AOI211_X1 g_118_53 (.ZN (n_118_53), .A (n_114_55), .B (n_108_58), .C1 (n_110_58), .C2 (n_115_54) );
AOI211_X1 g_120_52 (.ZN (n_120_52), .A (n_116_54), .B (n_110_57), .C1 (n_109_60), .C2 (n_113_55) );
AOI211_X1 g_122_51 (.ZN (n_122_51), .A (n_118_53), .B (n_112_56), .C1 (n_108_58), .C2 (n_112_57) );
AOI211_X1 g_124_50 (.ZN (n_124_50), .A (n_120_52), .B (n_114_55), .C1 (n_110_57), .C2 (n_110_58) );
AOI211_X1 g_126_49 (.ZN (n_126_49), .A (n_122_51), .B (n_116_54), .C1 (n_112_56), .C2 (n_109_60) );
AOI211_X1 g_128_48 (.ZN (n_128_48), .A (n_124_50), .B (n_118_53), .C1 (n_114_55), .C2 (n_108_58) );
AOI211_X1 g_130_47 (.ZN (n_130_47), .A (n_126_49), .B (n_120_52), .C1 (n_116_54), .C2 (n_110_57) );
AOI211_X1 g_132_46 (.ZN (n_132_46), .A (n_128_48), .B (n_122_51), .C1 (n_118_53), .C2 (n_112_56) );
AOI211_X1 g_134_45 (.ZN (n_134_45), .A (n_130_47), .B (n_124_50), .C1 (n_120_52), .C2 (n_114_55) );
AOI211_X1 g_136_44 (.ZN (n_136_44), .A (n_132_46), .B (n_126_49), .C1 (n_122_51), .C2 (n_116_54) );
AOI211_X1 g_138_43 (.ZN (n_138_43), .A (n_134_45), .B (n_128_48), .C1 (n_124_50), .C2 (n_118_53) );
AOI211_X1 g_140_42 (.ZN (n_140_42), .A (n_136_44), .B (n_130_47), .C1 (n_126_49), .C2 (n_120_52) );
AOI211_X1 g_139_44 (.ZN (n_139_44), .A (n_138_43), .B (n_132_46), .C1 (n_128_48), .C2 (n_122_51) );
AOI211_X1 g_141_43 (.ZN (n_141_43), .A (n_140_42), .B (n_134_45), .C1 (n_130_47), .C2 (n_124_50) );
AOI211_X1 g_143_42 (.ZN (n_143_42), .A (n_139_44), .B (n_136_44), .C1 (n_132_46), .C2 (n_126_49) );
AOI211_X1 g_145_43 (.ZN (n_145_43), .A (n_141_43), .B (n_138_43), .C1 (n_134_45), .C2 (n_128_48) );
AOI211_X1 g_144_41 (.ZN (n_144_41), .A (n_143_42), .B (n_140_42), .C1 (n_136_44), .C2 (n_130_47) );
AOI211_X1 g_142_42 (.ZN (n_142_42), .A (n_145_43), .B (n_139_44), .C1 (n_138_43), .C2 (n_132_46) );
AOI211_X1 g_140_43 (.ZN (n_140_43), .A (n_144_41), .B (n_141_43), .C1 (n_140_42), .C2 (n_134_45) );
AOI211_X1 g_138_44 (.ZN (n_138_44), .A (n_142_42), .B (n_143_42), .C1 (n_139_44), .C2 (n_136_44) );
AOI211_X1 g_136_45 (.ZN (n_136_45), .A (n_140_43), .B (n_145_43), .C1 (n_141_43), .C2 (n_138_43) );
AOI211_X1 g_134_46 (.ZN (n_134_46), .A (n_138_44), .B (n_144_41), .C1 (n_143_42), .C2 (n_140_42) );
AOI211_X1 g_132_47 (.ZN (n_132_47), .A (n_136_45), .B (n_142_42), .C1 (n_145_43), .C2 (n_139_44) );
AOI211_X1 g_130_48 (.ZN (n_130_48), .A (n_134_46), .B (n_140_43), .C1 (n_144_41), .C2 (n_141_43) );
AOI211_X1 g_128_49 (.ZN (n_128_49), .A (n_132_47), .B (n_138_44), .C1 (n_142_42), .C2 (n_143_42) );
AOI211_X1 g_126_50 (.ZN (n_126_50), .A (n_130_48), .B (n_136_45), .C1 (n_140_43), .C2 (n_145_43) );
AOI211_X1 g_124_51 (.ZN (n_124_51), .A (n_128_49), .B (n_134_46), .C1 (n_138_44), .C2 (n_144_41) );
AOI211_X1 g_122_52 (.ZN (n_122_52), .A (n_126_50), .B (n_132_47), .C1 (n_136_45), .C2 (n_142_42) );
AOI211_X1 g_120_53 (.ZN (n_120_53), .A (n_124_51), .B (n_130_48), .C1 (n_134_46), .C2 (n_140_43) );
AOI211_X1 g_118_54 (.ZN (n_118_54), .A (n_122_52), .B (n_128_49), .C1 (n_132_47), .C2 (n_138_44) );
AOI211_X1 g_116_55 (.ZN (n_116_55), .A (n_120_53), .B (n_126_50), .C1 (n_130_48), .C2 (n_136_45) );
AOI211_X1 g_114_56 (.ZN (n_114_56), .A (n_118_54), .B (n_124_51), .C1 (n_128_49), .C2 (n_134_46) );
AOI211_X1 g_113_58 (.ZN (n_113_58), .A (n_116_55), .B (n_122_52), .C1 (n_126_50), .C2 (n_132_47) );
AOI211_X1 g_111_57 (.ZN (n_111_57), .A (n_114_56), .B (n_120_53), .C1 (n_124_51), .C2 (n_130_48) );
AOI211_X1 g_113_56 (.ZN (n_113_56), .A (n_113_58), .B (n_118_54), .C1 (n_122_52), .C2 (n_128_49) );
AOI211_X1 g_115_55 (.ZN (n_115_55), .A (n_111_57), .B (n_116_55), .C1 (n_120_53), .C2 (n_126_50) );
AOI211_X1 g_117_54 (.ZN (n_117_54), .A (n_113_56), .B (n_114_56), .C1 (n_118_54), .C2 (n_124_51) );
AOI211_X1 g_119_53 (.ZN (n_119_53), .A (n_115_55), .B (n_113_58), .C1 (n_116_55), .C2 (n_122_52) );
AOI211_X1 g_121_52 (.ZN (n_121_52), .A (n_117_54), .B (n_111_57), .C1 (n_114_56), .C2 (n_120_53) );
AOI211_X1 g_123_51 (.ZN (n_123_51), .A (n_119_53), .B (n_113_56), .C1 (n_113_58), .C2 (n_118_54) );
AOI211_X1 g_125_50 (.ZN (n_125_50), .A (n_121_52), .B (n_115_55), .C1 (n_111_57), .C2 (n_116_55) );
AOI211_X1 g_127_49 (.ZN (n_127_49), .A (n_123_51), .B (n_117_54), .C1 (n_113_56), .C2 (n_114_56) );
AOI211_X1 g_129_48 (.ZN (n_129_48), .A (n_125_50), .B (n_119_53), .C1 (n_115_55), .C2 (n_113_58) );
AOI211_X1 g_131_47 (.ZN (n_131_47), .A (n_127_49), .B (n_121_52), .C1 (n_117_54), .C2 (n_111_57) );
AOI211_X1 g_133_46 (.ZN (n_133_46), .A (n_129_48), .B (n_123_51), .C1 (n_119_53), .C2 (n_113_56) );
AOI211_X1 g_135_45 (.ZN (n_135_45), .A (n_131_47), .B (n_125_50), .C1 (n_121_52), .C2 (n_115_55) );
AOI211_X1 g_137_44 (.ZN (n_137_44), .A (n_133_46), .B (n_127_49), .C1 (n_123_51), .C2 (n_117_54) );
AOI211_X1 g_139_43 (.ZN (n_139_43), .A (n_135_45), .B (n_129_48), .C1 (n_125_50), .C2 (n_119_53) );
AOI211_X1 g_141_42 (.ZN (n_141_42), .A (n_137_44), .B (n_131_47), .C1 (n_127_49), .C2 (n_121_52) );
AOI211_X1 g_143_41 (.ZN (n_143_41), .A (n_139_43), .B (n_133_46), .C1 (n_129_48), .C2 (n_123_51) );
AOI211_X1 g_145_40 (.ZN (n_145_40), .A (n_141_42), .B (n_135_45), .C1 (n_131_47), .C2 (n_125_50) );
AOI211_X1 g_147_41 (.ZN (n_147_41), .A (n_143_41), .B (n_137_44), .C1 (n_133_46), .C2 (n_127_49) );
AOI211_X1 g_145_42 (.ZN (n_145_42), .A (n_145_40), .B (n_139_43), .C1 (n_135_45), .C2 (n_129_48) );
AOI211_X1 g_143_43 (.ZN (n_143_43), .A (n_147_41), .B (n_141_42), .C1 (n_137_44), .C2 (n_131_47) );
AOI211_X1 g_141_44 (.ZN (n_141_44), .A (n_145_42), .B (n_143_41), .C1 (n_139_43), .C2 (n_133_46) );
AOI211_X1 g_139_45 (.ZN (n_139_45), .A (n_143_43), .B (n_145_40), .C1 (n_141_42), .C2 (n_135_45) );
AOI211_X1 g_137_46 (.ZN (n_137_46), .A (n_141_44), .B (n_147_41), .C1 (n_143_41), .C2 (n_137_44) );
AOI211_X1 g_135_47 (.ZN (n_135_47), .A (n_139_45), .B (n_145_42), .C1 (n_145_40), .C2 (n_139_43) );
AOI211_X1 g_133_48 (.ZN (n_133_48), .A (n_137_46), .B (n_143_43), .C1 (n_147_41), .C2 (n_141_42) );
AOI211_X1 g_131_49 (.ZN (n_131_49), .A (n_135_47), .B (n_141_44), .C1 (n_145_42), .C2 (n_143_41) );
AOI211_X1 g_129_50 (.ZN (n_129_50), .A (n_133_48), .B (n_139_45), .C1 (n_143_43), .C2 (n_145_40) );
AOI211_X1 g_127_51 (.ZN (n_127_51), .A (n_131_49), .B (n_137_46), .C1 (n_141_44), .C2 (n_147_41) );
AOI211_X1 g_125_52 (.ZN (n_125_52), .A (n_129_50), .B (n_135_47), .C1 (n_139_45), .C2 (n_145_42) );
AOI211_X1 g_123_53 (.ZN (n_123_53), .A (n_127_51), .B (n_133_48), .C1 (n_137_46), .C2 (n_143_43) );
AOI211_X1 g_121_54 (.ZN (n_121_54), .A (n_125_52), .B (n_131_49), .C1 (n_135_47), .C2 (n_141_44) );
AOI211_X1 g_119_55 (.ZN (n_119_55), .A (n_123_53), .B (n_129_50), .C1 (n_133_48), .C2 (n_139_45) );
AOI211_X1 g_117_56 (.ZN (n_117_56), .A (n_121_54), .B (n_127_51), .C1 (n_131_49), .C2 (n_137_46) );
AOI211_X1 g_115_57 (.ZN (n_115_57), .A (n_119_55), .B (n_125_52), .C1 (n_129_50), .C2 (n_135_47) );
AOI211_X1 g_114_59 (.ZN (n_114_59), .A (n_117_56), .B (n_123_53), .C1 (n_127_51), .C2 (n_133_48) );
AOI211_X1 g_113_57 (.ZN (n_113_57), .A (n_115_57), .B (n_121_54), .C1 (n_125_52), .C2 (n_131_49) );
AOI211_X1 g_115_56 (.ZN (n_115_56), .A (n_114_59), .B (n_119_55), .C1 (n_123_53), .C2 (n_129_50) );
AOI211_X1 g_117_55 (.ZN (n_117_55), .A (n_113_57), .B (n_117_56), .C1 (n_121_54), .C2 (n_127_51) );
AOI211_X1 g_119_54 (.ZN (n_119_54), .A (n_115_56), .B (n_115_57), .C1 (n_119_55), .C2 (n_125_52) );
AOI211_X1 g_121_53 (.ZN (n_121_53), .A (n_117_55), .B (n_114_59), .C1 (n_117_56), .C2 (n_123_53) );
AOI211_X1 g_123_52 (.ZN (n_123_52), .A (n_119_54), .B (n_113_57), .C1 (n_115_57), .C2 (n_121_54) );
AOI211_X1 g_125_51 (.ZN (n_125_51), .A (n_121_53), .B (n_115_56), .C1 (n_114_59), .C2 (n_119_55) );
AOI211_X1 g_127_50 (.ZN (n_127_50), .A (n_123_52), .B (n_117_55), .C1 (n_113_57), .C2 (n_117_56) );
AOI211_X1 g_129_49 (.ZN (n_129_49), .A (n_125_51), .B (n_119_54), .C1 (n_115_56), .C2 (n_115_57) );
AOI211_X1 g_131_48 (.ZN (n_131_48), .A (n_127_50), .B (n_121_53), .C1 (n_117_55), .C2 (n_114_59) );
AOI211_X1 g_133_47 (.ZN (n_133_47), .A (n_129_49), .B (n_123_52), .C1 (n_119_54), .C2 (n_113_57) );
AOI211_X1 g_135_46 (.ZN (n_135_46), .A (n_131_48), .B (n_125_51), .C1 (n_121_53), .C2 (n_115_56) );
AOI211_X1 g_137_45 (.ZN (n_137_45), .A (n_133_47), .B (n_127_50), .C1 (n_123_52), .C2 (n_117_55) );
AOI211_X1 g_136_47 (.ZN (n_136_47), .A (n_135_46), .B (n_129_49), .C1 (n_125_51), .C2 (n_119_54) );
AOI211_X1 g_138_46 (.ZN (n_138_46), .A (n_137_45), .B (n_131_48), .C1 (n_127_50), .C2 (n_121_53) );
AOI211_X1 g_140_45 (.ZN (n_140_45), .A (n_136_47), .B (n_133_47), .C1 (n_129_49), .C2 (n_123_52) );
AOI211_X1 g_142_44 (.ZN (n_142_44), .A (n_138_46), .B (n_135_46), .C1 (n_131_48), .C2 (n_125_51) );
AOI211_X1 g_144_43 (.ZN (n_144_43), .A (n_140_45), .B (n_137_45), .C1 (n_133_47), .C2 (n_127_50) );
AOI211_X1 g_146_42 (.ZN (n_146_42), .A (n_142_44), .B (n_136_47), .C1 (n_135_46), .C2 (n_129_49) );
AOI211_X1 g_147_44 (.ZN (n_147_44), .A (n_144_43), .B (n_138_46), .C1 (n_137_45), .C2 (n_131_48) );
AOI211_X1 g_149_45 (.ZN (n_149_45), .A (n_146_42), .B (n_140_45), .C1 (n_136_47), .C2 (n_133_47) );
AOI211_X1 g_148_43 (.ZN (n_148_43), .A (n_147_44), .B (n_142_44), .C1 (n_138_46), .C2 (n_135_46) );
AOI211_X1 g_146_44 (.ZN (n_146_44), .A (n_149_45), .B (n_144_43), .C1 (n_140_45), .C2 (n_137_45) );
AOI211_X1 g_147_46 (.ZN (n_147_46), .A (n_148_43), .B (n_146_42), .C1 (n_142_44), .C2 (n_136_47) );
AOI211_X1 g_145_45 (.ZN (n_145_45), .A (n_146_44), .B (n_147_44), .C1 (n_144_43), .C2 (n_138_46) );
AOI211_X1 g_146_43 (.ZN (n_146_43), .A (n_147_46), .B (n_149_45), .C1 (n_146_42), .C2 (n_140_45) );
AOI211_X1 g_144_42 (.ZN (n_144_42), .A (n_145_45), .B (n_148_43), .C1 (n_147_44), .C2 (n_142_44) );
AOI211_X1 g_143_44 (.ZN (n_143_44), .A (n_146_43), .B (n_146_44), .C1 (n_149_45), .C2 (n_144_43) );
AOI211_X1 g_141_45 (.ZN (n_141_45), .A (n_144_42), .B (n_147_46), .C1 (n_148_43), .C2 (n_146_42) );
AOI211_X1 g_142_43 (.ZN (n_142_43), .A (n_143_44), .B (n_145_45), .C1 (n_146_44), .C2 (n_147_44) );
AOI211_X1 g_144_44 (.ZN (n_144_44), .A (n_141_45), .B (n_146_43), .C1 (n_147_46), .C2 (n_149_45) );
AOI211_X1 g_143_46 (.ZN (n_143_46), .A (n_142_43), .B (n_144_42), .C1 (n_145_45), .C2 (n_148_43) );
AOI211_X1 g_145_47 (.ZN (n_145_47), .A (n_144_44), .B (n_143_44), .C1 (n_146_43), .C2 (n_146_44) );
AOI211_X1 g_144_45 (.ZN (n_144_45), .A (n_143_46), .B (n_141_45), .C1 (n_144_42), .C2 (n_147_46) );
AOI211_X1 g_142_46 (.ZN (n_142_46), .A (n_145_47), .B (n_142_43), .C1 (n_143_44), .C2 (n_145_45) );
AOI211_X1 g_140_47 (.ZN (n_140_47), .A (n_144_45), .B (n_144_44), .C1 (n_141_45), .C2 (n_146_43) );
AOI211_X1 g_138_48 (.ZN (n_138_48), .A (n_142_46), .B (n_143_46), .C1 (n_142_43), .C2 (n_144_42) );
AOI211_X1 g_139_46 (.ZN (n_139_46), .A (n_140_47), .B (n_145_47), .C1 (n_144_44), .C2 (n_143_44) );
AOI211_X1 g_140_44 (.ZN (n_140_44), .A (n_138_48), .B (n_144_45), .C1 (n_143_46), .C2 (n_141_45) );
AOI211_X1 g_138_45 (.ZN (n_138_45), .A (n_139_46), .B (n_142_46), .C1 (n_145_47), .C2 (n_142_43) );
AOI211_X1 g_136_46 (.ZN (n_136_46), .A (n_140_44), .B (n_140_47), .C1 (n_144_45), .C2 (n_144_44) );
AOI211_X1 g_134_47 (.ZN (n_134_47), .A (n_138_45), .B (n_138_48), .C1 (n_142_46), .C2 (n_143_46) );
AOI211_X1 g_132_48 (.ZN (n_132_48), .A (n_136_46), .B (n_139_46), .C1 (n_140_47), .C2 (n_145_47) );
AOI211_X1 g_130_49 (.ZN (n_130_49), .A (n_134_47), .B (n_140_44), .C1 (n_138_48), .C2 (n_144_45) );
AOI211_X1 g_128_50 (.ZN (n_128_50), .A (n_132_48), .B (n_138_45), .C1 (n_139_46), .C2 (n_142_46) );
AOI211_X1 g_126_51 (.ZN (n_126_51), .A (n_130_49), .B (n_136_46), .C1 (n_140_44), .C2 (n_140_47) );
AOI211_X1 g_124_52 (.ZN (n_124_52), .A (n_128_50), .B (n_134_47), .C1 (n_138_45), .C2 (n_138_48) );
AOI211_X1 g_122_53 (.ZN (n_122_53), .A (n_126_51), .B (n_132_48), .C1 (n_136_46), .C2 (n_139_46) );
AOI211_X1 g_120_54 (.ZN (n_120_54), .A (n_124_52), .B (n_130_49), .C1 (n_134_47), .C2 (n_140_44) );
AOI211_X1 g_118_55 (.ZN (n_118_55), .A (n_122_53), .B (n_128_50), .C1 (n_132_48), .C2 (n_138_45) );
AOI211_X1 g_116_56 (.ZN (n_116_56), .A (n_120_54), .B (n_126_51), .C1 (n_130_49), .C2 (n_136_46) );
AOI211_X1 g_114_57 (.ZN (n_114_57), .A (n_118_55), .B (n_124_52), .C1 (n_128_50), .C2 (n_134_47) );
AOI211_X1 g_112_58 (.ZN (n_112_58), .A (n_116_56), .B (n_122_53), .C1 (n_126_51), .C2 (n_132_48) );
AOI211_X1 g_110_59 (.ZN (n_110_59), .A (n_114_57), .B (n_120_54), .C1 (n_124_52), .C2 (n_130_49) );
AOI211_X1 g_112_60 (.ZN (n_112_60), .A (n_112_58), .B (n_118_55), .C1 (n_122_53), .C2 (n_128_50) );
AOI211_X1 g_111_58 (.ZN (n_111_58), .A (n_110_59), .B (n_116_56), .C1 (n_120_54), .C2 (n_126_51) );
AOI211_X1 g_109_59 (.ZN (n_109_59), .A (n_112_60), .B (n_114_57), .C1 (n_118_55), .C2 (n_124_52) );
AOI211_X1 g_107_60 (.ZN (n_107_60), .A (n_111_58), .B (n_112_58), .C1 (n_116_56), .C2 (n_122_53) );
AOI211_X1 g_109_61 (.ZN (n_109_61), .A (n_109_59), .B (n_110_59), .C1 (n_114_57), .C2 (n_120_54) );
AOI211_X1 g_111_60 (.ZN (n_111_60), .A (n_107_60), .B (n_112_60), .C1 (n_112_58), .C2 (n_118_55) );
AOI211_X1 g_113_59 (.ZN (n_113_59), .A (n_109_61), .B (n_111_58), .C1 (n_110_59), .C2 (n_116_56) );
AOI211_X1 g_115_58 (.ZN (n_115_58), .A (n_111_60), .B (n_109_59), .C1 (n_112_60), .C2 (n_114_57) );
AOI211_X1 g_117_57 (.ZN (n_117_57), .A (n_113_59), .B (n_107_60), .C1 (n_111_58), .C2 (n_112_58) );
AOI211_X1 g_119_56 (.ZN (n_119_56), .A (n_115_58), .B (n_109_61), .C1 (n_109_59), .C2 (n_110_59) );
AOI211_X1 g_121_55 (.ZN (n_121_55), .A (n_117_57), .B (n_111_60), .C1 (n_107_60), .C2 (n_112_60) );
AOI211_X1 g_123_54 (.ZN (n_123_54), .A (n_119_56), .B (n_113_59), .C1 (n_109_61), .C2 (n_111_58) );
AOI211_X1 g_125_53 (.ZN (n_125_53), .A (n_121_55), .B (n_115_58), .C1 (n_111_60), .C2 (n_109_59) );
AOI211_X1 g_127_52 (.ZN (n_127_52), .A (n_123_54), .B (n_117_57), .C1 (n_113_59), .C2 (n_107_60) );
AOI211_X1 g_129_51 (.ZN (n_129_51), .A (n_125_53), .B (n_119_56), .C1 (n_115_58), .C2 (n_109_61) );
AOI211_X1 g_131_50 (.ZN (n_131_50), .A (n_127_52), .B (n_121_55), .C1 (n_117_57), .C2 (n_111_60) );
AOI211_X1 g_133_49 (.ZN (n_133_49), .A (n_129_51), .B (n_123_54), .C1 (n_119_56), .C2 (n_113_59) );
AOI211_X1 g_135_48 (.ZN (n_135_48), .A (n_131_50), .B (n_125_53), .C1 (n_121_55), .C2 (n_115_58) );
AOI211_X1 g_137_47 (.ZN (n_137_47), .A (n_133_49), .B (n_127_52), .C1 (n_123_54), .C2 (n_117_57) );
AOI211_X1 g_136_49 (.ZN (n_136_49), .A (n_135_48), .B (n_129_51), .C1 (n_125_53), .C2 (n_119_56) );
AOI211_X1 g_134_48 (.ZN (n_134_48), .A (n_137_47), .B (n_131_50), .C1 (n_127_52), .C2 (n_121_55) );
AOI211_X1 g_132_49 (.ZN (n_132_49), .A (n_136_49), .B (n_133_49), .C1 (n_129_51), .C2 (n_123_54) );
AOI211_X1 g_130_50 (.ZN (n_130_50), .A (n_134_48), .B (n_135_48), .C1 (n_131_50), .C2 (n_125_53) );
AOI211_X1 g_128_51 (.ZN (n_128_51), .A (n_132_49), .B (n_137_47), .C1 (n_133_49), .C2 (n_127_52) );
AOI211_X1 g_126_52 (.ZN (n_126_52), .A (n_130_50), .B (n_136_49), .C1 (n_135_48), .C2 (n_129_51) );
AOI211_X1 g_124_53 (.ZN (n_124_53), .A (n_128_51), .B (n_134_48), .C1 (n_137_47), .C2 (n_131_50) );
AOI211_X1 g_122_54 (.ZN (n_122_54), .A (n_126_52), .B (n_132_49), .C1 (n_136_49), .C2 (n_133_49) );
AOI211_X1 g_120_55 (.ZN (n_120_55), .A (n_124_53), .B (n_130_50), .C1 (n_134_48), .C2 (n_135_48) );
AOI211_X1 g_118_56 (.ZN (n_118_56), .A (n_122_54), .B (n_128_51), .C1 (n_132_49), .C2 (n_137_47) );
AOI211_X1 g_116_57 (.ZN (n_116_57), .A (n_120_55), .B (n_126_52), .C1 (n_130_50), .C2 (n_136_49) );
AOI211_X1 g_114_58 (.ZN (n_114_58), .A (n_118_56), .B (n_124_53), .C1 (n_128_51), .C2 (n_134_48) );
AOI211_X1 g_112_59 (.ZN (n_112_59), .A (n_116_57), .B (n_122_54), .C1 (n_126_52), .C2 (n_132_49) );
AOI211_X1 g_110_60 (.ZN (n_110_60), .A (n_114_58), .B (n_120_55), .C1 (n_124_53), .C2 (n_130_50) );
AOI211_X1 g_109_58 (.ZN (n_109_58), .A (n_112_59), .B (n_118_56), .C1 (n_122_54), .C2 (n_128_51) );
AOI211_X1 g_111_59 (.ZN (n_111_59), .A (n_110_60), .B (n_116_57), .C1 (n_120_55), .C2 (n_126_52) );
AOI211_X1 g_110_61 (.ZN (n_110_61), .A (n_109_58), .B (n_114_58), .C1 (n_118_56), .C2 (n_124_53) );
AOI211_X1 g_108_60 (.ZN (n_108_60), .A (n_111_59), .B (n_112_59), .C1 (n_116_57), .C2 (n_122_54) );
AOI211_X1 g_106_59 (.ZN (n_106_59), .A (n_110_61), .B (n_110_60), .C1 (n_114_58), .C2 (n_120_55) );
AOI211_X1 g_104_60 (.ZN (n_104_60), .A (n_108_60), .B (n_109_58), .C1 (n_112_59), .C2 (n_118_56) );
AOI211_X1 g_105_58 (.ZN (n_105_58), .A (n_106_59), .B (n_111_59), .C1 (n_110_60), .C2 (n_116_57) );
AOI211_X1 g_107_59 (.ZN (n_107_59), .A (n_104_60), .B (n_110_61), .C1 (n_109_58), .C2 (n_114_58) );
AOI211_X1 g_106_61 (.ZN (n_106_61), .A (n_105_58), .B (n_108_60), .C1 (n_111_59), .C2 (n_112_59) );
AOI211_X1 g_108_62 (.ZN (n_108_62), .A (n_107_59), .B (n_106_59), .C1 (n_110_61), .C2 (n_110_60) );
AOI211_X1 g_110_63 (.ZN (n_110_63), .A (n_106_61), .B (n_104_60), .C1 (n_108_60), .C2 (n_109_58) );
AOI211_X1 g_111_61 (.ZN (n_111_61), .A (n_108_62), .B (n_105_58), .C1 (n_106_59), .C2 (n_111_59) );
AOI211_X1 g_113_60 (.ZN (n_113_60), .A (n_110_63), .B (n_107_59), .C1 (n_104_60), .C2 (n_110_61) );
AOI211_X1 g_115_59 (.ZN (n_115_59), .A (n_111_61), .B (n_106_61), .C1 (n_105_58), .C2 (n_108_60) );
AOI211_X1 g_117_58 (.ZN (n_117_58), .A (n_113_60), .B (n_108_62), .C1 (n_107_59), .C2 (n_106_59) );
AOI211_X1 g_119_57 (.ZN (n_119_57), .A (n_115_59), .B (n_110_63), .C1 (n_106_61), .C2 (n_104_60) );
AOI211_X1 g_121_56 (.ZN (n_121_56), .A (n_117_58), .B (n_111_61), .C1 (n_108_62), .C2 (n_105_58) );
AOI211_X1 g_123_55 (.ZN (n_123_55), .A (n_119_57), .B (n_113_60), .C1 (n_110_63), .C2 (n_107_59) );
AOI211_X1 g_125_54 (.ZN (n_125_54), .A (n_121_56), .B (n_115_59), .C1 (n_111_61), .C2 (n_106_61) );
AOI211_X1 g_127_53 (.ZN (n_127_53), .A (n_123_55), .B (n_117_58), .C1 (n_113_60), .C2 (n_108_62) );
AOI211_X1 g_129_52 (.ZN (n_129_52), .A (n_125_54), .B (n_119_57), .C1 (n_115_59), .C2 (n_110_63) );
AOI211_X1 g_131_51 (.ZN (n_131_51), .A (n_127_53), .B (n_121_56), .C1 (n_117_58), .C2 (n_111_61) );
AOI211_X1 g_133_50 (.ZN (n_133_50), .A (n_129_52), .B (n_123_55), .C1 (n_119_57), .C2 (n_113_60) );
AOI211_X1 g_135_49 (.ZN (n_135_49), .A (n_131_51), .B (n_125_54), .C1 (n_121_56), .C2 (n_115_59) );
AOI211_X1 g_137_48 (.ZN (n_137_48), .A (n_133_50), .B (n_127_53), .C1 (n_123_55), .C2 (n_117_58) );
AOI211_X1 g_139_47 (.ZN (n_139_47), .A (n_135_49), .B (n_129_52), .C1 (n_125_54), .C2 (n_119_57) );
AOI211_X1 g_141_46 (.ZN (n_141_46), .A (n_137_48), .B (n_131_51), .C1 (n_127_53), .C2 (n_121_56) );
AOI211_X1 g_143_45 (.ZN (n_143_45), .A (n_139_47), .B (n_133_50), .C1 (n_129_52), .C2 (n_123_55) );
AOI211_X1 g_145_44 (.ZN (n_145_44), .A (n_141_46), .B (n_135_49), .C1 (n_131_51), .C2 (n_125_54) );
AOI211_X1 g_147_45 (.ZN (n_147_45), .A (n_143_45), .B (n_137_48), .C1 (n_133_50), .C2 (n_127_53) );
AOI211_X1 g_145_46 (.ZN (n_145_46), .A (n_145_44), .B (n_139_47), .C1 (n_135_49), .C2 (n_129_52) );
AOI211_X1 g_143_47 (.ZN (n_143_47), .A (n_147_45), .B (n_141_46), .C1 (n_137_48), .C2 (n_131_51) );
AOI211_X1 g_142_45 (.ZN (n_142_45), .A (n_145_46), .B (n_143_45), .C1 (n_139_47), .C2 (n_133_50) );
AOI211_X1 g_140_46 (.ZN (n_140_46), .A (n_143_47), .B (n_145_44), .C1 (n_141_46), .C2 (n_135_49) );
AOI211_X1 g_138_47 (.ZN (n_138_47), .A (n_142_45), .B (n_147_45), .C1 (n_143_45), .C2 (n_137_48) );
AOI211_X1 g_136_48 (.ZN (n_136_48), .A (n_140_46), .B (n_145_46), .C1 (n_145_44), .C2 (n_139_47) );
AOI211_X1 g_134_49 (.ZN (n_134_49), .A (n_138_47), .B (n_143_47), .C1 (n_147_45), .C2 (n_141_46) );
AOI211_X1 g_132_50 (.ZN (n_132_50), .A (n_136_48), .B (n_142_45), .C1 (n_145_46), .C2 (n_143_45) );
AOI211_X1 g_130_51 (.ZN (n_130_51), .A (n_134_49), .B (n_140_46), .C1 (n_143_47), .C2 (n_145_44) );
AOI211_X1 g_128_52 (.ZN (n_128_52), .A (n_132_50), .B (n_138_47), .C1 (n_142_45), .C2 (n_147_45) );
AOI211_X1 g_126_53 (.ZN (n_126_53), .A (n_130_51), .B (n_136_48), .C1 (n_140_46), .C2 (n_145_46) );
AOI211_X1 g_124_54 (.ZN (n_124_54), .A (n_128_52), .B (n_134_49), .C1 (n_138_47), .C2 (n_143_47) );
AOI211_X1 g_122_55 (.ZN (n_122_55), .A (n_126_53), .B (n_132_50), .C1 (n_136_48), .C2 (n_142_45) );
AOI211_X1 g_120_56 (.ZN (n_120_56), .A (n_124_54), .B (n_130_51), .C1 (n_134_49), .C2 (n_140_46) );
AOI211_X1 g_118_57 (.ZN (n_118_57), .A (n_122_55), .B (n_128_52), .C1 (n_132_50), .C2 (n_138_47) );
AOI211_X1 g_116_58 (.ZN (n_116_58), .A (n_120_56), .B (n_126_53), .C1 (n_130_51), .C2 (n_136_48) );
AOI211_X1 g_115_60 (.ZN (n_115_60), .A (n_118_57), .B (n_124_54), .C1 (n_128_52), .C2 (n_134_49) );
AOI211_X1 g_117_59 (.ZN (n_117_59), .A (n_116_58), .B (n_122_55), .C1 (n_126_53), .C2 (n_132_50) );
AOI211_X1 g_119_58 (.ZN (n_119_58), .A (n_115_60), .B (n_120_56), .C1 (n_124_54), .C2 (n_130_51) );
AOI211_X1 g_121_57 (.ZN (n_121_57), .A (n_117_59), .B (n_118_57), .C1 (n_122_55), .C2 (n_128_52) );
AOI211_X1 g_123_56 (.ZN (n_123_56), .A (n_119_58), .B (n_116_58), .C1 (n_120_56), .C2 (n_126_53) );
AOI211_X1 g_125_55 (.ZN (n_125_55), .A (n_121_57), .B (n_115_60), .C1 (n_118_57), .C2 (n_124_54) );
AOI211_X1 g_127_54 (.ZN (n_127_54), .A (n_123_56), .B (n_117_59), .C1 (n_116_58), .C2 (n_122_55) );
AOI211_X1 g_129_53 (.ZN (n_129_53), .A (n_125_55), .B (n_119_58), .C1 (n_115_60), .C2 (n_120_56) );
AOI211_X1 g_131_52 (.ZN (n_131_52), .A (n_127_54), .B (n_121_57), .C1 (n_117_59), .C2 (n_118_57) );
AOI211_X1 g_133_51 (.ZN (n_133_51), .A (n_129_53), .B (n_123_56), .C1 (n_119_58), .C2 (n_116_58) );
AOI211_X1 g_135_50 (.ZN (n_135_50), .A (n_131_52), .B (n_125_55), .C1 (n_121_57), .C2 (n_115_60) );
AOI211_X1 g_137_49 (.ZN (n_137_49), .A (n_133_51), .B (n_127_54), .C1 (n_123_56), .C2 (n_117_59) );
AOI211_X1 g_139_48 (.ZN (n_139_48), .A (n_135_50), .B (n_129_53), .C1 (n_125_55), .C2 (n_119_58) );
AOI211_X1 g_141_47 (.ZN (n_141_47), .A (n_137_49), .B (n_131_52), .C1 (n_127_54), .C2 (n_121_57) );
AOI211_X1 g_140_49 (.ZN (n_140_49), .A (n_139_48), .B (n_133_51), .C1 (n_129_53), .C2 (n_123_56) );
AOI211_X1 g_142_48 (.ZN (n_142_48), .A (n_141_47), .B (n_135_50), .C1 (n_131_52), .C2 (n_125_55) );
AOI211_X1 g_144_47 (.ZN (n_144_47), .A (n_140_49), .B (n_137_49), .C1 (n_133_51), .C2 (n_127_54) );
AOI211_X1 g_146_46 (.ZN (n_146_46), .A (n_142_48), .B (n_139_48), .C1 (n_135_50), .C2 (n_129_53) );
AOI211_X1 g_147_48 (.ZN (n_147_48), .A (n_144_47), .B (n_141_47), .C1 (n_137_49), .C2 (n_131_52) );
AOI211_X1 g_149_49 (.ZN (n_149_49), .A (n_146_46), .B (n_140_49), .C1 (n_139_48), .C2 (n_133_51) );
AOI211_X1 g_148_47 (.ZN (n_148_47), .A (n_147_48), .B (n_142_48), .C1 (n_141_47), .C2 (n_135_50) );
AOI211_X1 g_146_48 (.ZN (n_146_48), .A (n_149_49), .B (n_144_47), .C1 (n_140_49), .C2 (n_137_49) );
AOI211_X1 g_147_50 (.ZN (n_147_50), .A (n_148_47), .B (n_146_46), .C1 (n_142_48), .C2 (n_139_48) );
AOI211_X1 g_145_49 (.ZN (n_145_49), .A (n_146_48), .B (n_147_48), .C1 (n_144_47), .C2 (n_141_47) );
AOI211_X1 g_146_47 (.ZN (n_146_47), .A (n_147_50), .B (n_149_49), .C1 (n_146_46), .C2 (n_140_49) );
AOI211_X1 g_144_46 (.ZN (n_144_46), .A (n_145_49), .B (n_148_47), .C1 (n_147_48), .C2 (n_142_48) );
AOI211_X1 g_143_48 (.ZN (n_143_48), .A (n_146_47), .B (n_146_48), .C1 (n_149_49), .C2 (n_144_47) );
AOI211_X1 g_141_49 (.ZN (n_141_49), .A (n_144_46), .B (n_147_50), .C1 (n_148_47), .C2 (n_146_46) );
AOI211_X1 g_142_47 (.ZN (n_142_47), .A (n_143_48), .B (n_145_49), .C1 (n_146_48), .C2 (n_147_48) );
AOI211_X1 g_144_48 (.ZN (n_144_48), .A (n_141_49), .B (n_146_47), .C1 (n_147_50), .C2 (n_149_49) );
AOI211_X1 g_143_50 (.ZN (n_143_50), .A (n_142_47), .B (n_144_46), .C1 (n_145_49), .C2 (n_148_47) );
AOI211_X1 g_145_51 (.ZN (n_145_51), .A (n_144_48), .B (n_143_48), .C1 (n_146_47), .C2 (n_146_48) );
AOI211_X1 g_144_49 (.ZN (n_144_49), .A (n_143_50), .B (n_141_49), .C1 (n_144_46), .C2 (n_147_50) );
AOI211_X1 g_142_50 (.ZN (n_142_50), .A (n_145_51), .B (n_142_47), .C1 (n_143_48), .C2 (n_145_49) );
AOI211_X1 g_141_48 (.ZN (n_141_48), .A (n_144_49), .B (n_144_48), .C1 (n_141_49), .C2 (n_146_47) );
AOI211_X1 g_139_49 (.ZN (n_139_49), .A (n_142_50), .B (n_143_50), .C1 (n_142_47), .C2 (n_144_46) );
AOI211_X1 g_137_50 (.ZN (n_137_50), .A (n_141_48), .B (n_145_51), .C1 (n_144_48), .C2 (n_143_48) );
AOI211_X1 g_135_51 (.ZN (n_135_51), .A (n_139_49), .B (n_144_49), .C1 (n_143_50), .C2 (n_141_49) );
AOI211_X1 g_133_52 (.ZN (n_133_52), .A (n_137_50), .B (n_142_50), .C1 (n_145_51), .C2 (n_142_47) );
AOI211_X1 g_134_50 (.ZN (n_134_50), .A (n_135_51), .B (n_141_48), .C1 (n_144_49), .C2 (n_144_48) );
AOI211_X1 g_132_51 (.ZN (n_132_51), .A (n_133_52), .B (n_139_49), .C1 (n_142_50), .C2 (n_143_50) );
AOI211_X1 g_130_52 (.ZN (n_130_52), .A (n_134_50), .B (n_137_50), .C1 (n_141_48), .C2 (n_145_51) );
AOI211_X1 g_128_53 (.ZN (n_128_53), .A (n_132_51), .B (n_135_51), .C1 (n_139_49), .C2 (n_144_49) );
AOI211_X1 g_126_54 (.ZN (n_126_54), .A (n_130_52), .B (n_133_52), .C1 (n_137_50), .C2 (n_142_50) );
AOI211_X1 g_124_55 (.ZN (n_124_55), .A (n_128_53), .B (n_134_50), .C1 (n_135_51), .C2 (n_141_48) );
AOI211_X1 g_122_56 (.ZN (n_122_56), .A (n_126_54), .B (n_132_51), .C1 (n_133_52), .C2 (n_139_49) );
AOI211_X1 g_120_57 (.ZN (n_120_57), .A (n_124_55), .B (n_130_52), .C1 (n_134_50), .C2 (n_137_50) );
AOI211_X1 g_118_58 (.ZN (n_118_58), .A (n_122_56), .B (n_128_53), .C1 (n_132_51), .C2 (n_135_51) );
AOI211_X1 g_116_59 (.ZN (n_116_59), .A (n_120_57), .B (n_126_54), .C1 (n_130_52), .C2 (n_133_52) );
AOI211_X1 g_114_60 (.ZN (n_114_60), .A (n_118_58), .B (n_124_55), .C1 (n_128_53), .C2 (n_134_50) );
AOI211_X1 g_112_61 (.ZN (n_112_61), .A (n_116_59), .B (n_122_56), .C1 (n_126_54), .C2 (n_132_51) );
AOI211_X1 g_110_62 (.ZN (n_110_62), .A (n_114_60), .B (n_120_57), .C1 (n_124_55), .C2 (n_130_52) );
AOI211_X1 g_108_61 (.ZN (n_108_61), .A (n_112_61), .B (n_118_58), .C1 (n_122_56), .C2 (n_128_53) );
AOI211_X1 g_106_60 (.ZN (n_106_60), .A (n_110_62), .B (n_116_59), .C1 (n_120_57), .C2 (n_126_54) );
AOI211_X1 g_104_59 (.ZN (n_104_59), .A (n_108_61), .B (n_114_60), .C1 (n_118_58), .C2 (n_124_55) );
AOI211_X1 g_102_60 (.ZN (n_102_60), .A (n_106_60), .B (n_112_61), .C1 (n_116_59), .C2 (n_122_56) );
AOI211_X1 g_100_61 (.ZN (n_100_61), .A (n_104_59), .B (n_110_62), .C1 (n_114_60), .C2 (n_120_57) );
AOI211_X1 g_99_63 (.ZN (n_99_63), .A (n_102_60), .B (n_108_61), .C1 (n_112_61), .C2 (n_118_58) );
AOI211_X1 g_97_62 (.ZN (n_97_62), .A (n_100_61), .B (n_106_60), .C1 (n_110_62), .C2 (n_116_59) );
AOI211_X1 g_99_61 (.ZN (n_99_61), .A (n_99_63), .B (n_104_59), .C1 (n_108_61), .C2 (n_114_60) );
AOI211_X1 g_101_60 (.ZN (n_101_60), .A (n_97_62), .B (n_102_60), .C1 (n_106_60), .C2 (n_112_61) );
AOI211_X1 g_103_59 (.ZN (n_103_59), .A (n_99_61), .B (n_100_61), .C1 (n_104_59), .C2 (n_110_62) );
AOI211_X1 g_102_61 (.ZN (n_102_61), .A (n_101_60), .B (n_99_63), .C1 (n_102_60), .C2 (n_108_61) );
AOI211_X1 g_100_62 (.ZN (n_100_62), .A (n_103_59), .B (n_97_62), .C1 (n_100_61), .C2 (n_106_60) );
AOI211_X1 g_98_63 (.ZN (n_98_63), .A (n_102_61), .B (n_99_61), .C1 (n_99_63), .C2 (n_104_59) );
AOI211_X1 g_96_64 (.ZN (n_96_64), .A (n_100_62), .B (n_101_60), .C1 (n_97_62), .C2 (n_102_60) );
AOI211_X1 g_94_65 (.ZN (n_94_65), .A (n_98_63), .B (n_103_59), .C1 (n_99_61), .C2 (n_100_61) );
AOI211_X1 g_95_63 (.ZN (n_95_63), .A (n_96_64), .B (n_102_61), .C1 (n_101_60), .C2 (n_99_63) );
AOI211_X1 g_93_64 (.ZN (n_93_64), .A (n_94_65), .B (n_100_62), .C1 (n_103_59), .C2 (n_97_62) );
AOI211_X1 g_91_65 (.ZN (n_91_65), .A (n_95_63), .B (n_98_63), .C1 (n_102_61), .C2 (n_99_61) );
AOI211_X1 g_89_66 (.ZN (n_89_66), .A (n_93_64), .B (n_96_64), .C1 (n_100_62), .C2 (n_101_60) );
AOI211_X1 g_87_67 (.ZN (n_87_67), .A (n_91_65), .B (n_94_65), .C1 (n_98_63), .C2 (n_103_59) );
AOI211_X1 g_85_68 (.ZN (n_85_68), .A (n_89_66), .B (n_95_63), .C1 (n_96_64), .C2 (n_102_61) );
AOI211_X1 g_83_69 (.ZN (n_83_69), .A (n_87_67), .B (n_93_64), .C1 (n_94_65), .C2 (n_100_62) );
AOI211_X1 g_81_70 (.ZN (n_81_70), .A (n_85_68), .B (n_91_65), .C1 (n_95_63), .C2 (n_98_63) );
AOI211_X1 g_79_71 (.ZN (n_79_71), .A (n_83_69), .B (n_89_66), .C1 (n_93_64), .C2 (n_96_64) );
AOI211_X1 g_77_72 (.ZN (n_77_72), .A (n_81_70), .B (n_87_67), .C1 (n_91_65), .C2 (n_94_65) );
AOI211_X1 g_75_73 (.ZN (n_75_73), .A (n_79_71), .B (n_85_68), .C1 (n_89_66), .C2 (n_95_63) );
AOI211_X1 g_73_74 (.ZN (n_73_74), .A (n_77_72), .B (n_83_69), .C1 (n_87_67), .C2 (n_93_64) );
AOI211_X1 g_71_75 (.ZN (n_71_75), .A (n_75_73), .B (n_81_70), .C1 (n_85_68), .C2 (n_91_65) );
AOI211_X1 g_69_76 (.ZN (n_69_76), .A (n_73_74), .B (n_79_71), .C1 (n_83_69), .C2 (n_89_66) );
AOI211_X1 g_67_77 (.ZN (n_67_77), .A (n_71_75), .B (n_77_72), .C1 (n_81_70), .C2 (n_87_67) );
AOI211_X1 g_66_79 (.ZN (n_66_79), .A (n_69_76), .B (n_75_73), .C1 (n_79_71), .C2 (n_85_68) );
AOI211_X1 g_68_78 (.ZN (n_68_78), .A (n_67_77), .B (n_73_74), .C1 (n_77_72), .C2 (n_83_69) );
AOI211_X1 g_70_77 (.ZN (n_70_77), .A (n_66_79), .B (n_71_75), .C1 (n_75_73), .C2 (n_81_70) );
AOI211_X1 g_72_76 (.ZN (n_72_76), .A (n_68_78), .B (n_69_76), .C1 (n_73_74), .C2 (n_79_71) );
AOI211_X1 g_74_75 (.ZN (n_74_75), .A (n_70_77), .B (n_67_77), .C1 (n_71_75), .C2 (n_77_72) );
AOI211_X1 g_76_74 (.ZN (n_76_74), .A (n_72_76), .B (n_66_79), .C1 (n_69_76), .C2 (n_75_73) );
AOI211_X1 g_78_73 (.ZN (n_78_73), .A (n_74_75), .B (n_68_78), .C1 (n_67_77), .C2 (n_73_74) );
AOI211_X1 g_80_72 (.ZN (n_80_72), .A (n_76_74), .B (n_70_77), .C1 (n_66_79), .C2 (n_71_75) );
AOI211_X1 g_82_71 (.ZN (n_82_71), .A (n_78_73), .B (n_72_76), .C1 (n_68_78), .C2 (n_69_76) );
AOI211_X1 g_84_70 (.ZN (n_84_70), .A (n_80_72), .B (n_74_75), .C1 (n_70_77), .C2 (n_67_77) );
AOI211_X1 g_86_69 (.ZN (n_86_69), .A (n_82_71), .B (n_76_74), .C1 (n_72_76), .C2 (n_66_79) );
AOI211_X1 g_88_68 (.ZN (n_88_68), .A (n_84_70), .B (n_78_73), .C1 (n_74_75), .C2 (n_68_78) );
AOI211_X1 g_90_67 (.ZN (n_90_67), .A (n_86_69), .B (n_80_72), .C1 (n_76_74), .C2 (n_70_77) );
AOI211_X1 g_92_66 (.ZN (n_92_66), .A (n_88_68), .B (n_82_71), .C1 (n_78_73), .C2 (n_72_76) );
AOI211_X1 g_91_68 (.ZN (n_91_68), .A (n_90_67), .B (n_84_70), .C1 (n_80_72), .C2 (n_74_75) );
AOI211_X1 g_89_67 (.ZN (n_89_67), .A (n_92_66), .B (n_86_69), .C1 (n_82_71), .C2 (n_76_74) );
AOI211_X1 g_91_66 (.ZN (n_91_66), .A (n_91_68), .B (n_88_68), .C1 (n_84_70), .C2 (n_78_73) );
AOI211_X1 g_93_65 (.ZN (n_93_65), .A (n_89_67), .B (n_90_67), .C1 (n_86_69), .C2 (n_80_72) );
AOI211_X1 g_95_64 (.ZN (n_95_64), .A (n_91_66), .B (n_92_66), .C1 (n_88_68), .C2 (n_82_71) );
AOI211_X1 g_97_63 (.ZN (n_97_63), .A (n_93_65), .B (n_91_68), .C1 (n_90_67), .C2 (n_84_70) );
AOI211_X1 g_96_65 (.ZN (n_96_65), .A (n_95_64), .B (n_89_67), .C1 (n_92_66), .C2 (n_86_69) );
AOI211_X1 g_98_64 (.ZN (n_98_64), .A (n_97_63), .B (n_91_66), .C1 (n_91_68), .C2 (n_88_68) );
AOI211_X1 g_100_63 (.ZN (n_100_63), .A (n_96_65), .B (n_93_65), .C1 (n_89_67), .C2 (n_90_67) );
AOI211_X1 g_102_62 (.ZN (n_102_62), .A (n_98_64), .B (n_95_64), .C1 (n_91_66), .C2 (n_92_66) );
AOI211_X1 g_104_61 (.ZN (n_104_61), .A (n_100_63), .B (n_97_63), .C1 (n_93_65), .C2 (n_91_68) );
AOI211_X1 g_106_62 (.ZN (n_106_62), .A (n_102_62), .B (n_96_65), .C1 (n_95_64), .C2 (n_89_67) );
AOI211_X1 g_105_60 (.ZN (n_105_60), .A (n_104_61), .B (n_98_64), .C1 (n_97_63), .C2 (n_91_66) );
AOI211_X1 g_103_61 (.ZN (n_103_61), .A (n_106_62), .B (n_100_63), .C1 (n_96_65), .C2 (n_93_65) );
AOI211_X1 g_101_62 (.ZN (n_101_62), .A (n_105_60), .B (n_102_62), .C1 (n_98_64), .C2 (n_95_64) );
AOI211_X1 g_100_64 (.ZN (n_100_64), .A (n_103_61), .B (n_104_61), .C1 (n_100_63), .C2 (n_97_63) );
AOI211_X1 g_102_63 (.ZN (n_102_63), .A (n_101_62), .B (n_106_62), .C1 (n_102_62), .C2 (n_96_65) );
AOI211_X1 g_104_62 (.ZN (n_104_62), .A (n_100_64), .B (n_105_60), .C1 (n_104_61), .C2 (n_98_64) );
AOI211_X1 g_103_64 (.ZN (n_103_64), .A (n_102_63), .B (n_103_61), .C1 (n_106_62), .C2 (n_100_63) );
AOI211_X1 g_101_63 (.ZN (n_101_63), .A (n_104_62), .B (n_101_62), .C1 (n_105_60), .C2 (n_102_62) );
AOI211_X1 g_103_62 (.ZN (n_103_62), .A (n_103_64), .B (n_100_64), .C1 (n_103_61), .C2 (n_104_61) );
AOI211_X1 g_105_61 (.ZN (n_105_61), .A (n_101_63), .B (n_102_63), .C1 (n_101_62), .C2 (n_106_62) );
AOI211_X1 g_104_63 (.ZN (n_104_63), .A (n_103_62), .B (n_104_62), .C1 (n_100_64), .C2 (n_105_60) );
AOI211_X1 g_102_64 (.ZN (n_102_64), .A (n_105_61), .B (n_103_64), .C1 (n_102_63), .C2 (n_103_61) );
AOI211_X1 g_100_65 (.ZN (n_100_65), .A (n_104_63), .B (n_101_63), .C1 (n_104_62), .C2 (n_101_62) );
AOI211_X1 g_98_66 (.ZN (n_98_66), .A (n_102_64), .B (n_103_62), .C1 (n_103_64), .C2 (n_100_64) );
AOI211_X1 g_99_64 (.ZN (n_99_64), .A (n_100_65), .B (n_105_61), .C1 (n_101_63), .C2 (n_102_63) );
AOI211_X1 g_97_65 (.ZN (n_97_65), .A (n_98_66), .B (n_104_63), .C1 (n_103_62), .C2 (n_104_62) );
AOI211_X1 g_95_66 (.ZN (n_95_66), .A (n_99_64), .B (n_102_64), .C1 (n_105_61), .C2 (n_103_64) );
AOI211_X1 g_93_67 (.ZN (n_93_67), .A (n_97_65), .B (n_100_65), .C1 (n_104_63), .C2 (n_101_63) );
AOI211_X1 g_92_69 (.ZN (n_92_69), .A (n_95_66), .B (n_98_66), .C1 (n_102_64), .C2 (n_103_62) );
AOI211_X1 g_91_67 (.ZN (n_91_67), .A (n_93_67), .B (n_99_64), .C1 (n_100_65), .C2 (n_105_61) );
AOI211_X1 g_93_66 (.ZN (n_93_66), .A (n_92_69), .B (n_97_65), .C1 (n_98_66), .C2 (n_104_63) );
AOI211_X1 g_95_65 (.ZN (n_95_65), .A (n_91_67), .B (n_95_66), .C1 (n_99_64), .C2 (n_102_64) );
AOI211_X1 g_97_64 (.ZN (n_97_64), .A (n_93_66), .B (n_93_67), .C1 (n_97_65), .C2 (n_100_65) );
AOI211_X1 g_96_66 (.ZN (n_96_66), .A (n_95_65), .B (n_92_69), .C1 (n_95_66), .C2 (n_98_66) );
AOI211_X1 g_98_65 (.ZN (n_98_65), .A (n_97_64), .B (n_91_67), .C1 (n_93_67), .C2 (n_99_64) );
AOI211_X1 g_97_67 (.ZN (n_97_67), .A (n_96_66), .B (n_93_66), .C1 (n_92_69), .C2 (n_97_65) );
AOI211_X1 g_99_66 (.ZN (n_99_66), .A (n_98_65), .B (n_95_65), .C1 (n_91_67), .C2 (n_95_66) );
AOI211_X1 g_101_65 (.ZN (n_101_65), .A (n_97_67), .B (n_97_64), .C1 (n_93_66), .C2 (n_93_67) );
AOI211_X1 g_100_67 (.ZN (n_100_67), .A (n_99_66), .B (n_96_66), .C1 (n_95_65), .C2 (n_92_69) );
AOI211_X1 g_99_65 (.ZN (n_99_65), .A (n_101_65), .B (n_98_65), .C1 (n_97_64), .C2 (n_91_67) );
AOI211_X1 g_101_64 (.ZN (n_101_64), .A (n_100_67), .B (n_97_67), .C1 (n_96_66), .C2 (n_93_66) );
AOI211_X1 g_103_63 (.ZN (n_103_63), .A (n_99_65), .B (n_99_66), .C1 (n_98_65), .C2 (n_95_65) );
AOI211_X1 g_105_62 (.ZN (n_105_62), .A (n_101_64), .B (n_101_65), .C1 (n_97_67), .C2 (n_97_64) );
AOI211_X1 g_107_61 (.ZN (n_107_61), .A (n_103_63), .B (n_100_67), .C1 (n_99_66), .C2 (n_96_66) );
AOI211_X1 g_106_63 (.ZN (n_106_63), .A (n_105_62), .B (n_99_65), .C1 (n_101_65), .C2 (n_98_65) );
AOI211_X1 g_104_64 (.ZN (n_104_64), .A (n_107_61), .B (n_101_64), .C1 (n_100_67), .C2 (n_97_67) );
AOI211_X1 g_102_65 (.ZN (n_102_65), .A (n_106_63), .B (n_103_63), .C1 (n_99_65), .C2 (n_99_66) );
AOI211_X1 g_100_66 (.ZN (n_100_66), .A (n_104_64), .B (n_105_62), .C1 (n_101_64), .C2 (n_101_65) );
AOI211_X1 g_98_67 (.ZN (n_98_67), .A (n_102_65), .B (n_107_61), .C1 (n_103_63), .C2 (n_100_67) );
AOI211_X1 g_96_68 (.ZN (n_96_68), .A (n_100_66), .B (n_106_63), .C1 (n_105_62), .C2 (n_99_65) );
AOI211_X1 g_97_66 (.ZN (n_97_66), .A (n_98_67), .B (n_104_64), .C1 (n_107_61), .C2 (n_101_64) );
AOI211_X1 g_95_67 (.ZN (n_95_67), .A (n_96_68), .B (n_102_65), .C1 (n_106_63), .C2 (n_103_63) );
AOI211_X1 g_93_68 (.ZN (n_93_68), .A (n_97_66), .B (n_100_66), .C1 (n_104_64), .C2 (n_105_62) );
AOI211_X1 g_94_66 (.ZN (n_94_66), .A (n_95_67), .B (n_98_67), .C1 (n_102_65), .C2 (n_107_61) );
AOI211_X1 g_92_67 (.ZN (n_92_67), .A (n_93_68), .B (n_96_68), .C1 (n_100_66), .C2 (n_106_63) );
AOI211_X1 g_90_68 (.ZN (n_90_68), .A (n_94_66), .B (n_97_66), .C1 (n_98_67), .C2 (n_104_64) );
AOI211_X1 g_88_69 (.ZN (n_88_69), .A (n_92_67), .B (n_95_67), .C1 (n_96_68), .C2 (n_102_65) );
AOI211_X1 g_86_70 (.ZN (n_86_70), .A (n_90_68), .B (n_93_68), .C1 (n_97_66), .C2 (n_100_66) );
AOI211_X1 g_87_68 (.ZN (n_87_68), .A (n_88_69), .B (n_94_66), .C1 (n_95_67), .C2 (n_98_67) );
AOI211_X1 g_85_69 (.ZN (n_85_69), .A (n_86_70), .B (n_92_67), .C1 (n_93_68), .C2 (n_96_68) );
AOI211_X1 g_83_70 (.ZN (n_83_70), .A (n_87_68), .B (n_90_68), .C1 (n_94_66), .C2 (n_97_66) );
AOI211_X1 g_81_71 (.ZN (n_81_71), .A (n_85_69), .B (n_88_69), .C1 (n_92_67), .C2 (n_95_67) );
AOI211_X1 g_79_72 (.ZN (n_79_72), .A (n_83_70), .B (n_86_70), .C1 (n_90_68), .C2 (n_93_68) );
AOI211_X1 g_77_73 (.ZN (n_77_73), .A (n_81_71), .B (n_87_68), .C1 (n_88_69), .C2 (n_94_66) );
AOI211_X1 g_75_74 (.ZN (n_75_74), .A (n_79_72), .B (n_85_69), .C1 (n_86_70), .C2 (n_92_67) );
AOI211_X1 g_73_75 (.ZN (n_73_75), .A (n_77_73), .B (n_83_70), .C1 (n_87_68), .C2 (n_90_68) );
AOI211_X1 g_71_76 (.ZN (n_71_76), .A (n_75_74), .B (n_81_71), .C1 (n_85_69), .C2 (n_88_69) );
AOI211_X1 g_69_77 (.ZN (n_69_77), .A (n_73_75), .B (n_79_72), .C1 (n_83_70), .C2 (n_86_70) );
AOI211_X1 g_67_78 (.ZN (n_67_78), .A (n_71_76), .B (n_77_73), .C1 (n_81_71), .C2 (n_87_68) );
AOI211_X1 g_65_79 (.ZN (n_65_79), .A (n_69_77), .B (n_75_74), .C1 (n_79_72), .C2 (n_85_69) );
AOI211_X1 g_63_80 (.ZN (n_63_80), .A (n_67_78), .B (n_73_75), .C1 (n_77_73), .C2 (n_83_70) );
AOI211_X1 g_61_81 (.ZN (n_61_81), .A (n_65_79), .B (n_71_76), .C1 (n_75_74), .C2 (n_81_71) );
AOI211_X1 g_59_80 (.ZN (n_59_80), .A (n_63_80), .B (n_69_77), .C1 (n_73_75), .C2 (n_79_72) );
AOI211_X1 g_57_81 (.ZN (n_57_81), .A (n_61_81), .B (n_67_78), .C1 (n_71_76), .C2 (n_77_73) );
AOI211_X1 g_55_82 (.ZN (n_55_82), .A (n_59_80), .B (n_65_79), .C1 (n_69_77), .C2 (n_75_74) );
AOI211_X1 g_53_83 (.ZN (n_53_83), .A (n_57_81), .B (n_63_80), .C1 (n_67_78), .C2 (n_73_75) );
AOI211_X1 g_51_84 (.ZN (n_51_84), .A (n_55_82), .B (n_61_81), .C1 (n_65_79), .C2 (n_71_76) );
AOI211_X1 g_49_85 (.ZN (n_49_85), .A (n_53_83), .B (n_59_80), .C1 (n_63_80), .C2 (n_69_77) );
AOI211_X1 g_47_86 (.ZN (n_47_86), .A (n_51_84), .B (n_57_81), .C1 (n_61_81), .C2 (n_67_78) );
AOI211_X1 g_45_87 (.ZN (n_45_87), .A (n_49_85), .B (n_55_82), .C1 (n_59_80), .C2 (n_65_79) );
AOI211_X1 g_43_88 (.ZN (n_43_88), .A (n_47_86), .B (n_53_83), .C1 (n_57_81), .C2 (n_63_80) );
AOI211_X1 g_41_89 (.ZN (n_41_89), .A (n_45_87), .B (n_51_84), .C1 (n_55_82), .C2 (n_61_81) );
AOI211_X1 g_39_90 (.ZN (n_39_90), .A (n_43_88), .B (n_49_85), .C1 (n_53_83), .C2 (n_59_80) );
AOI211_X1 g_37_91 (.ZN (n_37_91), .A (n_41_89), .B (n_47_86), .C1 (n_51_84), .C2 (n_57_81) );
AOI211_X1 g_35_92 (.ZN (n_35_92), .A (n_39_90), .B (n_45_87), .C1 (n_49_85), .C2 (n_55_82) );
AOI211_X1 g_36_90 (.ZN (n_36_90), .A (n_37_91), .B (n_43_88), .C1 (n_47_86), .C2 (n_53_83) );
AOI211_X1 g_34_91 (.ZN (n_34_91), .A (n_35_92), .B (n_41_89), .C1 (n_45_87), .C2 (n_51_84) );
AOI211_X1 g_33_93 (.ZN (n_33_93), .A (n_36_90), .B (n_39_90), .C1 (n_43_88), .C2 (n_49_85) );
AOI211_X1 g_31_94 (.ZN (n_31_94), .A (n_34_91), .B (n_37_91), .C1 (n_41_89), .C2 (n_47_86) );
AOI211_X1 g_32_92 (.ZN (n_32_92), .A (n_33_93), .B (n_35_92), .C1 (n_39_90), .C2 (n_45_87) );
AOI211_X1 g_33_90 (.ZN (n_33_90), .A (n_31_94), .B (n_36_90), .C1 (n_37_91), .C2 (n_43_88) );
AOI211_X1 g_31_91 (.ZN (n_31_91), .A (n_32_92), .B (n_34_91), .C1 (n_35_92), .C2 (n_41_89) );
AOI211_X1 g_29_92 (.ZN (n_29_92), .A (n_33_90), .B (n_33_93), .C1 (n_36_90), .C2 (n_39_90) );
AOI211_X1 g_28_94 (.ZN (n_28_94), .A (n_31_91), .B (n_31_94), .C1 (n_34_91), .C2 (n_37_91) );
AOI211_X1 g_30_93 (.ZN (n_30_93), .A (n_29_92), .B (n_32_92), .C1 (n_33_93), .C2 (n_35_92) );
AOI211_X1 g_29_95 (.ZN (n_29_95), .A (n_28_94), .B (n_33_90), .C1 (n_31_94), .C2 (n_36_90) );
AOI211_X1 g_27_94 (.ZN (n_27_94), .A (n_30_93), .B (n_31_91), .C1 (n_32_92), .C2 (n_34_91) );
AOI211_X1 g_25_95 (.ZN (n_25_95), .A (n_29_95), .B (n_29_92), .C1 (n_33_90), .C2 (n_33_93) );
AOI211_X1 g_23_96 (.ZN (n_23_96), .A (n_27_94), .B (n_28_94), .C1 (n_31_91), .C2 (n_31_94) );
AOI211_X1 g_21_97 (.ZN (n_21_97), .A (n_25_95), .B (n_30_93), .C1 (n_29_92), .C2 (n_32_92) );
AOI211_X1 g_23_98 (.ZN (n_23_98), .A (n_23_96), .B (n_29_95), .C1 (n_28_94), .C2 (n_33_90) );
AOI211_X1 g_25_97 (.ZN (n_25_97), .A (n_21_97), .B (n_27_94), .C1 (n_30_93), .C2 (n_31_91) );
AOI211_X1 g_27_96 (.ZN (n_27_96), .A (n_23_98), .B (n_25_95), .C1 (n_29_95), .C2 (n_29_92) );
AOI211_X1 g_26_98 (.ZN (n_26_98), .A (n_25_97), .B (n_23_96), .C1 (n_27_94), .C2 (n_28_94) );
AOI211_X1 g_25_96 (.ZN (n_25_96), .A (n_27_96), .B (n_21_97), .C1 (n_25_95), .C2 (n_30_93) );
AOI211_X1 g_23_95 (.ZN (n_23_95), .A (n_26_98), .B (n_23_98), .C1 (n_23_96), .C2 (n_29_95) );
AOI211_X1 g_25_94 (.ZN (n_25_94), .A (n_25_96), .B (n_25_97), .C1 (n_21_97), .C2 (n_27_94) );
AOI211_X1 g_24_96 (.ZN (n_24_96), .A (n_23_95), .B (n_27_96), .C1 (n_23_98), .C2 (n_25_95) );
AOI211_X1 g_26_95 (.ZN (n_26_95), .A (n_25_94), .B (n_26_98), .C1 (n_25_97), .C2 (n_23_96) );
AOI211_X1 g_27_97 (.ZN (n_27_97), .A (n_24_96), .B (n_25_96), .C1 (n_27_96), .C2 (n_21_97) );
AOI211_X1 g_28_95 (.ZN (n_28_95), .A (n_26_95), .B (n_23_95), .C1 (n_26_98), .C2 (n_23_98) );
AOI211_X1 g_30_94 (.ZN (n_30_94), .A (n_27_97), .B (n_25_94), .C1 (n_25_96), .C2 (n_25_97) );
AOI211_X1 g_32_93 (.ZN (n_32_93), .A (n_28_95), .B (n_24_96), .C1 (n_23_95), .C2 (n_27_96) );
AOI211_X1 g_34_92 (.ZN (n_34_92), .A (n_30_94), .B (n_26_95), .C1 (n_25_94), .C2 (n_26_98) );
AOI211_X1 g_36_91 (.ZN (n_36_91), .A (n_32_93), .B (n_27_97), .C1 (n_24_96), .C2 (n_25_96) );
AOI211_X1 g_38_90 (.ZN (n_38_90), .A (n_34_92), .B (n_28_95), .C1 (n_26_95), .C2 (n_23_95) );
AOI211_X1 g_40_89 (.ZN (n_40_89), .A (n_36_91), .B (n_30_94), .C1 (n_27_97), .C2 (n_25_94) );
AOI211_X1 g_42_88 (.ZN (n_42_88), .A (n_38_90), .B (n_32_93), .C1 (n_28_95), .C2 (n_24_96) );
AOI211_X1 g_44_87 (.ZN (n_44_87), .A (n_40_89), .B (n_34_92), .C1 (n_30_94), .C2 (n_26_95) );
AOI211_X1 g_46_86 (.ZN (n_46_86), .A (n_42_88), .B (n_36_91), .C1 (n_32_93), .C2 (n_27_97) );
AOI211_X1 g_48_85 (.ZN (n_48_85), .A (n_44_87), .B (n_38_90), .C1 (n_34_92), .C2 (n_28_95) );
AOI211_X1 g_50_84 (.ZN (n_50_84), .A (n_46_86), .B (n_40_89), .C1 (n_36_91), .C2 (n_30_94) );
AOI211_X1 g_52_83 (.ZN (n_52_83), .A (n_48_85), .B (n_42_88), .C1 (n_38_90), .C2 (n_32_93) );
AOI211_X1 g_54_82 (.ZN (n_54_82), .A (n_50_84), .B (n_44_87), .C1 (n_40_89), .C2 (n_34_92) );
AOI211_X1 g_53_84 (.ZN (n_53_84), .A (n_52_83), .B (n_46_86), .C1 (n_42_88), .C2 (n_36_91) );
AOI211_X1 g_51_85 (.ZN (n_51_85), .A (n_54_82), .B (n_48_85), .C1 (n_44_87), .C2 (n_38_90) );
AOI211_X1 g_49_86 (.ZN (n_49_86), .A (n_53_84), .B (n_50_84), .C1 (n_46_86), .C2 (n_40_89) );
AOI211_X1 g_47_87 (.ZN (n_47_87), .A (n_51_85), .B (n_52_83), .C1 (n_48_85), .C2 (n_42_88) );
AOI211_X1 g_45_88 (.ZN (n_45_88), .A (n_49_86), .B (n_54_82), .C1 (n_50_84), .C2 (n_44_87) );
AOI211_X1 g_43_87 (.ZN (n_43_87), .A (n_47_87), .B (n_53_84), .C1 (n_52_83), .C2 (n_46_86) );
AOI211_X1 g_41_88 (.ZN (n_41_88), .A (n_45_88), .B (n_51_85), .C1 (n_54_82), .C2 (n_48_85) );
AOI211_X1 g_39_89 (.ZN (n_39_89), .A (n_43_87), .B (n_49_86), .C1 (n_53_84), .C2 (n_50_84) );
AOI211_X1 g_38_91 (.ZN (n_38_91), .A (n_41_88), .B (n_47_87), .C1 (n_51_85), .C2 (n_52_83) );
AOI211_X1 g_40_90 (.ZN (n_40_90), .A (n_39_89), .B (n_45_88), .C1 (n_49_86), .C2 (n_54_82) );
AOI211_X1 g_42_89 (.ZN (n_42_89), .A (n_38_91), .B (n_43_87), .C1 (n_47_87), .C2 (n_53_84) );
AOI211_X1 g_44_88 (.ZN (n_44_88), .A (n_40_90), .B (n_41_88), .C1 (n_45_88), .C2 (n_51_85) );
AOI211_X1 g_46_87 (.ZN (n_46_87), .A (n_42_89), .B (n_39_89), .C1 (n_43_87), .C2 (n_49_86) );
AOI211_X1 g_48_86 (.ZN (n_48_86), .A (n_44_88), .B (n_38_91), .C1 (n_41_88), .C2 (n_47_87) );
AOI211_X1 g_47_88 (.ZN (n_47_88), .A (n_46_87), .B (n_40_90), .C1 (n_39_89), .C2 (n_45_88) );
AOI211_X1 g_49_87 (.ZN (n_49_87), .A (n_48_86), .B (n_42_89), .C1 (n_38_91), .C2 (n_43_87) );
AOI211_X1 g_51_86 (.ZN (n_51_86), .A (n_47_88), .B (n_44_88), .C1 (n_40_90), .C2 (n_41_88) );
AOI211_X1 g_53_85 (.ZN (n_53_85), .A (n_49_87), .B (n_46_87), .C1 (n_42_89), .C2 (n_39_89) );
AOI211_X1 g_55_84 (.ZN (n_55_84), .A (n_51_86), .B (n_48_86), .C1 (n_44_88), .C2 (n_38_91) );
AOI211_X1 g_57_83 (.ZN (n_57_83), .A (n_53_85), .B (n_47_88), .C1 (n_46_87), .C2 (n_40_90) );
AOI211_X1 g_59_82 (.ZN (n_59_82), .A (n_55_84), .B (n_49_87), .C1 (n_48_86), .C2 (n_42_89) );
AOI211_X1 g_58_84 (.ZN (n_58_84), .A (n_57_83), .B (n_51_86), .C1 (n_47_88), .C2 (n_44_88) );
AOI211_X1 g_56_83 (.ZN (n_56_83), .A (n_59_82), .B (n_53_85), .C1 (n_49_87), .C2 (n_46_87) );
AOI211_X1 g_58_82 (.ZN (n_58_82), .A (n_58_84), .B (n_55_84), .C1 (n_51_86), .C2 (n_48_86) );
AOI211_X1 g_60_81 (.ZN (n_60_81), .A (n_56_83), .B (n_57_83), .C1 (n_53_85), .C2 (n_47_88) );
AOI211_X1 g_62_80 (.ZN (n_62_80), .A (n_58_82), .B (n_59_82), .C1 (n_55_84), .C2 (n_49_87) );
AOI211_X1 g_64_79 (.ZN (n_64_79), .A (n_60_81), .B (n_58_84), .C1 (n_57_83), .C2 (n_51_86) );
AOI211_X1 g_63_81 (.ZN (n_63_81), .A (n_62_80), .B (n_56_83), .C1 (n_59_82), .C2 (n_53_85) );
AOI211_X1 g_65_80 (.ZN (n_65_80), .A (n_64_79), .B (n_58_82), .C1 (n_58_84), .C2 (n_55_84) );
AOI211_X1 g_67_79 (.ZN (n_67_79), .A (n_63_81), .B (n_60_81), .C1 (n_56_83), .C2 (n_57_83) );
AOI211_X1 g_69_78 (.ZN (n_69_78), .A (n_65_80), .B (n_62_80), .C1 (n_58_82), .C2 (n_59_82) );
AOI211_X1 g_71_77 (.ZN (n_71_77), .A (n_67_79), .B (n_64_79), .C1 (n_60_81), .C2 (n_58_84) );
AOI211_X1 g_73_76 (.ZN (n_73_76), .A (n_69_78), .B (n_63_81), .C1 (n_62_80), .C2 (n_56_83) );
AOI211_X1 g_75_75 (.ZN (n_75_75), .A (n_71_77), .B (n_65_80), .C1 (n_64_79), .C2 (n_58_82) );
AOI211_X1 g_77_74 (.ZN (n_77_74), .A (n_73_76), .B (n_67_79), .C1 (n_63_81), .C2 (n_60_81) );
AOI211_X1 g_79_73 (.ZN (n_79_73), .A (n_75_75), .B (n_69_78), .C1 (n_65_80), .C2 (n_62_80) );
AOI211_X1 g_81_72 (.ZN (n_81_72), .A (n_77_74), .B (n_71_77), .C1 (n_67_79), .C2 (n_64_79) );
AOI211_X1 g_83_71 (.ZN (n_83_71), .A (n_79_73), .B (n_73_76), .C1 (n_69_78), .C2 (n_63_81) );
AOI211_X1 g_85_70 (.ZN (n_85_70), .A (n_81_72), .B (n_75_75), .C1 (n_71_77), .C2 (n_65_80) );
AOI211_X1 g_87_69 (.ZN (n_87_69), .A (n_83_71), .B (n_77_74), .C1 (n_73_76), .C2 (n_67_79) );
AOI211_X1 g_89_68 (.ZN (n_89_68), .A (n_85_70), .B (n_79_73), .C1 (n_75_75), .C2 (n_69_78) );
AOI211_X1 g_90_70 (.ZN (n_90_70), .A (n_87_69), .B (n_81_72), .C1 (n_77_74), .C2 (n_71_77) );
AOI211_X1 g_88_71 (.ZN (n_88_71), .A (n_89_68), .B (n_83_71), .C1 (n_79_73), .C2 (n_73_76) );
AOI211_X1 g_89_69 (.ZN (n_89_69), .A (n_90_70), .B (n_85_70), .C1 (n_81_72), .C2 (n_75_75) );
AOI211_X1 g_87_70 (.ZN (n_87_70), .A (n_88_71), .B (n_87_69), .C1 (n_83_71), .C2 (n_77_74) );
AOI211_X1 g_85_71 (.ZN (n_85_71), .A (n_89_69), .B (n_89_68), .C1 (n_85_70), .C2 (n_79_73) );
AOI211_X1 g_83_72 (.ZN (n_83_72), .A (n_87_70), .B (n_90_70), .C1 (n_87_69), .C2 (n_81_72) );
AOI211_X1 g_81_73 (.ZN (n_81_73), .A (n_85_71), .B (n_88_71), .C1 (n_89_68), .C2 (n_83_71) );
AOI211_X1 g_79_74 (.ZN (n_79_74), .A (n_83_72), .B (n_89_69), .C1 (n_90_70), .C2 (n_85_70) );
AOI211_X1 g_77_75 (.ZN (n_77_75), .A (n_81_73), .B (n_87_70), .C1 (n_88_71), .C2 (n_87_69) );
AOI211_X1 g_75_76 (.ZN (n_75_76), .A (n_79_74), .B (n_85_71), .C1 (n_89_69), .C2 (n_89_68) );
AOI211_X1 g_73_77 (.ZN (n_73_77), .A (n_77_75), .B (n_83_72), .C1 (n_87_70), .C2 (n_90_70) );
AOI211_X1 g_71_78 (.ZN (n_71_78), .A (n_75_76), .B (n_81_73), .C1 (n_85_71), .C2 (n_88_71) );
AOI211_X1 g_69_79 (.ZN (n_69_79), .A (n_73_77), .B (n_79_74), .C1 (n_83_72), .C2 (n_89_69) );
AOI211_X1 g_67_80 (.ZN (n_67_80), .A (n_71_78), .B (n_77_75), .C1 (n_81_73), .C2 (n_87_70) );
AOI211_X1 g_65_81 (.ZN (n_65_81), .A (n_69_79), .B (n_75_76), .C1 (n_79_74), .C2 (n_85_71) );
AOI211_X1 g_63_82 (.ZN (n_63_82), .A (n_67_80), .B (n_73_77), .C1 (n_77_75), .C2 (n_83_72) );
AOI211_X1 g_64_80 (.ZN (n_64_80), .A (n_65_81), .B (n_71_78), .C1 (n_75_76), .C2 (n_81_73) );
AOI211_X1 g_62_81 (.ZN (n_62_81), .A (n_63_82), .B (n_69_79), .C1 (n_73_77), .C2 (n_79_74) );
AOI211_X1 g_60_82 (.ZN (n_60_82), .A (n_64_80), .B (n_67_80), .C1 (n_71_78), .C2 (n_77_75) );
AOI211_X1 g_58_83 (.ZN (n_58_83), .A (n_62_81), .B (n_65_81), .C1 (n_69_79), .C2 (n_75_76) );
AOI211_X1 g_56_84 (.ZN (n_56_84), .A (n_60_82), .B (n_63_82), .C1 (n_67_80), .C2 (n_73_77) );
AOI211_X1 g_54_85 (.ZN (n_54_85), .A (n_58_83), .B (n_64_80), .C1 (n_65_81), .C2 (n_71_78) );
AOI211_X1 g_52_86 (.ZN (n_52_86), .A (n_56_84), .B (n_62_81), .C1 (n_63_82), .C2 (n_69_79) );
AOI211_X1 g_50_87 (.ZN (n_50_87), .A (n_54_85), .B (n_60_82), .C1 (n_64_80), .C2 (n_67_80) );
AOI211_X1 g_48_88 (.ZN (n_48_88), .A (n_52_86), .B (n_58_83), .C1 (n_62_81), .C2 (n_65_81) );
AOI211_X1 g_46_89 (.ZN (n_46_89), .A (n_50_87), .B (n_56_84), .C1 (n_60_82), .C2 (n_63_82) );
AOI211_X1 g_44_90 (.ZN (n_44_90), .A (n_48_88), .B (n_54_85), .C1 (n_58_83), .C2 (n_64_80) );
AOI211_X1 g_42_91 (.ZN (n_42_91), .A (n_46_89), .B (n_52_86), .C1 (n_56_84), .C2 (n_62_81) );
AOI211_X1 g_43_89 (.ZN (n_43_89), .A (n_44_90), .B (n_50_87), .C1 (n_54_85), .C2 (n_60_82) );
AOI211_X1 g_41_90 (.ZN (n_41_90), .A (n_42_91), .B (n_48_88), .C1 (n_52_86), .C2 (n_58_83) );
AOI211_X1 g_39_91 (.ZN (n_39_91), .A (n_43_89), .B (n_46_89), .C1 (n_50_87), .C2 (n_56_84) );
AOI211_X1 g_37_92 (.ZN (n_37_92), .A (n_41_90), .B (n_44_90), .C1 (n_48_88), .C2 (n_54_85) );
AOI211_X1 g_35_91 (.ZN (n_35_91), .A (n_39_91), .B (n_42_91), .C1 (n_46_89), .C2 (n_52_86) );
AOI211_X1 g_33_92 (.ZN (n_33_92), .A (n_37_92), .B (n_43_89), .C1 (n_44_90), .C2 (n_50_87) );
AOI211_X1 g_31_93 (.ZN (n_31_93), .A (n_35_91), .B (n_41_90), .C1 (n_42_91), .C2 (n_48_88) );
AOI211_X1 g_29_94 (.ZN (n_29_94), .A (n_33_92), .B (n_39_91), .C1 (n_43_89), .C2 (n_46_89) );
AOI211_X1 g_27_95 (.ZN (n_27_95), .A (n_31_93), .B (n_37_92), .C1 (n_41_90), .C2 (n_44_90) );
AOI211_X1 g_29_96 (.ZN (n_29_96), .A (n_29_94), .B (n_35_91), .C1 (n_39_91), .C2 (n_42_91) );
AOI211_X1 g_31_95 (.ZN (n_31_95), .A (n_27_95), .B (n_33_92), .C1 (n_37_92), .C2 (n_43_89) );
AOI211_X1 g_33_94 (.ZN (n_33_94), .A (n_29_96), .B (n_31_93), .C1 (n_35_91), .C2 (n_41_90) );
AOI211_X1 g_35_93 (.ZN (n_35_93), .A (n_31_95), .B (n_29_94), .C1 (n_33_92), .C2 (n_39_91) );
AOI211_X1 g_34_95 (.ZN (n_34_95), .A (n_33_94), .B (n_27_95), .C1 (n_31_93), .C2 (n_37_92) );
AOI211_X1 g_32_94 (.ZN (n_32_94), .A (n_35_93), .B (n_29_96), .C1 (n_29_94), .C2 (n_35_91) );
AOI211_X1 g_34_93 (.ZN (n_34_93), .A (n_34_95), .B (n_31_95), .C1 (n_27_95), .C2 (n_33_92) );
AOI211_X1 g_36_92 (.ZN (n_36_92), .A (n_32_94), .B (n_33_94), .C1 (n_29_96), .C2 (n_31_93) );
AOI211_X1 g_35_94 (.ZN (n_35_94), .A (n_34_93), .B (n_35_93), .C1 (n_31_95), .C2 (n_29_94) );
AOI211_X1 g_37_93 (.ZN (n_37_93), .A (n_36_92), .B (n_34_95), .C1 (n_33_94), .C2 (n_27_95) );
AOI211_X1 g_39_92 (.ZN (n_39_92), .A (n_35_94), .B (n_32_94), .C1 (n_35_93), .C2 (n_29_96) );
AOI211_X1 g_41_91 (.ZN (n_41_91), .A (n_37_93), .B (n_34_93), .C1 (n_34_95), .C2 (n_31_95) );
AOI211_X1 g_43_90 (.ZN (n_43_90), .A (n_39_92), .B (n_36_92), .C1 (n_32_94), .C2 (n_33_94) );
AOI211_X1 g_45_89 (.ZN (n_45_89), .A (n_41_91), .B (n_35_94), .C1 (n_34_93), .C2 (n_35_93) );
AOI211_X1 g_44_91 (.ZN (n_44_91), .A (n_43_90), .B (n_37_93), .C1 (n_36_92), .C2 (n_34_95) );
AOI211_X1 g_42_90 (.ZN (n_42_90), .A (n_45_89), .B (n_39_92), .C1 (n_35_94), .C2 (n_32_94) );
AOI211_X1 g_44_89 (.ZN (n_44_89), .A (n_44_91), .B (n_41_91), .C1 (n_37_93), .C2 (n_34_93) );
AOI211_X1 g_46_88 (.ZN (n_46_88), .A (n_42_90), .B (n_43_90), .C1 (n_39_92), .C2 (n_36_92) );
AOI211_X1 g_48_87 (.ZN (n_48_87), .A (n_44_89), .B (n_45_89), .C1 (n_41_91), .C2 (n_35_94) );
AOI211_X1 g_50_86 (.ZN (n_50_86), .A (n_46_88), .B (n_44_91), .C1 (n_43_90), .C2 (n_37_93) );
AOI211_X1 g_52_85 (.ZN (n_52_85), .A (n_48_87), .B (n_42_90), .C1 (n_45_89), .C2 (n_39_92) );
AOI211_X1 g_54_84 (.ZN (n_54_84), .A (n_50_86), .B (n_44_89), .C1 (n_44_91), .C2 (n_41_91) );
AOI211_X1 g_56_85 (.ZN (n_56_85), .A (n_52_85), .B (n_46_88), .C1 (n_42_90), .C2 (n_43_90) );
AOI211_X1 g_54_86 (.ZN (n_54_86), .A (n_54_84), .B (n_48_87), .C1 (n_44_89), .C2 (n_45_89) );
AOI211_X1 g_52_87 (.ZN (n_52_87), .A (n_56_85), .B (n_50_86), .C1 (n_46_88), .C2 (n_44_91) );
AOI211_X1 g_50_88 (.ZN (n_50_88), .A (n_54_86), .B (n_52_85), .C1 (n_48_87), .C2 (n_42_90) );
AOI211_X1 g_48_89 (.ZN (n_48_89), .A (n_52_87), .B (n_54_84), .C1 (n_50_86), .C2 (n_44_89) );
AOI211_X1 g_46_90 (.ZN (n_46_90), .A (n_50_88), .B (n_56_85), .C1 (n_52_85), .C2 (n_46_88) );
AOI211_X1 g_45_92 (.ZN (n_45_92), .A (n_48_89), .B (n_54_86), .C1 (n_54_84), .C2 (n_48_87) );
AOI211_X1 g_43_91 (.ZN (n_43_91), .A (n_46_90), .B (n_52_87), .C1 (n_56_85), .C2 (n_50_86) );
AOI211_X1 g_45_90 (.ZN (n_45_90), .A (n_45_92), .B (n_50_88), .C1 (n_54_86), .C2 (n_52_85) );
AOI211_X1 g_47_89 (.ZN (n_47_89), .A (n_43_91), .B (n_48_89), .C1 (n_52_87), .C2 (n_54_84) );
AOI211_X1 g_49_88 (.ZN (n_49_88), .A (n_45_90), .B (n_46_90), .C1 (n_50_88), .C2 (n_56_85) );
AOI211_X1 g_51_87 (.ZN (n_51_87), .A (n_47_89), .B (n_45_92), .C1 (n_48_89), .C2 (n_54_86) );
AOI211_X1 g_53_86 (.ZN (n_53_86), .A (n_49_88), .B (n_43_91), .C1 (n_46_90), .C2 (n_52_87) );
AOI211_X1 g_55_85 (.ZN (n_55_85), .A (n_51_87), .B (n_45_90), .C1 (n_45_92), .C2 (n_50_88) );
AOI211_X1 g_57_84 (.ZN (n_57_84), .A (n_53_86), .B (n_47_89), .C1 (n_43_91), .C2 (n_48_89) );
AOI211_X1 g_59_83 (.ZN (n_59_83), .A (n_55_85), .B (n_49_88), .C1 (n_45_90), .C2 (n_46_90) );
AOI211_X1 g_61_82 (.ZN (n_61_82), .A (n_57_84), .B (n_51_87), .C1 (n_47_89), .C2 (n_45_92) );
AOI211_X1 g_60_84 (.ZN (n_60_84), .A (n_59_83), .B (n_53_86), .C1 (n_49_88), .C2 (n_43_91) );
AOI211_X1 g_62_83 (.ZN (n_62_83), .A (n_61_82), .B (n_55_85), .C1 (n_51_87), .C2 (n_45_90) );
AOI211_X1 g_64_82 (.ZN (n_64_82), .A (n_60_84), .B (n_57_84), .C1 (n_53_86), .C2 (n_47_89) );
AOI211_X1 g_66_81 (.ZN (n_66_81), .A (n_62_83), .B (n_59_83), .C1 (n_55_85), .C2 (n_49_88) );
AOI211_X1 g_68_80 (.ZN (n_68_80), .A (n_64_82), .B (n_61_82), .C1 (n_57_84), .C2 (n_51_87) );
AOI211_X1 g_70_79 (.ZN (n_70_79), .A (n_66_81), .B (n_60_84), .C1 (n_59_83), .C2 (n_53_86) );
AOI211_X1 g_72_78 (.ZN (n_72_78), .A (n_68_80), .B (n_62_83), .C1 (n_61_82), .C2 (n_55_85) );
AOI211_X1 g_74_77 (.ZN (n_74_77), .A (n_70_79), .B (n_64_82), .C1 (n_60_84), .C2 (n_57_84) );
AOI211_X1 g_76_76 (.ZN (n_76_76), .A (n_72_78), .B (n_66_81), .C1 (n_62_83), .C2 (n_59_83) );
AOI211_X1 g_78_75 (.ZN (n_78_75), .A (n_74_77), .B (n_68_80), .C1 (n_64_82), .C2 (n_61_82) );
AOI211_X1 g_80_74 (.ZN (n_80_74), .A (n_76_76), .B (n_70_79), .C1 (n_66_81), .C2 (n_60_84) );
AOI211_X1 g_82_73 (.ZN (n_82_73), .A (n_78_75), .B (n_72_78), .C1 (n_68_80), .C2 (n_62_83) );
AOI211_X1 g_84_72 (.ZN (n_84_72), .A (n_80_74), .B (n_74_77), .C1 (n_70_79), .C2 (n_64_82) );
AOI211_X1 g_86_71 (.ZN (n_86_71), .A (n_82_73), .B (n_76_76), .C1 (n_72_78), .C2 (n_66_81) );
AOI211_X1 g_88_70 (.ZN (n_88_70), .A (n_84_72), .B (n_78_75), .C1 (n_74_77), .C2 (n_68_80) );
AOI211_X1 g_90_69 (.ZN (n_90_69), .A (n_86_71), .B (n_80_74), .C1 (n_76_76), .C2 (n_70_79) );
AOI211_X1 g_92_68 (.ZN (n_92_68), .A (n_88_70), .B (n_82_73), .C1 (n_78_75), .C2 (n_72_78) );
AOI211_X1 g_94_67 (.ZN (n_94_67), .A (n_90_69), .B (n_84_72), .C1 (n_80_74), .C2 (n_74_77) );
AOI211_X1 g_93_69 (.ZN (n_93_69), .A (n_92_68), .B (n_86_71), .C1 (n_82_73), .C2 (n_76_76) );
AOI211_X1 g_95_68 (.ZN (n_95_68), .A (n_94_67), .B (n_88_70), .C1 (n_84_72), .C2 (n_78_75) );
AOI211_X1 g_94_70 (.ZN (n_94_70), .A (n_93_69), .B (n_90_69), .C1 (n_86_71), .C2 (n_80_74) );
AOI211_X1 g_96_69 (.ZN (n_96_69), .A (n_95_68), .B (n_92_68), .C1 (n_88_70), .C2 (n_82_73) );
AOI211_X1 g_94_68 (.ZN (n_94_68), .A (n_94_70), .B (n_94_67), .C1 (n_90_69), .C2 (n_84_72) );
AOI211_X1 g_96_67 (.ZN (n_96_67), .A (n_96_69), .B (n_93_69), .C1 (n_92_68), .C2 (n_86_71) );
AOI211_X1 g_98_68 (.ZN (n_98_68), .A (n_94_68), .B (n_95_68), .C1 (n_94_67), .C2 (n_88_70) );
AOI211_X1 g_97_70 (.ZN (n_97_70), .A (n_96_67), .B (n_94_70), .C1 (n_93_69), .C2 (n_90_69) );
AOI211_X1 g_95_69 (.ZN (n_95_69), .A (n_98_68), .B (n_96_69), .C1 (n_95_68), .C2 (n_92_68) );
AOI211_X1 g_97_68 (.ZN (n_97_68), .A (n_97_70), .B (n_94_68), .C1 (n_94_70), .C2 (n_94_67) );
AOI211_X1 g_99_67 (.ZN (n_99_67), .A (n_95_69), .B (n_96_67), .C1 (n_96_69), .C2 (n_93_69) );
AOI211_X1 g_101_66 (.ZN (n_101_66), .A (n_97_68), .B (n_98_68), .C1 (n_94_68), .C2 (n_95_68) );
AOI211_X1 g_103_65 (.ZN (n_103_65), .A (n_99_67), .B (n_97_70), .C1 (n_96_67), .C2 (n_94_70) );
AOI211_X1 g_105_64 (.ZN (n_105_64), .A (n_101_66), .B (n_95_69), .C1 (n_98_68), .C2 (n_96_69) );
AOI211_X1 g_107_63 (.ZN (n_107_63), .A (n_103_65), .B (n_97_68), .C1 (n_97_70), .C2 (n_94_68) );
AOI211_X1 g_109_62 (.ZN (n_109_62), .A (n_105_64), .B (n_99_67), .C1 (n_95_69), .C2 (n_96_67) );
AOI211_X1 g_108_64 (.ZN (n_108_64), .A (n_107_63), .B (n_101_66), .C1 (n_97_68), .C2 (n_98_68) );
AOI211_X1 g_107_62 (.ZN (n_107_62), .A (n_109_62), .B (n_103_65), .C1 (n_99_67), .C2 (n_97_70) );
AOI211_X1 g_105_63 (.ZN (n_105_63), .A (n_108_64), .B (n_105_64), .C1 (n_101_66), .C2 (n_95_69) );
AOI211_X1 g_106_65 (.ZN (n_106_65), .A (n_107_62), .B (n_107_63), .C1 (n_103_65), .C2 (n_97_68) );
AOI211_X1 g_104_66 (.ZN (n_104_66), .A (n_105_63), .B (n_109_62), .C1 (n_105_64), .C2 (n_99_67) );
AOI211_X1 g_102_67 (.ZN (n_102_67), .A (n_106_65), .B (n_108_64), .C1 (n_107_63), .C2 (n_101_66) );
AOI211_X1 g_100_68 (.ZN (n_100_68), .A (n_104_66), .B (n_107_62), .C1 (n_109_62), .C2 (n_103_65) );
AOI211_X1 g_98_69 (.ZN (n_98_69), .A (n_102_67), .B (n_105_63), .C1 (n_108_64), .C2 (n_105_64) );
AOI211_X1 g_96_70 (.ZN (n_96_70), .A (n_100_68), .B (n_106_65), .C1 (n_107_62), .C2 (n_107_63) );
AOI211_X1 g_94_69 (.ZN (n_94_69), .A (n_98_69), .B (n_104_66), .C1 (n_105_63), .C2 (n_109_62) );
AOI211_X1 g_92_70 (.ZN (n_92_70), .A (n_96_70), .B (n_102_67), .C1 (n_106_65), .C2 (n_108_64) );
AOI211_X1 g_94_71 (.ZN (n_94_71), .A (n_94_69), .B (n_100_68), .C1 (n_104_66), .C2 (n_107_62) );
AOI211_X1 g_96_72 (.ZN (n_96_72), .A (n_92_70), .B (n_98_69), .C1 (n_102_67), .C2 (n_105_63) );
AOI211_X1 g_95_70 (.ZN (n_95_70), .A (n_94_71), .B (n_96_70), .C1 (n_100_68), .C2 (n_106_65) );
AOI211_X1 g_97_69 (.ZN (n_97_69), .A (n_96_72), .B (n_94_69), .C1 (n_98_69), .C2 (n_104_66) );
AOI211_X1 g_99_68 (.ZN (n_99_68), .A (n_95_70), .B (n_92_70), .C1 (n_96_70), .C2 (n_102_67) );
AOI211_X1 g_101_67 (.ZN (n_101_67), .A (n_97_69), .B (n_94_71), .C1 (n_94_69), .C2 (n_100_68) );
AOI211_X1 g_103_66 (.ZN (n_103_66), .A (n_99_68), .B (n_96_72), .C1 (n_92_70), .C2 (n_98_69) );
AOI211_X1 g_105_65 (.ZN (n_105_65), .A (n_101_67), .B (n_95_70), .C1 (n_94_71), .C2 (n_96_70) );
AOI211_X1 g_107_64 (.ZN (n_107_64), .A (n_103_66), .B (n_97_69), .C1 (n_96_72), .C2 (n_94_69) );
AOI211_X1 g_109_63 (.ZN (n_109_63), .A (n_105_65), .B (n_99_68), .C1 (n_95_70), .C2 (n_92_70) );
AOI211_X1 g_111_62 (.ZN (n_111_62), .A (n_107_64), .B (n_101_67), .C1 (n_97_69), .C2 (n_94_71) );
AOI211_X1 g_113_61 (.ZN (n_113_61), .A (n_109_63), .B (n_103_66), .C1 (n_99_68), .C2 (n_96_72) );
AOI211_X1 g_112_63 (.ZN (n_112_63), .A (n_111_62), .B (n_105_65), .C1 (n_101_67), .C2 (n_95_70) );
AOI211_X1 g_114_62 (.ZN (n_114_62), .A (n_113_61), .B (n_107_64), .C1 (n_103_66), .C2 (n_97_69) );
AOI211_X1 g_116_61 (.ZN (n_116_61), .A (n_112_63), .B (n_109_63), .C1 (n_105_65), .C2 (n_99_68) );
AOI211_X1 g_118_60 (.ZN (n_118_60), .A (n_114_62), .B (n_111_62), .C1 (n_107_64), .C2 (n_101_67) );
AOI211_X1 g_120_59 (.ZN (n_120_59), .A (n_116_61), .B (n_113_61), .C1 (n_109_63), .C2 (n_103_66) );
AOI211_X1 g_122_58 (.ZN (n_122_58), .A (n_118_60), .B (n_112_63), .C1 (n_111_62), .C2 (n_105_65) );
AOI211_X1 g_124_57 (.ZN (n_124_57), .A (n_120_59), .B (n_114_62), .C1 (n_113_61), .C2 (n_107_64) );
AOI211_X1 g_126_56 (.ZN (n_126_56), .A (n_122_58), .B (n_116_61), .C1 (n_112_63), .C2 (n_109_63) );
AOI211_X1 g_128_55 (.ZN (n_128_55), .A (n_124_57), .B (n_118_60), .C1 (n_114_62), .C2 (n_111_62) );
AOI211_X1 g_130_54 (.ZN (n_130_54), .A (n_126_56), .B (n_120_59), .C1 (n_116_61), .C2 (n_113_61) );
AOI211_X1 g_132_53 (.ZN (n_132_53), .A (n_128_55), .B (n_122_58), .C1 (n_118_60), .C2 (n_112_63) );
AOI211_X1 g_134_52 (.ZN (n_134_52), .A (n_130_54), .B (n_124_57), .C1 (n_120_59), .C2 (n_114_62) );
AOI211_X1 g_136_51 (.ZN (n_136_51), .A (n_132_53), .B (n_126_56), .C1 (n_122_58), .C2 (n_116_61) );
AOI211_X1 g_138_50 (.ZN (n_138_50), .A (n_134_52), .B (n_128_55), .C1 (n_124_57), .C2 (n_118_60) );
AOI211_X1 g_140_51 (.ZN (n_140_51), .A (n_136_51), .B (n_130_54), .C1 (n_126_56), .C2 (n_120_59) );
AOI211_X1 g_138_52 (.ZN (n_138_52), .A (n_138_50), .B (n_132_53), .C1 (n_128_55), .C2 (n_122_58) );
AOI211_X1 g_139_50 (.ZN (n_139_50), .A (n_140_51), .B (n_134_52), .C1 (n_130_54), .C2 (n_124_57) );
AOI211_X1 g_140_48 (.ZN (n_140_48), .A (n_138_52), .B (n_136_51), .C1 (n_132_53), .C2 (n_126_56) );
AOI211_X1 g_138_49 (.ZN (n_138_49), .A (n_139_50), .B (n_138_50), .C1 (n_134_52), .C2 (n_128_55) );
AOI211_X1 g_136_50 (.ZN (n_136_50), .A (n_140_48), .B (n_140_51), .C1 (n_136_51), .C2 (n_130_54) );
AOI211_X1 g_134_51 (.ZN (n_134_51), .A (n_138_49), .B (n_138_52), .C1 (n_138_50), .C2 (n_132_53) );
AOI211_X1 g_132_52 (.ZN (n_132_52), .A (n_136_50), .B (n_139_50), .C1 (n_140_51), .C2 (n_134_52) );
AOI211_X1 g_130_53 (.ZN (n_130_53), .A (n_134_51), .B (n_140_48), .C1 (n_138_52), .C2 (n_136_51) );
AOI211_X1 g_128_54 (.ZN (n_128_54), .A (n_132_52), .B (n_138_49), .C1 (n_139_50), .C2 (n_138_50) );
AOI211_X1 g_126_55 (.ZN (n_126_55), .A (n_130_53), .B (n_136_50), .C1 (n_140_48), .C2 (n_140_51) );
AOI211_X1 g_124_56 (.ZN (n_124_56), .A (n_128_54), .B (n_134_51), .C1 (n_138_49), .C2 (n_138_52) );
AOI211_X1 g_122_57 (.ZN (n_122_57), .A (n_126_55), .B (n_132_52), .C1 (n_136_50), .C2 (n_139_50) );
AOI211_X1 g_120_58 (.ZN (n_120_58), .A (n_124_56), .B (n_130_53), .C1 (n_134_51), .C2 (n_140_48) );
AOI211_X1 g_118_59 (.ZN (n_118_59), .A (n_122_57), .B (n_128_54), .C1 (n_132_52), .C2 (n_138_49) );
AOI211_X1 g_116_60 (.ZN (n_116_60), .A (n_120_58), .B (n_126_55), .C1 (n_130_53), .C2 (n_136_50) );
AOI211_X1 g_114_61 (.ZN (n_114_61), .A (n_118_59), .B (n_124_56), .C1 (n_128_54), .C2 (n_134_51) );
AOI211_X1 g_112_62 (.ZN (n_112_62), .A (n_116_60), .B (n_122_57), .C1 (n_126_55), .C2 (n_132_52) );
AOI211_X1 g_111_64 (.ZN (n_111_64), .A (n_114_61), .B (n_120_58), .C1 (n_124_56), .C2 (n_130_53) );
AOI211_X1 g_113_63 (.ZN (n_113_63), .A (n_112_62), .B (n_118_59), .C1 (n_122_57), .C2 (n_128_54) );
AOI211_X1 g_115_62 (.ZN (n_115_62), .A (n_111_64), .B (n_116_60), .C1 (n_120_58), .C2 (n_126_55) );
AOI211_X1 g_117_61 (.ZN (n_117_61), .A (n_113_63), .B (n_114_61), .C1 (n_118_59), .C2 (n_124_56) );
AOI211_X1 g_119_60 (.ZN (n_119_60), .A (n_115_62), .B (n_112_62), .C1 (n_116_60), .C2 (n_122_57) );
AOI211_X1 g_121_59 (.ZN (n_121_59), .A (n_117_61), .B (n_111_64), .C1 (n_114_61), .C2 (n_120_58) );
AOI211_X1 g_123_58 (.ZN (n_123_58), .A (n_119_60), .B (n_113_63), .C1 (n_112_62), .C2 (n_118_59) );
AOI211_X1 g_125_57 (.ZN (n_125_57), .A (n_121_59), .B (n_115_62), .C1 (n_111_64), .C2 (n_116_60) );
AOI211_X1 g_127_56 (.ZN (n_127_56), .A (n_123_58), .B (n_117_61), .C1 (n_113_63), .C2 (n_114_61) );
AOI211_X1 g_129_55 (.ZN (n_129_55), .A (n_125_57), .B (n_119_60), .C1 (n_115_62), .C2 (n_112_62) );
AOI211_X1 g_131_54 (.ZN (n_131_54), .A (n_127_56), .B (n_121_59), .C1 (n_117_61), .C2 (n_111_64) );
AOI211_X1 g_133_53 (.ZN (n_133_53), .A (n_129_55), .B (n_123_58), .C1 (n_119_60), .C2 (n_113_63) );
AOI211_X1 g_135_52 (.ZN (n_135_52), .A (n_131_54), .B (n_125_57), .C1 (n_121_59), .C2 (n_115_62) );
AOI211_X1 g_137_51 (.ZN (n_137_51), .A (n_133_53), .B (n_127_56), .C1 (n_123_58), .C2 (n_117_61) );
AOI211_X1 g_136_53 (.ZN (n_136_53), .A (n_135_52), .B (n_129_55), .C1 (n_125_57), .C2 (n_119_60) );
AOI211_X1 g_134_54 (.ZN (n_134_54), .A (n_137_51), .B (n_131_54), .C1 (n_127_56), .C2 (n_121_59) );
AOI211_X1 g_132_55 (.ZN (n_132_55), .A (n_136_53), .B (n_133_53), .C1 (n_129_55), .C2 (n_123_58) );
AOI211_X1 g_131_53 (.ZN (n_131_53), .A (n_134_54), .B (n_135_52), .C1 (n_131_54), .C2 (n_125_57) );
AOI211_X1 g_129_54 (.ZN (n_129_54), .A (n_132_55), .B (n_137_51), .C1 (n_133_53), .C2 (n_127_56) );
AOI211_X1 g_127_55 (.ZN (n_127_55), .A (n_131_53), .B (n_136_53), .C1 (n_135_52), .C2 (n_129_55) );
AOI211_X1 g_125_56 (.ZN (n_125_56), .A (n_129_54), .B (n_134_54), .C1 (n_137_51), .C2 (n_131_54) );
AOI211_X1 g_123_57 (.ZN (n_123_57), .A (n_127_55), .B (n_132_55), .C1 (n_136_53), .C2 (n_133_53) );
AOI211_X1 g_121_58 (.ZN (n_121_58), .A (n_125_56), .B (n_131_53), .C1 (n_134_54), .C2 (n_135_52) );
AOI211_X1 g_119_59 (.ZN (n_119_59), .A (n_123_57), .B (n_129_54), .C1 (n_132_55), .C2 (n_137_51) );
AOI211_X1 g_117_60 (.ZN (n_117_60), .A (n_121_58), .B (n_127_55), .C1 (n_131_53), .C2 (n_136_53) );
AOI211_X1 g_115_61 (.ZN (n_115_61), .A (n_119_59), .B (n_125_56), .C1 (n_129_54), .C2 (n_134_54) );
AOI211_X1 g_113_62 (.ZN (n_113_62), .A (n_117_60), .B (n_123_57), .C1 (n_127_55), .C2 (n_132_55) );
AOI211_X1 g_111_63 (.ZN (n_111_63), .A (n_115_61), .B (n_121_58), .C1 (n_125_56), .C2 (n_131_53) );
AOI211_X1 g_109_64 (.ZN (n_109_64), .A (n_113_62), .B (n_119_59), .C1 (n_123_57), .C2 (n_129_54) );
AOI211_X1 g_107_65 (.ZN (n_107_65), .A (n_111_63), .B (n_117_60), .C1 (n_121_58), .C2 (n_127_55) );
AOI211_X1 g_108_63 (.ZN (n_108_63), .A (n_109_64), .B (n_115_61), .C1 (n_119_59), .C2 (n_125_56) );
AOI211_X1 g_106_64 (.ZN (n_106_64), .A (n_107_65), .B (n_113_62), .C1 (n_117_60), .C2 (n_123_57) );
AOI211_X1 g_104_65 (.ZN (n_104_65), .A (n_108_63), .B (n_111_63), .C1 (n_115_61), .C2 (n_121_58) );
AOI211_X1 g_102_66 (.ZN (n_102_66), .A (n_106_64), .B (n_109_64), .C1 (n_113_62), .C2 (n_119_59) );
AOI211_X1 g_101_68 (.ZN (n_101_68), .A (n_104_65), .B (n_107_65), .C1 (n_111_63), .C2 (n_117_60) );
AOI211_X1 g_99_69 (.ZN (n_99_69), .A (n_102_66), .B (n_108_63), .C1 (n_109_64), .C2 (n_115_61) );
AOI211_X1 g_98_71 (.ZN (n_98_71), .A (n_101_68), .B (n_106_64), .C1 (n_107_65), .C2 (n_113_62) );
AOI211_X1 g_100_70 (.ZN (n_100_70), .A (n_99_69), .B (n_104_65), .C1 (n_108_63), .C2 (n_111_63) );
AOI211_X1 g_102_69 (.ZN (n_102_69), .A (n_98_71), .B (n_102_66), .C1 (n_106_64), .C2 (n_109_64) );
AOI211_X1 g_103_67 (.ZN (n_103_67), .A (n_100_70), .B (n_101_68), .C1 (n_104_65), .C2 (n_107_65) );
AOI211_X1 g_105_66 (.ZN (n_105_66), .A (n_102_69), .B (n_99_69), .C1 (n_102_66), .C2 (n_108_63) );
AOI211_X1 g_104_68 (.ZN (n_104_68), .A (n_103_67), .B (n_98_71), .C1 (n_101_68), .C2 (n_106_64) );
AOI211_X1 g_106_67 (.ZN (n_106_67), .A (n_105_66), .B (n_100_70), .C1 (n_99_69), .C2 (n_104_65) );
AOI211_X1 g_108_66 (.ZN (n_108_66), .A (n_104_68), .B (n_102_69), .C1 (n_98_71), .C2 (n_102_66) );
AOI211_X1 g_110_65 (.ZN (n_110_65), .A (n_106_67), .B (n_103_67), .C1 (n_100_70), .C2 (n_101_68) );
AOI211_X1 g_112_64 (.ZN (n_112_64), .A (n_108_66), .B (n_105_66), .C1 (n_102_69), .C2 (n_99_69) );
AOI211_X1 g_114_63 (.ZN (n_114_63), .A (n_110_65), .B (n_104_68), .C1 (n_103_67), .C2 (n_98_71) );
AOI211_X1 g_116_62 (.ZN (n_116_62), .A (n_112_64), .B (n_106_67), .C1 (n_105_66), .C2 (n_100_70) );
AOI211_X1 g_118_61 (.ZN (n_118_61), .A (n_114_63), .B (n_108_66), .C1 (n_104_68), .C2 (n_102_69) );
AOI211_X1 g_120_60 (.ZN (n_120_60), .A (n_116_62), .B (n_110_65), .C1 (n_106_67), .C2 (n_103_67) );
AOI211_X1 g_122_59 (.ZN (n_122_59), .A (n_118_61), .B (n_112_64), .C1 (n_108_66), .C2 (n_105_66) );
AOI211_X1 g_124_58 (.ZN (n_124_58), .A (n_120_60), .B (n_114_63), .C1 (n_110_65), .C2 (n_104_68) );
AOI211_X1 g_126_57 (.ZN (n_126_57), .A (n_122_59), .B (n_116_62), .C1 (n_112_64), .C2 (n_106_67) );
AOI211_X1 g_128_56 (.ZN (n_128_56), .A (n_124_58), .B (n_118_61), .C1 (n_114_63), .C2 (n_108_66) );
AOI211_X1 g_130_55 (.ZN (n_130_55), .A (n_126_57), .B (n_120_60), .C1 (n_116_62), .C2 (n_110_65) );
AOI211_X1 g_132_54 (.ZN (n_132_54), .A (n_128_56), .B (n_122_59), .C1 (n_118_61), .C2 (n_112_64) );
AOI211_X1 g_134_53 (.ZN (n_134_53), .A (n_130_55), .B (n_124_58), .C1 (n_120_60), .C2 (n_114_63) );
AOI211_X1 g_136_52 (.ZN (n_136_52), .A (n_132_54), .B (n_126_57), .C1 (n_122_59), .C2 (n_116_62) );
AOI211_X1 g_138_51 (.ZN (n_138_51), .A (n_134_53), .B (n_128_56), .C1 (n_124_58), .C2 (n_118_61) );
AOI211_X1 g_140_50 (.ZN (n_140_50), .A (n_136_52), .B (n_130_55), .C1 (n_126_57), .C2 (n_120_60) );
AOI211_X1 g_142_49 (.ZN (n_142_49), .A (n_138_51), .B (n_132_54), .C1 (n_128_56), .C2 (n_122_59) );
AOI211_X1 g_141_51 (.ZN (n_141_51), .A (n_140_50), .B (n_134_53), .C1 (n_130_55), .C2 (n_124_58) );
AOI211_X1 g_139_52 (.ZN (n_139_52), .A (n_142_49), .B (n_136_52), .C1 (n_132_54), .C2 (n_126_57) );
AOI211_X1 g_137_53 (.ZN (n_137_53), .A (n_141_51), .B (n_138_51), .C1 (n_134_53), .C2 (n_128_56) );
AOI211_X1 g_135_54 (.ZN (n_135_54), .A (n_139_52), .B (n_140_50), .C1 (n_136_52), .C2 (n_130_55) );
AOI211_X1 g_133_55 (.ZN (n_133_55), .A (n_137_53), .B (n_142_49), .C1 (n_138_51), .C2 (n_132_54) );
AOI211_X1 g_131_56 (.ZN (n_131_56), .A (n_135_54), .B (n_141_51), .C1 (n_140_50), .C2 (n_134_53) );
AOI211_X1 g_129_57 (.ZN (n_129_57), .A (n_133_55), .B (n_139_52), .C1 (n_142_49), .C2 (n_136_52) );
AOI211_X1 g_127_58 (.ZN (n_127_58), .A (n_131_56), .B (n_137_53), .C1 (n_141_51), .C2 (n_138_51) );
AOI211_X1 g_125_59 (.ZN (n_125_59), .A (n_129_57), .B (n_135_54), .C1 (n_139_52), .C2 (n_140_50) );
AOI211_X1 g_123_60 (.ZN (n_123_60), .A (n_127_58), .B (n_133_55), .C1 (n_137_53), .C2 (n_142_49) );
AOI211_X1 g_121_61 (.ZN (n_121_61), .A (n_125_59), .B (n_131_56), .C1 (n_135_54), .C2 (n_141_51) );
AOI211_X1 g_119_62 (.ZN (n_119_62), .A (n_123_60), .B (n_129_57), .C1 (n_133_55), .C2 (n_139_52) );
AOI211_X1 g_117_63 (.ZN (n_117_63), .A (n_121_61), .B (n_127_58), .C1 (n_131_56), .C2 (n_137_53) );
AOI211_X1 g_115_64 (.ZN (n_115_64), .A (n_119_62), .B (n_125_59), .C1 (n_129_57), .C2 (n_135_54) );
AOI211_X1 g_113_65 (.ZN (n_113_65), .A (n_117_63), .B (n_123_60), .C1 (n_127_58), .C2 (n_133_55) );
AOI211_X1 g_111_66 (.ZN (n_111_66), .A (n_115_64), .B (n_121_61), .C1 (n_125_59), .C2 (n_131_56) );
AOI211_X1 g_110_64 (.ZN (n_110_64), .A (n_113_65), .B (n_119_62), .C1 (n_123_60), .C2 (n_129_57) );
AOI211_X1 g_108_65 (.ZN (n_108_65), .A (n_111_66), .B (n_117_63), .C1 (n_121_61), .C2 (n_127_58) );
AOI211_X1 g_106_66 (.ZN (n_106_66), .A (n_110_64), .B (n_115_64), .C1 (n_119_62), .C2 (n_125_59) );
AOI211_X1 g_104_67 (.ZN (n_104_67), .A (n_108_65), .B (n_113_65), .C1 (n_117_63), .C2 (n_123_60) );
AOI211_X1 g_102_68 (.ZN (n_102_68), .A (n_106_66), .B (n_111_66), .C1 (n_115_64), .C2 (n_121_61) );
AOI211_X1 g_100_69 (.ZN (n_100_69), .A (n_104_67), .B (n_110_64), .C1 (n_113_65), .C2 (n_119_62) );
AOI211_X1 g_98_70 (.ZN (n_98_70), .A (n_102_68), .B (n_108_65), .C1 (n_111_66), .C2 (n_117_63) );
AOI211_X1 g_96_71 (.ZN (n_96_71), .A (n_100_69), .B (n_106_66), .C1 (n_110_64), .C2 (n_115_64) );
AOI211_X1 g_94_72 (.ZN (n_94_72), .A (n_98_70), .B (n_104_67), .C1 (n_108_65), .C2 (n_113_65) );
AOI211_X1 g_93_70 (.ZN (n_93_70), .A (n_96_71), .B (n_102_68), .C1 (n_106_66), .C2 (n_111_66) );
AOI211_X1 g_91_69 (.ZN (n_91_69), .A (n_94_72), .B (n_100_69), .C1 (n_104_67), .C2 (n_110_64) );
AOI211_X1 g_92_71 (.ZN (n_92_71), .A (n_93_70), .B (n_98_70), .C1 (n_102_68), .C2 (n_108_65) );
AOI211_X1 g_90_72 (.ZN (n_90_72), .A (n_91_69), .B (n_96_71), .C1 (n_100_69), .C2 (n_106_66) );
AOI211_X1 g_91_70 (.ZN (n_91_70), .A (n_92_71), .B (n_94_72), .C1 (n_98_70), .C2 (n_104_67) );
AOI211_X1 g_89_71 (.ZN (n_89_71), .A (n_90_72), .B (n_93_70), .C1 (n_96_71), .C2 (n_102_68) );
AOI211_X1 g_87_72 (.ZN (n_87_72), .A (n_91_70), .B (n_91_69), .C1 (n_94_72), .C2 (n_100_69) );
AOI211_X1 g_85_73 (.ZN (n_85_73), .A (n_89_71), .B (n_92_71), .C1 (n_93_70), .C2 (n_98_70) );
AOI211_X1 g_84_71 (.ZN (n_84_71), .A (n_87_72), .B (n_90_72), .C1 (n_91_69), .C2 (n_96_71) );
AOI211_X1 g_82_72 (.ZN (n_82_72), .A (n_85_73), .B (n_91_70), .C1 (n_92_71), .C2 (n_94_72) );
AOI211_X1 g_80_73 (.ZN (n_80_73), .A (n_84_71), .B (n_89_71), .C1 (n_90_72), .C2 (n_93_70) );
AOI211_X1 g_78_74 (.ZN (n_78_74), .A (n_82_72), .B (n_87_72), .C1 (n_91_70), .C2 (n_91_69) );
AOI211_X1 g_76_75 (.ZN (n_76_75), .A (n_80_73), .B (n_85_73), .C1 (n_89_71), .C2 (n_92_71) );
AOI211_X1 g_74_76 (.ZN (n_74_76), .A (n_78_74), .B (n_84_71), .C1 (n_87_72), .C2 (n_90_72) );
AOI211_X1 g_72_77 (.ZN (n_72_77), .A (n_76_75), .B (n_82_72), .C1 (n_85_73), .C2 (n_91_70) );
AOI211_X1 g_70_78 (.ZN (n_70_78), .A (n_74_76), .B (n_80_73), .C1 (n_84_71), .C2 (n_89_71) );
AOI211_X1 g_68_79 (.ZN (n_68_79), .A (n_72_77), .B (n_78_74), .C1 (n_82_72), .C2 (n_87_72) );
AOI211_X1 g_66_80 (.ZN (n_66_80), .A (n_70_78), .B (n_76_75), .C1 (n_80_73), .C2 (n_85_73) );
AOI211_X1 g_64_81 (.ZN (n_64_81), .A (n_68_79), .B (n_74_76), .C1 (n_78_74), .C2 (n_84_71) );
AOI211_X1 g_62_82 (.ZN (n_62_82), .A (n_66_80), .B (n_72_77), .C1 (n_76_75), .C2 (n_82_72) );
AOI211_X1 g_60_83 (.ZN (n_60_83), .A (n_64_81), .B (n_70_78), .C1 (n_74_76), .C2 (n_80_73) );
AOI211_X1 g_59_85 (.ZN (n_59_85), .A (n_62_82), .B (n_68_79), .C1 (n_72_77), .C2 (n_78_74) );
AOI211_X1 g_61_84 (.ZN (n_61_84), .A (n_60_83), .B (n_66_80), .C1 (n_70_78), .C2 (n_76_75) );
AOI211_X1 g_63_83 (.ZN (n_63_83), .A (n_59_85), .B (n_64_81), .C1 (n_68_79), .C2 (n_74_76) );
AOI211_X1 g_65_82 (.ZN (n_65_82), .A (n_61_84), .B (n_62_82), .C1 (n_66_80), .C2 (n_72_77) );
AOI211_X1 g_67_81 (.ZN (n_67_81), .A (n_63_83), .B (n_60_83), .C1 (n_64_81), .C2 (n_70_78) );
AOI211_X1 g_69_80 (.ZN (n_69_80), .A (n_65_82), .B (n_59_85), .C1 (n_62_82), .C2 (n_68_79) );
AOI211_X1 g_71_79 (.ZN (n_71_79), .A (n_67_81), .B (n_61_84), .C1 (n_60_83), .C2 (n_66_80) );
AOI211_X1 g_73_78 (.ZN (n_73_78), .A (n_69_80), .B (n_63_83), .C1 (n_59_85), .C2 (n_64_81) );
AOI211_X1 g_75_77 (.ZN (n_75_77), .A (n_71_79), .B (n_65_82), .C1 (n_61_84), .C2 (n_62_82) );
AOI211_X1 g_77_76 (.ZN (n_77_76), .A (n_73_78), .B (n_67_81), .C1 (n_63_83), .C2 (n_60_83) );
AOI211_X1 g_79_75 (.ZN (n_79_75), .A (n_75_77), .B (n_69_80), .C1 (n_65_82), .C2 (n_59_85) );
AOI211_X1 g_81_74 (.ZN (n_81_74), .A (n_77_76), .B (n_71_79), .C1 (n_67_81), .C2 (n_61_84) );
AOI211_X1 g_83_73 (.ZN (n_83_73), .A (n_79_75), .B (n_73_78), .C1 (n_69_80), .C2 (n_63_83) );
AOI211_X1 g_85_72 (.ZN (n_85_72), .A (n_81_74), .B (n_75_77), .C1 (n_71_79), .C2 (n_65_82) );
AOI211_X1 g_87_71 (.ZN (n_87_71), .A (n_83_73), .B (n_77_76), .C1 (n_73_78), .C2 (n_67_81) );
AOI211_X1 g_89_70 (.ZN (n_89_70), .A (n_85_72), .B (n_79_75), .C1 (n_75_77), .C2 (n_69_80) );
AOI211_X1 g_91_71 (.ZN (n_91_71), .A (n_87_71), .B (n_81_74), .C1 (n_77_76), .C2 (n_71_79) );
AOI211_X1 g_89_72 (.ZN (n_89_72), .A (n_89_70), .B (n_83_73), .C1 (n_79_75), .C2 (n_73_78) );
AOI211_X1 g_87_73 (.ZN (n_87_73), .A (n_91_71), .B (n_85_72), .C1 (n_81_74), .C2 (n_75_77) );
AOI211_X1 g_85_74 (.ZN (n_85_74), .A (n_89_72), .B (n_87_71), .C1 (n_83_73), .C2 (n_77_76) );
AOI211_X1 g_86_72 (.ZN (n_86_72), .A (n_87_73), .B (n_89_70), .C1 (n_85_72), .C2 (n_79_75) );
AOI211_X1 g_84_73 (.ZN (n_84_73), .A (n_85_74), .B (n_91_71), .C1 (n_87_71), .C2 (n_81_74) );
AOI211_X1 g_82_74 (.ZN (n_82_74), .A (n_86_72), .B (n_89_72), .C1 (n_89_70), .C2 (n_83_73) );
AOI211_X1 g_80_75 (.ZN (n_80_75), .A (n_84_73), .B (n_87_73), .C1 (n_91_71), .C2 (n_85_72) );
AOI211_X1 g_78_76 (.ZN (n_78_76), .A (n_82_74), .B (n_85_74), .C1 (n_89_72), .C2 (n_87_71) );
AOI211_X1 g_76_77 (.ZN (n_76_77), .A (n_80_75), .B (n_86_72), .C1 (n_87_73), .C2 (n_89_70) );
AOI211_X1 g_74_78 (.ZN (n_74_78), .A (n_78_76), .B (n_84_73), .C1 (n_85_74), .C2 (n_91_71) );
AOI211_X1 g_72_79 (.ZN (n_72_79), .A (n_76_77), .B (n_82_74), .C1 (n_86_72), .C2 (n_89_72) );
AOI211_X1 g_70_80 (.ZN (n_70_80), .A (n_74_78), .B (n_80_75), .C1 (n_84_73), .C2 (n_87_73) );
AOI211_X1 g_68_81 (.ZN (n_68_81), .A (n_72_79), .B (n_78_76), .C1 (n_82_74), .C2 (n_85_74) );
AOI211_X1 g_66_82 (.ZN (n_66_82), .A (n_70_80), .B (n_76_77), .C1 (n_80_75), .C2 (n_86_72) );
AOI211_X1 g_64_83 (.ZN (n_64_83), .A (n_68_81), .B (n_74_78), .C1 (n_78_76), .C2 (n_84_73) );
AOI211_X1 g_62_84 (.ZN (n_62_84), .A (n_66_82), .B (n_72_79), .C1 (n_76_77), .C2 (n_82_74) );
AOI211_X1 g_60_85 (.ZN (n_60_85), .A (n_64_83), .B (n_70_80), .C1 (n_74_78), .C2 (n_80_75) );
AOI211_X1 g_61_83 (.ZN (n_61_83), .A (n_62_84), .B (n_68_81), .C1 (n_72_79), .C2 (n_78_76) );
AOI211_X1 g_59_84 (.ZN (n_59_84), .A (n_60_85), .B (n_66_82), .C1 (n_70_80), .C2 (n_76_77) );
AOI211_X1 g_57_85 (.ZN (n_57_85), .A (n_61_83), .B (n_64_83), .C1 (n_68_81), .C2 (n_74_78) );
AOI211_X1 g_55_86 (.ZN (n_55_86), .A (n_59_84), .B (n_62_84), .C1 (n_66_82), .C2 (n_72_79) );
AOI211_X1 g_53_87 (.ZN (n_53_87), .A (n_57_85), .B (n_60_85), .C1 (n_64_83), .C2 (n_70_80) );
AOI211_X1 g_51_88 (.ZN (n_51_88), .A (n_55_86), .B (n_61_83), .C1 (n_62_84), .C2 (n_68_81) );
AOI211_X1 g_49_89 (.ZN (n_49_89), .A (n_53_87), .B (n_59_84), .C1 (n_60_85), .C2 (n_66_82) );
AOI211_X1 g_47_90 (.ZN (n_47_90), .A (n_51_88), .B (n_57_85), .C1 (n_61_83), .C2 (n_64_83) );
AOI211_X1 g_45_91 (.ZN (n_45_91), .A (n_49_89), .B (n_55_86), .C1 (n_59_84), .C2 (n_62_84) );
AOI211_X1 g_43_92 (.ZN (n_43_92), .A (n_47_90), .B (n_53_87), .C1 (n_57_85), .C2 (n_60_85) );
AOI211_X1 g_41_93 (.ZN (n_41_93), .A (n_45_91), .B (n_51_88), .C1 (n_55_86), .C2 (n_61_83) );
AOI211_X1 g_40_91 (.ZN (n_40_91), .A (n_43_92), .B (n_49_89), .C1 (n_53_87), .C2 (n_59_84) );
AOI211_X1 g_38_92 (.ZN (n_38_92), .A (n_41_93), .B (n_47_90), .C1 (n_51_88), .C2 (n_57_85) );
AOI211_X1 g_36_93 (.ZN (n_36_93), .A (n_40_91), .B (n_45_91), .C1 (n_49_89), .C2 (n_55_86) );
AOI211_X1 g_34_94 (.ZN (n_34_94), .A (n_38_92), .B (n_43_92), .C1 (n_47_90), .C2 (n_53_87) );
AOI211_X1 g_32_95 (.ZN (n_32_95), .A (n_36_93), .B (n_41_93), .C1 (n_45_91), .C2 (n_51_88) );
AOI211_X1 g_30_96 (.ZN (n_30_96), .A (n_34_94), .B (n_40_91), .C1 (n_43_92), .C2 (n_49_89) );
AOI211_X1 g_28_97 (.ZN (n_28_97), .A (n_32_95), .B (n_38_92), .C1 (n_41_93), .C2 (n_47_90) );
AOI211_X1 g_26_96 (.ZN (n_26_96), .A (n_30_96), .B (n_36_93), .C1 (n_40_91), .C2 (n_45_91) );
AOI211_X1 g_24_97 (.ZN (n_24_97), .A (n_28_97), .B (n_34_94), .C1 (n_38_92), .C2 (n_43_92) );
AOI211_X1 g_22_98 (.ZN (n_22_98), .A (n_26_96), .B (n_32_95), .C1 (n_36_93), .C2 (n_41_93) );
AOI211_X1 g_21_96 (.ZN (n_21_96), .A (n_24_97), .B (n_30_96), .C1 (n_34_94), .C2 (n_40_91) );
AOI211_X1 g_19_97 (.ZN (n_19_97), .A (n_22_98), .B (n_28_97), .C1 (n_32_95), .C2 (n_38_92) );
AOI211_X1 g_17_98 (.ZN (n_17_98), .A (n_21_96), .B (n_26_96), .C1 (n_30_96), .C2 (n_36_93) );
AOI211_X1 g_15_99 (.ZN (n_15_99), .A (n_19_97), .B (n_24_97), .C1 (n_28_97), .C2 (n_34_94) );
AOI211_X1 g_16_97 (.ZN (n_16_97), .A (n_17_98), .B (n_22_98), .C1 (n_26_96), .C2 (n_32_95) );
AOI211_X1 g_14_98 (.ZN (n_14_98), .A (n_15_99), .B (n_21_96), .C1 (n_24_97), .C2 (n_30_96) );
AOI211_X1 g_12_99 (.ZN (n_12_99), .A (n_16_97), .B (n_19_97), .C1 (n_22_98), .C2 (n_28_97) );
AOI211_X1 g_11_101 (.ZN (n_11_101), .A (n_14_98), .B (n_17_98), .C1 (n_21_96), .C2 (n_26_96) );
AOI211_X1 g_13_100 (.ZN (n_13_100), .A (n_12_99), .B (n_15_99), .C1 (n_19_97), .C2 (n_24_97) );
AOI211_X1 g_12_102 (.ZN (n_12_102), .A (n_11_101), .B (n_16_97), .C1 (n_17_98), .C2 (n_22_98) );
AOI211_X1 g_11_100 (.ZN (n_11_100), .A (n_13_100), .B (n_14_98), .C1 (n_15_99), .C2 (n_21_96) );
AOI211_X1 g_13_99 (.ZN (n_13_99), .A (n_12_102), .B (n_12_99), .C1 (n_16_97), .C2 (n_19_97) );
AOI211_X1 g_15_98 (.ZN (n_15_98), .A (n_11_100), .B (n_11_101), .C1 (n_14_98), .C2 (n_17_98) );
AOI211_X1 g_17_99 (.ZN (n_17_99), .A (n_13_99), .B (n_13_100), .C1 (n_12_99), .C2 (n_15_99) );
AOI211_X1 g_15_100 (.ZN (n_15_100), .A (n_15_98), .B (n_12_102), .C1 (n_11_101), .C2 (n_16_97) );
AOI211_X1 g_13_101 (.ZN (n_13_101), .A (n_17_99), .B (n_11_100), .C1 (n_13_100), .C2 (n_14_98) );
AOI211_X1 g_14_99 (.ZN (n_14_99), .A (n_15_100), .B (n_13_99), .C1 (n_12_102), .C2 (n_12_99) );
AOI211_X1 g_12_100 (.ZN (n_12_100), .A (n_13_101), .B (n_15_98), .C1 (n_11_100), .C2 (n_11_101) );
AOI211_X1 g_11_102 (.ZN (n_11_102), .A (n_14_99), .B (n_17_99), .C1 (n_13_99), .C2 (n_13_100) );
AOI211_X1 g_10_104 (.ZN (n_10_104), .A (n_12_100), .B (n_15_100), .C1 (n_15_98), .C2 (n_12_102) );
AOI211_X1 g_8_103 (.ZN (n_8_103), .A (n_11_102), .B (n_13_101), .C1 (n_17_99), .C2 (n_11_100) );
AOI211_X1 g_10_102 (.ZN (n_10_102), .A (n_10_104), .B (n_14_99), .C1 (n_15_100), .C2 (n_13_99) );
AOI211_X1 g_12_101 (.ZN (n_12_101), .A (n_8_103), .B (n_12_100), .C1 (n_13_101), .C2 (n_15_98) );
AOI211_X1 g_14_100 (.ZN (n_14_100), .A (n_10_102), .B (n_11_102), .C1 (n_14_99), .C2 (n_17_99) );
AOI211_X1 g_16_99 (.ZN (n_16_99), .A (n_12_101), .B (n_10_104), .C1 (n_12_100), .C2 (n_15_100) );
AOI211_X1 g_18_98 (.ZN (n_18_98), .A (n_14_100), .B (n_8_103), .C1 (n_11_102), .C2 (n_13_101) );
AOI211_X1 g_20_99 (.ZN (n_20_99), .A (n_16_99), .B (n_10_102), .C1 (n_10_104), .C2 (n_14_99) );
AOI211_X1 g_18_100 (.ZN (n_18_100), .A (n_18_98), .B (n_12_101), .C1 (n_8_103), .C2 (n_12_100) );
AOI211_X1 g_16_101 (.ZN (n_16_101), .A (n_20_99), .B (n_14_100), .C1 (n_10_102), .C2 (n_11_102) );
AOI211_X1 g_14_102 (.ZN (n_14_102), .A (n_18_100), .B (n_16_99), .C1 (n_12_101), .C2 (n_10_104) );
AOI211_X1 g_12_103 (.ZN (n_12_103), .A (n_16_101), .B (n_18_98), .C1 (n_14_100), .C2 (n_8_103) );
AOI211_X1 g_11_105 (.ZN (n_11_105), .A (n_14_102), .B (n_20_99), .C1 (n_16_99), .C2 (n_10_102) );
AOI211_X1 g_10_103 (.ZN (n_10_103), .A (n_12_103), .B (n_18_100), .C1 (n_18_98), .C2 (n_12_101) );
AOI211_X1 g_8_104 (.ZN (n_8_104), .A (n_11_105), .B (n_16_101), .C1 (n_20_99), .C2 (n_14_100) );
AOI211_X1 g_6_105 (.ZN (n_6_105), .A (n_10_103), .B (n_14_102), .C1 (n_18_100), .C2 (n_16_99) );
AOI211_X1 g_4_106 (.ZN (n_4_106), .A (n_8_104), .B (n_12_103), .C1 (n_16_101), .C2 (n_18_98) );
AOI211_X1 g_3_108 (.ZN (n_3_108), .A (n_6_105), .B (n_11_105), .C1 (n_14_102), .C2 (n_20_99) );
AOI211_X1 g_2_106 (.ZN (n_2_106), .A (n_4_106), .B (n_10_103), .C1 (n_12_103), .C2 (n_18_100) );
AOI211_X1 g_1_108 (.ZN (n_1_108), .A (n_3_108), .B (n_8_104), .C1 (n_11_105), .C2 (n_16_101) );
AOI211_X1 g_3_107 (.ZN (n_3_107), .A (n_2_106), .B (n_6_105), .C1 (n_10_103), .C2 (n_14_102) );
AOI211_X1 g_4_105 (.ZN (n_4_105), .A (n_1_108), .B (n_4_106), .C1 (n_8_104), .C2 (n_12_103) );
AOI211_X1 g_6_104 (.ZN (n_6_104), .A (n_3_107), .B (n_3_108), .C1 (n_6_105), .C2 (n_11_105) );
AOI211_X1 g_5_106 (.ZN (n_5_106), .A (n_4_105), .B (n_2_106), .C1 (n_4_106), .C2 (n_10_103) );
AOI211_X1 g_7_105 (.ZN (n_7_105), .A (n_6_104), .B (n_1_108), .C1 (n_3_108), .C2 (n_8_104) );
AOI211_X1 g_9_104 (.ZN (n_9_104), .A (n_5_106), .B (n_3_107), .C1 (n_2_106), .C2 (n_6_105) );
AOI211_X1 g_11_103 (.ZN (n_11_103), .A (n_7_105), .B (n_4_105), .C1 (n_1_108), .C2 (n_4_106) );
AOI211_X1 g_13_102 (.ZN (n_13_102), .A (n_9_104), .B (n_6_104), .C1 (n_3_107), .C2 (n_3_108) );
AOI211_X1 g_15_101 (.ZN (n_15_101), .A (n_11_103), .B (n_5_106), .C1 (n_4_105), .C2 (n_2_106) );
AOI211_X1 g_17_100 (.ZN (n_17_100), .A (n_13_102), .B (n_7_105), .C1 (n_6_104), .C2 (n_1_108) );
AOI211_X1 g_19_99 (.ZN (n_19_99), .A (n_15_101), .B (n_9_104), .C1 (n_5_106), .C2 (n_3_107) );
AOI211_X1 g_21_98 (.ZN (n_21_98), .A (n_17_100), .B (n_11_103), .C1 (n_7_105), .C2 (n_4_105) );
AOI211_X1 g_23_97 (.ZN (n_23_97), .A (n_19_99), .B (n_13_102), .C1 (n_9_104), .C2 (n_6_104) );
AOI211_X1 g_24_99 (.ZN (n_24_99), .A (n_21_98), .B (n_15_101), .C1 (n_11_103), .C2 (n_5_106) );
AOI211_X1 g_22_100 (.ZN (n_22_100), .A (n_23_97), .B (n_17_100), .C1 (n_13_102), .C2 (n_7_105) );
AOI211_X1 g_20_101 (.ZN (n_20_101), .A (n_24_99), .B (n_19_99), .C1 (n_15_101), .C2 (n_9_104) );
AOI211_X1 g_21_99 (.ZN (n_21_99), .A (n_22_100), .B (n_21_98), .C1 (n_17_100), .C2 (n_11_103) );
AOI211_X1 g_22_97 (.ZN (n_22_97), .A (n_20_101), .B (n_23_97), .C1 (n_19_99), .C2 (n_13_102) );
AOI211_X1 g_20_98 (.ZN (n_20_98), .A (n_21_99), .B (n_24_99), .C1 (n_21_98), .C2 (n_15_101) );
AOI211_X1 g_18_99 (.ZN (n_18_99), .A (n_22_97), .B (n_22_100), .C1 (n_23_97), .C2 (n_17_100) );
AOI211_X1 g_16_100 (.ZN (n_16_100), .A (n_20_98), .B (n_20_101), .C1 (n_24_99), .C2 (n_19_99) );
AOI211_X1 g_14_101 (.ZN (n_14_101), .A (n_18_99), .B (n_21_99), .C1 (n_22_100), .C2 (n_21_98) );
AOI211_X1 g_13_103 (.ZN (n_13_103), .A (n_16_100), .B (n_22_97), .C1 (n_20_101), .C2 (n_23_97) );
AOI211_X1 g_15_102 (.ZN (n_15_102), .A (n_14_101), .B (n_20_98), .C1 (n_21_99), .C2 (n_24_99) );
AOI211_X1 g_17_101 (.ZN (n_17_101), .A (n_13_103), .B (n_18_99), .C1 (n_22_97), .C2 (n_22_100) );
AOI211_X1 g_19_100 (.ZN (n_19_100), .A (n_15_102), .B (n_16_100), .C1 (n_20_98), .C2 (n_20_101) );
AOI211_X1 g_18_102 (.ZN (n_18_102), .A (n_17_101), .B (n_14_101), .C1 (n_18_99), .C2 (n_21_99) );
AOI211_X1 g_16_103 (.ZN (n_16_103), .A (n_19_100), .B (n_13_103), .C1 (n_16_100), .C2 (n_22_97) );
AOI211_X1 g_14_104 (.ZN (n_14_104), .A (n_18_102), .B (n_15_102), .C1 (n_14_101), .C2 (n_20_98) );
AOI211_X1 g_12_105 (.ZN (n_12_105), .A (n_16_103), .B (n_17_101), .C1 (n_13_103), .C2 (n_18_99) );
AOI211_X1 g_10_106 (.ZN (n_10_106), .A (n_14_104), .B (n_19_100), .C1 (n_15_102), .C2 (n_16_100) );
AOI211_X1 g_11_104 (.ZN (n_11_104), .A (n_12_105), .B (n_18_102), .C1 (n_17_101), .C2 (n_14_101) );
AOI211_X1 g_9_105 (.ZN (n_9_105), .A (n_10_106), .B (n_16_103), .C1 (n_19_100), .C2 (n_13_103) );
AOI211_X1 g_7_106 (.ZN (n_7_106), .A (n_11_104), .B (n_14_104), .C1 (n_18_102), .C2 (n_15_102) );
AOI211_X1 g_5_107 (.ZN (n_5_107), .A (n_9_105), .B (n_12_105), .C1 (n_16_103), .C2 (n_17_101) );
AOI211_X1 g_4_109 (.ZN (n_4_109), .A (n_7_106), .B (n_10_106), .C1 (n_14_104), .C2 (n_19_100) );
AOI211_X1 g_2_110 (.ZN (n_2_110), .A (n_5_107), .B (n_11_104), .C1 (n_12_105), .C2 (n_18_102) );
AOI211_X1 g_1_112 (.ZN (n_1_112), .A (n_4_109), .B (n_9_105), .C1 (n_10_106), .C2 (n_16_103) );
AOI211_X1 g_3_111 (.ZN (n_3_111), .A (n_2_110), .B (n_7_106), .C1 (n_11_104), .C2 (n_14_104) );
AOI211_X1 g_5_110 (.ZN (n_5_110), .A (n_1_112), .B (n_5_107), .C1 (n_9_105), .C2 (n_12_105) );
AOI211_X1 g_3_109 (.ZN (n_3_109), .A (n_3_111), .B (n_4_109), .C1 (n_7_106), .C2 (n_10_106) );
AOI211_X1 g_4_107 (.ZN (n_4_107), .A (n_5_110), .B (n_2_110), .C1 (n_5_107), .C2 (n_11_104) );
AOI211_X1 g_6_108 (.ZN (n_6_108), .A (n_3_109), .B (n_1_112), .C1 (n_4_109), .C2 (n_9_105) );
AOI211_X1 g_8_107 (.ZN (n_8_107), .A (n_4_107), .B (n_3_111), .C1 (n_2_110), .C2 (n_7_106) );
AOI211_X1 g_6_106 (.ZN (n_6_106), .A (n_6_108), .B (n_5_110), .C1 (n_1_112), .C2 (n_5_107) );
AOI211_X1 g_8_105 (.ZN (n_8_105), .A (n_8_107), .B (n_3_109), .C1 (n_3_111), .C2 (n_4_109) );
AOI211_X1 g_7_107 (.ZN (n_7_107), .A (n_6_106), .B (n_4_107), .C1 (n_5_110), .C2 (n_2_110) );
AOI211_X1 g_9_106 (.ZN (n_9_106), .A (n_8_105), .B (n_6_108), .C1 (n_3_109), .C2 (n_1_112) );
AOI211_X1 g_8_108 (.ZN (n_8_108), .A (n_7_107), .B (n_8_107), .C1 (n_4_107), .C2 (n_3_111) );
AOI211_X1 g_6_107 (.ZN (n_6_107), .A (n_9_106), .B (n_6_106), .C1 (n_6_108), .C2 (n_5_110) );
AOI211_X1 g_8_106 (.ZN (n_8_106), .A (n_8_108), .B (n_8_105), .C1 (n_8_107), .C2 (n_3_109) );
AOI211_X1 g_10_105 (.ZN (n_10_105), .A (n_6_107), .B (n_7_107), .C1 (n_6_106), .C2 (n_4_107) );
AOI211_X1 g_12_104 (.ZN (n_12_104), .A (n_8_106), .B (n_9_106), .C1 (n_8_105), .C2 (n_6_108) );
AOI211_X1 g_14_103 (.ZN (n_14_103), .A (n_10_105), .B (n_8_108), .C1 (n_7_107), .C2 (n_8_107) );
AOI211_X1 g_16_102 (.ZN (n_16_102), .A (n_12_104), .B (n_6_107), .C1 (n_9_106), .C2 (n_6_106) );
AOI211_X1 g_18_101 (.ZN (n_18_101), .A (n_14_103), .B (n_8_106), .C1 (n_8_108), .C2 (n_8_105) );
AOI211_X1 g_20_100 (.ZN (n_20_100), .A (n_16_102), .B (n_10_105), .C1 (n_6_107), .C2 (n_7_107) );
AOI211_X1 g_22_99 (.ZN (n_22_99), .A (n_18_101), .B (n_12_104), .C1 (n_8_106), .C2 (n_9_106) );
AOI211_X1 g_24_98 (.ZN (n_24_98), .A (n_20_100), .B (n_14_103), .C1 (n_10_105), .C2 (n_8_108) );
AOI211_X1 g_26_97 (.ZN (n_26_97), .A (n_22_99), .B (n_16_102), .C1 (n_12_104), .C2 (n_6_107) );
AOI211_X1 g_28_96 (.ZN (n_28_96), .A (n_24_98), .B (n_18_101), .C1 (n_14_103), .C2 (n_8_106) );
AOI211_X1 g_30_95 (.ZN (n_30_95), .A (n_26_97), .B (n_20_100), .C1 (n_16_102), .C2 (n_10_105) );
AOI211_X1 g_32_96 (.ZN (n_32_96), .A (n_28_96), .B (n_22_99), .C1 (n_18_101), .C2 (n_12_104) );
AOI211_X1 g_30_97 (.ZN (n_30_97), .A (n_30_95), .B (n_24_98), .C1 (n_20_100), .C2 (n_14_103) );
AOI211_X1 g_28_98 (.ZN (n_28_98), .A (n_32_96), .B (n_26_97), .C1 (n_22_99), .C2 (n_16_102) );
AOI211_X1 g_26_99 (.ZN (n_26_99), .A (n_30_97), .B (n_28_96), .C1 (n_24_98), .C2 (n_18_101) );
AOI211_X1 g_24_100 (.ZN (n_24_100), .A (n_28_98), .B (n_30_95), .C1 (n_26_97), .C2 (n_20_100) );
AOI211_X1 g_25_98 (.ZN (n_25_98), .A (n_26_99), .B (n_32_96), .C1 (n_28_96), .C2 (n_22_99) );
AOI211_X1 g_23_99 (.ZN (n_23_99), .A (n_24_100), .B (n_30_97), .C1 (n_30_95), .C2 (n_24_98) );
AOI211_X1 g_21_100 (.ZN (n_21_100), .A (n_25_98), .B (n_28_98), .C1 (n_32_96), .C2 (n_26_97) );
AOI211_X1 g_19_101 (.ZN (n_19_101), .A (n_23_99), .B (n_26_99), .C1 (n_30_97), .C2 (n_28_96) );
AOI211_X1 g_17_102 (.ZN (n_17_102), .A (n_21_100), .B (n_24_100), .C1 (n_28_98), .C2 (n_30_95) );
AOI211_X1 g_15_103 (.ZN (n_15_103), .A (n_19_101), .B (n_25_98), .C1 (n_26_99), .C2 (n_32_96) );
AOI211_X1 g_13_104 (.ZN (n_13_104), .A (n_17_102), .B (n_23_99), .C1 (n_24_100), .C2 (n_30_97) );
AOI211_X1 g_12_106 (.ZN (n_12_106), .A (n_15_103), .B (n_21_100), .C1 (n_25_98), .C2 (n_28_98) );
AOI211_X1 g_10_107 (.ZN (n_10_107), .A (n_13_104), .B (n_19_101), .C1 (n_23_99), .C2 (n_26_99) );
AOI211_X1 g_9_109 (.ZN (n_9_109), .A (n_12_106), .B (n_17_102), .C1 (n_21_100), .C2 (n_24_100) );
AOI211_X1 g_7_108 (.ZN (n_7_108), .A (n_10_107), .B (n_15_103), .C1 (n_19_101), .C2 (n_25_98) );
AOI211_X1 g_5_109 (.ZN (n_5_109), .A (n_9_109), .B (n_13_104), .C1 (n_17_102), .C2 (n_23_99) );
AOI211_X1 g_4_111 (.ZN (n_4_111), .A (n_7_108), .B (n_12_106), .C1 (n_15_103), .C2 (n_21_100) );
AOI211_X1 g_3_113 (.ZN (n_3_113), .A (n_5_109), .B (n_10_107), .C1 (n_13_104), .C2 (n_19_101) );
AOI211_X1 g_5_114 (.ZN (n_5_114), .A (n_4_111), .B (n_9_109), .C1 (n_12_106), .C2 (n_17_102) );
AOI211_X1 g_3_115 (.ZN (n_3_115), .A (n_3_113), .B (n_7_108), .C1 (n_10_107), .C2 (n_15_103) );
AOI211_X1 g_1_116 (.ZN (n_1_116), .A (n_5_114), .B (n_5_109), .C1 (n_9_109), .C2 (n_13_104) );
AOI211_X1 g_2_114 (.ZN (n_2_114), .A (n_3_115), .B (n_4_111), .C1 (n_7_108), .C2 (n_12_106) );
AOI211_X1 g_4_113 (.ZN (n_4_113), .A (n_1_116), .B (n_3_113), .C1 (n_5_109), .C2 (n_10_107) );
AOI211_X1 g_6_112 (.ZN (n_6_112), .A (n_2_114), .B (n_5_114), .C1 (n_4_111), .C2 (n_9_109) );
AOI211_X1 g_7_110 (.ZN (n_7_110), .A (n_4_113), .B (n_3_115), .C1 (n_3_113), .C2 (n_7_108) );
AOI211_X1 g_5_111 (.ZN (n_5_111), .A (n_6_112), .B (n_1_116), .C1 (n_5_114), .C2 (n_5_109) );
AOI211_X1 g_6_109 (.ZN (n_6_109), .A (n_7_110), .B (n_2_114), .C1 (n_3_115), .C2 (n_4_111) );
AOI211_X1 g_4_110 (.ZN (n_4_110), .A (n_5_111), .B (n_4_113), .C1 (n_1_116), .C2 (n_3_113) );
AOI211_X1 g_5_108 (.ZN (n_5_108), .A (n_6_109), .B (n_6_112), .C1 (n_2_114), .C2 (n_5_114) );
AOI211_X1 g_6_110 (.ZN (n_6_110), .A (n_4_110), .B (n_7_110), .C1 (n_4_113), .C2 (n_3_115) );
AOI211_X1 g_5_112 (.ZN (n_5_112), .A (n_5_108), .B (n_5_111), .C1 (n_6_112), .C2 (n_1_116) );
AOI211_X1 g_7_111 (.ZN (n_7_111), .A (n_6_110), .B (n_6_109), .C1 (n_7_110), .C2 (n_2_114) );
AOI211_X1 g_8_109 (.ZN (n_8_109), .A (n_5_112), .B (n_4_110), .C1 (n_5_111), .C2 (n_4_113) );
AOI211_X1 g_9_107 (.ZN (n_9_107), .A (n_7_111), .B (n_5_108), .C1 (n_6_109), .C2 (n_6_112) );
AOI211_X1 g_11_106 (.ZN (n_11_106), .A (n_8_109), .B (n_6_110), .C1 (n_4_110), .C2 (n_7_110) );
AOI211_X1 g_13_105 (.ZN (n_13_105), .A (n_9_107), .B (n_5_112), .C1 (n_5_108), .C2 (n_5_111) );
AOI211_X1 g_15_104 (.ZN (n_15_104), .A (n_11_106), .B (n_7_111), .C1 (n_6_110), .C2 (n_6_109) );
AOI211_X1 g_17_103 (.ZN (n_17_103), .A (n_13_105), .B (n_8_109), .C1 (n_5_112), .C2 (n_4_110) );
AOI211_X1 g_19_102 (.ZN (n_19_102), .A (n_15_104), .B (n_9_107), .C1 (n_7_111), .C2 (n_5_108) );
AOI211_X1 g_21_101 (.ZN (n_21_101), .A (n_17_103), .B (n_11_106), .C1 (n_8_109), .C2 (n_6_110) );
AOI211_X1 g_23_100 (.ZN (n_23_100), .A (n_19_102), .B (n_13_105), .C1 (n_9_107), .C2 (n_5_112) );
AOI211_X1 g_25_99 (.ZN (n_25_99), .A (n_21_101), .B (n_15_104), .C1 (n_11_106), .C2 (n_7_111) );
AOI211_X1 g_27_98 (.ZN (n_27_98), .A (n_23_100), .B (n_17_103), .C1 (n_13_105), .C2 (n_8_109) );
AOI211_X1 g_29_97 (.ZN (n_29_97), .A (n_25_99), .B (n_19_102), .C1 (n_15_104), .C2 (n_9_107) );
AOI211_X1 g_31_96 (.ZN (n_31_96), .A (n_27_98), .B (n_21_101), .C1 (n_17_103), .C2 (n_11_106) );
AOI211_X1 g_33_95 (.ZN (n_33_95), .A (n_29_97), .B (n_23_100), .C1 (n_19_102), .C2 (n_13_105) );
AOI211_X1 g_32_97 (.ZN (n_32_97), .A (n_31_96), .B (n_25_99), .C1 (n_21_101), .C2 (n_15_104) );
AOI211_X1 g_34_96 (.ZN (n_34_96), .A (n_33_95), .B (n_27_98), .C1 (n_23_100), .C2 (n_17_103) );
AOI211_X1 g_36_95 (.ZN (n_36_95), .A (n_32_97), .B (n_29_97), .C1 (n_25_99), .C2 (n_19_102) );
AOI211_X1 g_38_94 (.ZN (n_38_94), .A (n_34_96), .B (n_31_96), .C1 (n_27_98), .C2 (n_21_101) );
AOI211_X1 g_40_93 (.ZN (n_40_93), .A (n_36_95), .B (n_33_95), .C1 (n_29_97), .C2 (n_23_100) );
AOI211_X1 g_42_92 (.ZN (n_42_92), .A (n_38_94), .B (n_32_97), .C1 (n_31_96), .C2 (n_25_99) );
AOI211_X1 g_44_93 (.ZN (n_44_93), .A (n_40_93), .B (n_34_96), .C1 (n_33_95), .C2 (n_27_98) );
AOI211_X1 g_46_92 (.ZN (n_46_92), .A (n_42_92), .B (n_36_95), .C1 (n_32_97), .C2 (n_29_97) );
AOI211_X1 g_48_91 (.ZN (n_48_91), .A (n_44_93), .B (n_38_94), .C1 (n_34_96), .C2 (n_31_96) );
AOI211_X1 g_50_90 (.ZN (n_50_90), .A (n_46_92), .B (n_40_93), .C1 (n_36_95), .C2 (n_33_95) );
AOI211_X1 g_52_89 (.ZN (n_52_89), .A (n_48_91), .B (n_42_92), .C1 (n_38_94), .C2 (n_32_97) );
AOI211_X1 g_54_88 (.ZN (n_54_88), .A (n_50_90), .B (n_44_93), .C1 (n_40_93), .C2 (n_34_96) );
AOI211_X1 g_56_87 (.ZN (n_56_87), .A (n_52_89), .B (n_46_92), .C1 (n_42_92), .C2 (n_36_95) );
AOI211_X1 g_58_86 (.ZN (n_58_86), .A (n_54_88), .B (n_48_91), .C1 (n_44_93), .C2 (n_38_94) );
AOI211_X1 g_60_87 (.ZN (n_60_87), .A (n_56_87), .B (n_50_90), .C1 (n_46_92), .C2 (n_40_93) );
AOI211_X1 g_61_85 (.ZN (n_61_85), .A (n_58_86), .B (n_52_89), .C1 (n_48_91), .C2 (n_42_92) );
AOI211_X1 g_63_84 (.ZN (n_63_84), .A (n_60_87), .B (n_54_88), .C1 (n_50_90), .C2 (n_44_93) );
AOI211_X1 g_65_83 (.ZN (n_65_83), .A (n_61_85), .B (n_56_87), .C1 (n_52_89), .C2 (n_46_92) );
AOI211_X1 g_67_82 (.ZN (n_67_82), .A (n_63_84), .B (n_58_86), .C1 (n_54_88), .C2 (n_48_91) );
AOI211_X1 g_69_81 (.ZN (n_69_81), .A (n_65_83), .B (n_60_87), .C1 (n_56_87), .C2 (n_50_90) );
AOI211_X1 g_71_80 (.ZN (n_71_80), .A (n_67_82), .B (n_61_85), .C1 (n_58_86), .C2 (n_52_89) );
AOI211_X1 g_73_79 (.ZN (n_73_79), .A (n_69_81), .B (n_63_84), .C1 (n_60_87), .C2 (n_54_88) );
AOI211_X1 g_75_78 (.ZN (n_75_78), .A (n_71_80), .B (n_65_83), .C1 (n_61_85), .C2 (n_56_87) );
AOI211_X1 g_77_77 (.ZN (n_77_77), .A (n_73_79), .B (n_67_82), .C1 (n_63_84), .C2 (n_58_86) );
AOI211_X1 g_79_76 (.ZN (n_79_76), .A (n_75_78), .B (n_69_81), .C1 (n_65_83), .C2 (n_60_87) );
AOI211_X1 g_81_75 (.ZN (n_81_75), .A (n_77_77), .B (n_71_80), .C1 (n_67_82), .C2 (n_61_85) );
AOI211_X1 g_83_74 (.ZN (n_83_74), .A (n_79_76), .B (n_73_79), .C1 (n_69_81), .C2 (n_63_84) );
AOI211_X1 g_82_76 (.ZN (n_82_76), .A (n_81_75), .B (n_75_78), .C1 (n_71_80), .C2 (n_65_83) );
AOI211_X1 g_84_75 (.ZN (n_84_75), .A (n_83_74), .B (n_77_77), .C1 (n_73_79), .C2 (n_67_82) );
AOI211_X1 g_86_74 (.ZN (n_86_74), .A (n_82_76), .B (n_79_76), .C1 (n_75_78), .C2 (n_69_81) );
AOI211_X1 g_88_73 (.ZN (n_88_73), .A (n_84_75), .B (n_81_75), .C1 (n_77_77), .C2 (n_71_80) );
AOI211_X1 g_87_75 (.ZN (n_87_75), .A (n_86_74), .B (n_83_74), .C1 (n_79_76), .C2 (n_73_79) );
AOI211_X1 g_86_73 (.ZN (n_86_73), .A (n_88_73), .B (n_82_76), .C1 (n_81_75), .C2 (n_75_78) );
AOI211_X1 g_88_72 (.ZN (n_88_72), .A (n_87_75), .B (n_84_75), .C1 (n_83_74), .C2 (n_77_77) );
AOI211_X1 g_90_71 (.ZN (n_90_71), .A (n_86_73), .B (n_86_74), .C1 (n_82_76), .C2 (n_79_76) );
AOI211_X1 g_92_72 (.ZN (n_92_72), .A (n_88_72), .B (n_88_73), .C1 (n_84_75), .C2 (n_81_75) );
AOI211_X1 g_90_73 (.ZN (n_90_73), .A (n_90_71), .B (n_87_75), .C1 (n_86_74), .C2 (n_83_74) );
AOI211_X1 g_88_74 (.ZN (n_88_74), .A (n_92_72), .B (n_86_73), .C1 (n_88_73), .C2 (n_82_76) );
AOI211_X1 g_86_75 (.ZN (n_86_75), .A (n_90_73), .B (n_88_72), .C1 (n_87_75), .C2 (n_84_75) );
AOI211_X1 g_84_74 (.ZN (n_84_74), .A (n_88_74), .B (n_90_71), .C1 (n_86_73), .C2 (n_86_74) );
AOI211_X1 g_82_75 (.ZN (n_82_75), .A (n_86_75), .B (n_92_72), .C1 (n_88_72), .C2 (n_88_73) );
AOI211_X1 g_80_76 (.ZN (n_80_76), .A (n_84_74), .B (n_90_73), .C1 (n_90_71), .C2 (n_87_75) );
AOI211_X1 g_78_77 (.ZN (n_78_77), .A (n_82_75), .B (n_88_74), .C1 (n_92_72), .C2 (n_86_73) );
AOI211_X1 g_76_78 (.ZN (n_76_78), .A (n_80_76), .B (n_86_75), .C1 (n_90_73), .C2 (n_88_72) );
AOI211_X1 g_74_79 (.ZN (n_74_79), .A (n_78_77), .B (n_84_74), .C1 (n_88_74), .C2 (n_90_71) );
AOI211_X1 g_72_80 (.ZN (n_72_80), .A (n_76_78), .B (n_82_75), .C1 (n_86_75), .C2 (n_92_72) );
AOI211_X1 g_70_81 (.ZN (n_70_81), .A (n_74_79), .B (n_80_76), .C1 (n_84_74), .C2 (n_90_73) );
AOI211_X1 g_68_82 (.ZN (n_68_82), .A (n_72_80), .B (n_78_77), .C1 (n_82_75), .C2 (n_88_74) );
AOI211_X1 g_66_83 (.ZN (n_66_83), .A (n_70_81), .B (n_76_78), .C1 (n_80_76), .C2 (n_86_75) );
AOI211_X1 g_64_84 (.ZN (n_64_84), .A (n_68_82), .B (n_74_79), .C1 (n_78_77), .C2 (n_84_74) );
AOI211_X1 g_62_85 (.ZN (n_62_85), .A (n_66_83), .B (n_72_80), .C1 (n_76_78), .C2 (n_82_75) );
AOI211_X1 g_60_86 (.ZN (n_60_86), .A (n_64_84), .B (n_70_81), .C1 (n_74_79), .C2 (n_80_76) );
AOI211_X1 g_58_85 (.ZN (n_58_85), .A (n_62_85), .B (n_68_82), .C1 (n_72_80), .C2 (n_78_77) );
AOI211_X1 g_56_86 (.ZN (n_56_86), .A (n_60_86), .B (n_66_83), .C1 (n_70_81), .C2 (n_76_78) );
AOI211_X1 g_54_87 (.ZN (n_54_87), .A (n_58_85), .B (n_64_84), .C1 (n_68_82), .C2 (n_74_79) );
AOI211_X1 g_52_88 (.ZN (n_52_88), .A (n_56_86), .B (n_62_85), .C1 (n_66_83), .C2 (n_72_80) );
AOI211_X1 g_50_89 (.ZN (n_50_89), .A (n_54_87), .B (n_60_86), .C1 (n_64_84), .C2 (n_70_81) );
AOI211_X1 g_48_90 (.ZN (n_48_90), .A (n_52_88), .B (n_58_85), .C1 (n_62_85), .C2 (n_68_82) );
AOI211_X1 g_46_91 (.ZN (n_46_91), .A (n_50_89), .B (n_56_86), .C1 (n_60_86), .C2 (n_66_83) );
AOI211_X1 g_44_92 (.ZN (n_44_92), .A (n_48_90), .B (n_54_87), .C1 (n_58_85), .C2 (n_64_84) );
AOI211_X1 g_42_93 (.ZN (n_42_93), .A (n_46_91), .B (n_52_88), .C1 (n_56_86), .C2 (n_62_85) );
AOI211_X1 g_40_92 (.ZN (n_40_92), .A (n_44_92), .B (n_50_89), .C1 (n_54_87), .C2 (n_60_86) );
AOI211_X1 g_38_93 (.ZN (n_38_93), .A (n_42_93), .B (n_48_90), .C1 (n_52_88), .C2 (n_58_85) );
AOI211_X1 g_36_94 (.ZN (n_36_94), .A (n_40_92), .B (n_46_91), .C1 (n_50_89), .C2 (n_56_86) );
AOI211_X1 g_35_96 (.ZN (n_35_96), .A (n_38_93), .B (n_44_92), .C1 (n_48_90), .C2 (n_54_87) );
AOI211_X1 g_37_95 (.ZN (n_37_95), .A (n_36_94), .B (n_42_93), .C1 (n_46_91), .C2 (n_52_88) );
AOI211_X1 g_39_94 (.ZN (n_39_94), .A (n_35_96), .B (n_40_92), .C1 (n_44_92), .C2 (n_50_89) );
AOI211_X1 g_41_95 (.ZN (n_41_95), .A (n_37_95), .B (n_38_93), .C1 (n_42_93), .C2 (n_48_90) );
AOI211_X1 g_43_94 (.ZN (n_43_94), .A (n_39_94), .B (n_36_94), .C1 (n_40_92), .C2 (n_46_91) );
AOI211_X1 g_45_93 (.ZN (n_45_93), .A (n_41_95), .B (n_35_96), .C1 (n_38_93), .C2 (n_44_92) );
AOI211_X1 g_47_92 (.ZN (n_47_92), .A (n_43_94), .B (n_37_95), .C1 (n_36_94), .C2 (n_42_93) );
AOI211_X1 g_49_91 (.ZN (n_49_91), .A (n_45_93), .B (n_39_94), .C1 (n_35_96), .C2 (n_40_92) );
AOI211_X1 g_51_90 (.ZN (n_51_90), .A (n_47_92), .B (n_41_95), .C1 (n_37_95), .C2 (n_38_93) );
AOI211_X1 g_53_89 (.ZN (n_53_89), .A (n_49_91), .B (n_43_94), .C1 (n_39_94), .C2 (n_36_94) );
AOI211_X1 g_55_88 (.ZN (n_55_88), .A (n_51_90), .B (n_45_93), .C1 (n_41_95), .C2 (n_35_96) );
AOI211_X1 g_57_87 (.ZN (n_57_87), .A (n_53_89), .B (n_47_92), .C1 (n_43_94), .C2 (n_37_95) );
AOI211_X1 g_59_86 (.ZN (n_59_86), .A (n_55_88), .B (n_49_91), .C1 (n_45_93), .C2 (n_39_94) );
AOI211_X1 g_58_88 (.ZN (n_58_88), .A (n_57_87), .B (n_51_90), .C1 (n_47_92), .C2 (n_41_95) );
AOI211_X1 g_57_86 (.ZN (n_57_86), .A (n_59_86), .B (n_53_89), .C1 (n_49_91), .C2 (n_43_94) );
AOI211_X1 g_55_87 (.ZN (n_55_87), .A (n_58_88), .B (n_55_88), .C1 (n_51_90), .C2 (n_45_93) );
AOI211_X1 g_53_88 (.ZN (n_53_88), .A (n_57_86), .B (n_57_87), .C1 (n_53_89), .C2 (n_47_92) );
AOI211_X1 g_51_89 (.ZN (n_51_89), .A (n_55_87), .B (n_59_86), .C1 (n_55_88), .C2 (n_49_91) );
AOI211_X1 g_49_90 (.ZN (n_49_90), .A (n_53_88), .B (n_58_88), .C1 (n_57_87), .C2 (n_51_90) );
AOI211_X1 g_47_91 (.ZN (n_47_91), .A (n_51_89), .B (n_57_86), .C1 (n_59_86), .C2 (n_53_89) );
AOI211_X1 g_46_93 (.ZN (n_46_93), .A (n_49_90), .B (n_55_87), .C1 (n_58_88), .C2 (n_55_88) );
AOI211_X1 g_48_92 (.ZN (n_48_92), .A (n_47_91), .B (n_53_88), .C1 (n_57_86), .C2 (n_57_87) );
AOI211_X1 g_50_91 (.ZN (n_50_91), .A (n_46_93), .B (n_51_89), .C1 (n_55_87), .C2 (n_59_86) );
AOI211_X1 g_52_90 (.ZN (n_52_90), .A (n_48_92), .B (n_49_90), .C1 (n_53_88), .C2 (n_58_88) );
AOI211_X1 g_54_89 (.ZN (n_54_89), .A (n_50_91), .B (n_47_91), .C1 (n_51_89), .C2 (n_57_86) );
AOI211_X1 g_56_88 (.ZN (n_56_88), .A (n_52_90), .B (n_46_93), .C1 (n_49_90), .C2 (n_55_87) );
AOI211_X1 g_58_87 (.ZN (n_58_87), .A (n_54_89), .B (n_48_92), .C1 (n_47_91), .C2 (n_53_88) );
AOI211_X1 g_57_89 (.ZN (n_57_89), .A (n_56_88), .B (n_50_91), .C1 (n_46_93), .C2 (n_51_89) );
AOI211_X1 g_59_88 (.ZN (n_59_88), .A (n_58_87), .B (n_52_90), .C1 (n_48_92), .C2 (n_49_90) );
AOI211_X1 g_61_87 (.ZN (n_61_87), .A (n_57_89), .B (n_54_89), .C1 (n_50_91), .C2 (n_47_91) );
AOI211_X1 g_63_86 (.ZN (n_63_86), .A (n_59_88), .B (n_56_88), .C1 (n_52_90), .C2 (n_46_93) );
AOI211_X1 g_65_85 (.ZN (n_65_85), .A (n_61_87), .B (n_58_87), .C1 (n_54_89), .C2 (n_48_92) );
AOI211_X1 g_67_84 (.ZN (n_67_84), .A (n_63_86), .B (n_57_89), .C1 (n_56_88), .C2 (n_50_91) );
AOI211_X1 g_69_83 (.ZN (n_69_83), .A (n_65_85), .B (n_59_88), .C1 (n_58_87), .C2 (n_52_90) );
AOI211_X1 g_71_82 (.ZN (n_71_82), .A (n_67_84), .B (n_61_87), .C1 (n_57_89), .C2 (n_54_89) );
AOI211_X1 g_73_81 (.ZN (n_73_81), .A (n_69_83), .B (n_63_86), .C1 (n_59_88), .C2 (n_56_88) );
AOI211_X1 g_75_80 (.ZN (n_75_80), .A (n_71_82), .B (n_65_85), .C1 (n_61_87), .C2 (n_58_87) );
AOI211_X1 g_77_79 (.ZN (n_77_79), .A (n_73_81), .B (n_67_84), .C1 (n_63_86), .C2 (n_57_89) );
AOI211_X1 g_79_78 (.ZN (n_79_78), .A (n_75_80), .B (n_69_83), .C1 (n_65_85), .C2 (n_59_88) );
AOI211_X1 g_81_77 (.ZN (n_81_77), .A (n_77_79), .B (n_71_82), .C1 (n_67_84), .C2 (n_61_87) );
AOI211_X1 g_83_76 (.ZN (n_83_76), .A (n_79_78), .B (n_73_81), .C1 (n_69_83), .C2 (n_63_86) );
AOI211_X1 g_85_75 (.ZN (n_85_75), .A (n_81_77), .B (n_75_80), .C1 (n_71_82), .C2 (n_65_85) );
AOI211_X1 g_87_74 (.ZN (n_87_74), .A (n_83_76), .B (n_77_79), .C1 (n_73_81), .C2 (n_67_84) );
AOI211_X1 g_89_73 (.ZN (n_89_73), .A (n_85_75), .B (n_79_78), .C1 (n_75_80), .C2 (n_69_83) );
AOI211_X1 g_91_72 (.ZN (n_91_72), .A (n_87_74), .B (n_81_77), .C1 (n_77_79), .C2 (n_71_82) );
AOI211_X1 g_93_71 (.ZN (n_93_71), .A (n_89_73), .B (n_83_76), .C1 (n_79_78), .C2 (n_73_81) );
AOI211_X1 g_92_73 (.ZN (n_92_73), .A (n_91_72), .B (n_85_75), .C1 (n_81_77), .C2 (n_75_80) );
AOI211_X1 g_90_74 (.ZN (n_90_74), .A (n_93_71), .B (n_87_74), .C1 (n_83_76), .C2 (n_77_79) );
AOI211_X1 g_88_75 (.ZN (n_88_75), .A (n_92_73), .B (n_89_73), .C1 (n_85_75), .C2 (n_79_78) );
AOI211_X1 g_86_76 (.ZN (n_86_76), .A (n_90_74), .B (n_91_72), .C1 (n_87_74), .C2 (n_81_77) );
AOI211_X1 g_84_77 (.ZN (n_84_77), .A (n_88_75), .B (n_93_71), .C1 (n_89_73), .C2 (n_83_76) );
AOI211_X1 g_83_75 (.ZN (n_83_75), .A (n_86_76), .B (n_92_73), .C1 (n_91_72), .C2 (n_85_75) );
AOI211_X1 g_81_76 (.ZN (n_81_76), .A (n_84_77), .B (n_90_74), .C1 (n_93_71), .C2 (n_87_74) );
AOI211_X1 g_79_77 (.ZN (n_79_77), .A (n_83_75), .B (n_88_75), .C1 (n_92_73), .C2 (n_89_73) );
AOI211_X1 g_77_78 (.ZN (n_77_78), .A (n_81_76), .B (n_86_76), .C1 (n_90_74), .C2 (n_91_72) );
AOI211_X1 g_75_79 (.ZN (n_75_79), .A (n_79_77), .B (n_84_77), .C1 (n_88_75), .C2 (n_93_71) );
AOI211_X1 g_73_80 (.ZN (n_73_80), .A (n_77_78), .B (n_83_75), .C1 (n_86_76), .C2 (n_92_73) );
AOI211_X1 g_71_81 (.ZN (n_71_81), .A (n_75_79), .B (n_81_76), .C1 (n_84_77), .C2 (n_90_74) );
AOI211_X1 g_69_82 (.ZN (n_69_82), .A (n_73_80), .B (n_79_77), .C1 (n_83_75), .C2 (n_88_75) );
AOI211_X1 g_67_83 (.ZN (n_67_83), .A (n_71_81), .B (n_77_78), .C1 (n_81_76), .C2 (n_86_76) );
AOI211_X1 g_65_84 (.ZN (n_65_84), .A (n_69_82), .B (n_75_79), .C1 (n_79_77), .C2 (n_84_77) );
AOI211_X1 g_63_85 (.ZN (n_63_85), .A (n_67_83), .B (n_73_80), .C1 (n_77_78), .C2 (n_83_75) );
AOI211_X1 g_61_86 (.ZN (n_61_86), .A (n_65_84), .B (n_71_81), .C1 (n_75_79), .C2 (n_81_76) );
AOI211_X1 g_59_87 (.ZN (n_59_87), .A (n_63_85), .B (n_69_82), .C1 (n_73_80), .C2 (n_79_77) );
AOI211_X1 g_57_88 (.ZN (n_57_88), .A (n_61_86), .B (n_67_83), .C1 (n_71_81), .C2 (n_77_78) );
AOI211_X1 g_55_89 (.ZN (n_55_89), .A (n_59_87), .B (n_65_84), .C1 (n_69_82), .C2 (n_75_79) );
AOI211_X1 g_53_90 (.ZN (n_53_90), .A (n_57_88), .B (n_63_85), .C1 (n_67_83), .C2 (n_73_80) );
AOI211_X1 g_51_91 (.ZN (n_51_91), .A (n_55_89), .B (n_61_86), .C1 (n_65_84), .C2 (n_71_81) );
AOI211_X1 g_49_92 (.ZN (n_49_92), .A (n_53_90), .B (n_59_87), .C1 (n_63_85), .C2 (n_69_82) );
AOI211_X1 g_47_93 (.ZN (n_47_93), .A (n_51_91), .B (n_57_88), .C1 (n_61_86), .C2 (n_67_83) );
AOI211_X1 g_45_94 (.ZN (n_45_94), .A (n_49_92), .B (n_55_89), .C1 (n_59_87), .C2 (n_65_84) );
AOI211_X1 g_43_93 (.ZN (n_43_93), .A (n_47_93), .B (n_53_90), .C1 (n_57_88), .C2 (n_63_85) );
AOI211_X1 g_41_92 (.ZN (n_41_92), .A (n_45_94), .B (n_51_91), .C1 (n_55_89), .C2 (n_61_86) );
AOI211_X1 g_39_93 (.ZN (n_39_93), .A (n_43_93), .B (n_49_92), .C1 (n_53_90), .C2 (n_59_87) );
AOI211_X1 g_37_94 (.ZN (n_37_94), .A (n_41_92), .B (n_47_93), .C1 (n_51_91), .C2 (n_57_88) );
AOI211_X1 g_35_95 (.ZN (n_35_95), .A (n_39_93), .B (n_45_94), .C1 (n_49_92), .C2 (n_55_89) );
AOI211_X1 g_33_96 (.ZN (n_33_96), .A (n_37_94), .B (n_43_93), .C1 (n_47_93), .C2 (n_53_90) );
AOI211_X1 g_31_97 (.ZN (n_31_97), .A (n_35_95), .B (n_41_92), .C1 (n_45_94), .C2 (n_51_91) );
AOI211_X1 g_29_98 (.ZN (n_29_98), .A (n_33_96), .B (n_39_93), .C1 (n_43_93), .C2 (n_49_92) );
AOI211_X1 g_27_99 (.ZN (n_27_99), .A (n_31_97), .B (n_37_94), .C1 (n_41_92), .C2 (n_47_93) );
AOI211_X1 g_25_100 (.ZN (n_25_100), .A (n_29_98), .B (n_35_95), .C1 (n_39_93), .C2 (n_45_94) );
AOI211_X1 g_23_101 (.ZN (n_23_101), .A (n_27_99), .B (n_33_96), .C1 (n_37_94), .C2 (n_43_93) );
AOI211_X1 g_21_102 (.ZN (n_21_102), .A (n_25_100), .B (n_31_97), .C1 (n_35_95), .C2 (n_41_92) );
AOI211_X1 g_19_103 (.ZN (n_19_103), .A (n_23_101), .B (n_29_98), .C1 (n_33_96), .C2 (n_39_93) );
AOI211_X1 g_17_104 (.ZN (n_17_104), .A (n_21_102), .B (n_27_99), .C1 (n_31_97), .C2 (n_37_94) );
AOI211_X1 g_15_105 (.ZN (n_15_105), .A (n_19_103), .B (n_25_100), .C1 (n_29_98), .C2 (n_35_95) );
AOI211_X1 g_13_106 (.ZN (n_13_106), .A (n_17_104), .B (n_23_101), .C1 (n_27_99), .C2 (n_33_96) );
AOI211_X1 g_11_107 (.ZN (n_11_107), .A (n_15_105), .B (n_21_102), .C1 (n_25_100), .C2 (n_31_97) );
AOI211_X1 g_9_108 (.ZN (n_9_108), .A (n_13_106), .B (n_19_103), .C1 (n_23_101), .C2 (n_29_98) );
AOI211_X1 g_7_109 (.ZN (n_7_109), .A (n_11_107), .B (n_17_104), .C1 (n_21_102), .C2 (n_27_99) );
AOI211_X1 g_6_111 (.ZN (n_6_111), .A (n_9_108), .B (n_15_105), .C1 (n_19_103), .C2 (n_25_100) );
AOI211_X1 g_8_110 (.ZN (n_8_110), .A (n_7_109), .B (n_13_106), .C1 (n_17_104), .C2 (n_23_101) );
AOI211_X1 g_10_109 (.ZN (n_10_109), .A (n_6_111), .B (n_11_107), .C1 (n_15_105), .C2 (n_21_102) );
AOI211_X1 g_12_108 (.ZN (n_12_108), .A (n_8_110), .B (n_9_108), .C1 (n_13_106), .C2 (n_19_103) );
AOI211_X1 g_14_107 (.ZN (n_14_107), .A (n_10_109), .B (n_7_109), .C1 (n_11_107), .C2 (n_17_104) );
AOI211_X1 g_16_106 (.ZN (n_16_106), .A (n_12_108), .B (n_6_111), .C1 (n_9_108), .C2 (n_15_105) );
AOI211_X1 g_14_105 (.ZN (n_14_105), .A (n_14_107), .B (n_8_110), .C1 (n_7_109), .C2 (n_13_106) );
AOI211_X1 g_16_104 (.ZN (n_16_104), .A (n_16_106), .B (n_10_109), .C1 (n_6_111), .C2 (n_11_107) );
AOI211_X1 g_18_103 (.ZN (n_18_103), .A (n_14_105), .B (n_12_108), .C1 (n_8_110), .C2 (n_9_108) );
AOI211_X1 g_20_102 (.ZN (n_20_102), .A (n_16_104), .B (n_14_107), .C1 (n_10_109), .C2 (n_7_109) );
AOI211_X1 g_22_101 (.ZN (n_22_101), .A (n_18_103), .B (n_16_106), .C1 (n_12_108), .C2 (n_6_111) );
AOI211_X1 g_21_103 (.ZN (n_21_103), .A (n_20_102), .B (n_14_105), .C1 (n_14_107), .C2 (n_8_110) );
AOI211_X1 g_23_102 (.ZN (n_23_102), .A (n_22_101), .B (n_16_104), .C1 (n_16_106), .C2 (n_10_109) );
AOI211_X1 g_25_101 (.ZN (n_25_101), .A (n_21_103), .B (n_18_103), .C1 (n_14_105), .C2 (n_12_108) );
AOI211_X1 g_27_100 (.ZN (n_27_100), .A (n_23_102), .B (n_20_102), .C1 (n_16_104), .C2 (n_14_107) );
AOI211_X1 g_29_99 (.ZN (n_29_99), .A (n_25_101), .B (n_22_101), .C1 (n_18_103), .C2 (n_16_106) );
AOI211_X1 g_31_98 (.ZN (n_31_98), .A (n_27_100), .B (n_21_103), .C1 (n_20_102), .C2 (n_14_105) );
AOI211_X1 g_33_97 (.ZN (n_33_97), .A (n_29_99), .B (n_23_102), .C1 (n_22_101), .C2 (n_16_104) );
AOI211_X1 g_32_99 (.ZN (n_32_99), .A (n_31_98), .B (n_25_101), .C1 (n_21_103), .C2 (n_18_103) );
AOI211_X1 g_30_98 (.ZN (n_30_98), .A (n_33_97), .B (n_27_100), .C1 (n_23_102), .C2 (n_20_102) );
AOI211_X1 g_28_99 (.ZN (n_28_99), .A (n_32_99), .B (n_29_99), .C1 (n_25_101), .C2 (n_22_101) );
AOI211_X1 g_26_100 (.ZN (n_26_100), .A (n_30_98), .B (n_31_98), .C1 (n_27_100), .C2 (n_21_103) );
AOI211_X1 g_24_101 (.ZN (n_24_101), .A (n_28_99), .B (n_33_97), .C1 (n_29_99), .C2 (n_23_102) );
AOI211_X1 g_22_102 (.ZN (n_22_102), .A (n_26_100), .B (n_32_99), .C1 (n_31_98), .C2 (n_25_101) );
AOI211_X1 g_20_103 (.ZN (n_20_103), .A (n_24_101), .B (n_30_98), .C1 (n_33_97), .C2 (n_27_100) );
AOI211_X1 g_18_104 (.ZN (n_18_104), .A (n_22_102), .B (n_28_99), .C1 (n_32_99), .C2 (n_29_99) );
AOI211_X1 g_16_105 (.ZN (n_16_105), .A (n_20_103), .B (n_26_100), .C1 (n_30_98), .C2 (n_31_98) );
AOI211_X1 g_14_106 (.ZN (n_14_106), .A (n_18_104), .B (n_24_101), .C1 (n_28_99), .C2 (n_33_97) );
AOI211_X1 g_12_107 (.ZN (n_12_107), .A (n_16_105), .B (n_22_102), .C1 (n_26_100), .C2 (n_32_99) );
AOI211_X1 g_10_108 (.ZN (n_10_108), .A (n_14_106), .B (n_20_103), .C1 (n_24_101), .C2 (n_30_98) );
AOI211_X1 g_9_110 (.ZN (n_9_110), .A (n_12_107), .B (n_18_104), .C1 (n_22_102), .C2 (n_28_99) );
AOI211_X1 g_11_109 (.ZN (n_11_109), .A (n_10_108), .B (n_16_105), .C1 (n_20_103), .C2 (n_26_100) );
AOI211_X1 g_13_108 (.ZN (n_13_108), .A (n_9_110), .B (n_14_106), .C1 (n_18_104), .C2 (n_24_101) );
AOI211_X1 g_15_107 (.ZN (n_15_107), .A (n_11_109), .B (n_12_107), .C1 (n_16_105), .C2 (n_22_102) );
AOI211_X1 g_17_106 (.ZN (n_17_106), .A (n_13_108), .B (n_10_108), .C1 (n_14_106), .C2 (n_20_103) );
AOI211_X1 g_19_105 (.ZN (n_19_105), .A (n_15_107), .B (n_9_110), .C1 (n_12_107), .C2 (n_18_104) );
AOI211_X1 g_21_104 (.ZN (n_21_104), .A (n_17_106), .B (n_11_109), .C1 (n_10_108), .C2 (n_16_105) );
AOI211_X1 g_23_103 (.ZN (n_23_103), .A (n_19_105), .B (n_13_108), .C1 (n_9_110), .C2 (n_14_106) );
AOI211_X1 g_25_102 (.ZN (n_25_102), .A (n_21_104), .B (n_15_107), .C1 (n_11_109), .C2 (n_12_107) );
AOI211_X1 g_27_101 (.ZN (n_27_101), .A (n_23_103), .B (n_17_106), .C1 (n_13_108), .C2 (n_10_108) );
AOI211_X1 g_29_100 (.ZN (n_29_100), .A (n_25_102), .B (n_19_105), .C1 (n_15_107), .C2 (n_9_110) );
AOI211_X1 g_31_99 (.ZN (n_31_99), .A (n_27_101), .B (n_21_104), .C1 (n_17_106), .C2 (n_11_109) );
AOI211_X1 g_33_98 (.ZN (n_33_98), .A (n_29_100), .B (n_23_103), .C1 (n_19_105), .C2 (n_13_108) );
AOI211_X1 g_35_97 (.ZN (n_35_97), .A (n_31_99), .B (n_25_102), .C1 (n_21_104), .C2 (n_15_107) );
AOI211_X1 g_37_96 (.ZN (n_37_96), .A (n_33_98), .B (n_27_101), .C1 (n_23_103), .C2 (n_17_106) );
AOI211_X1 g_39_95 (.ZN (n_39_95), .A (n_35_97), .B (n_29_100), .C1 (n_25_102), .C2 (n_19_105) );
AOI211_X1 g_41_94 (.ZN (n_41_94), .A (n_37_96), .B (n_31_99), .C1 (n_27_101), .C2 (n_21_104) );
AOI211_X1 g_43_95 (.ZN (n_43_95), .A (n_39_95), .B (n_33_98), .C1 (n_29_100), .C2 (n_23_103) );
AOI211_X1 g_41_96 (.ZN (n_41_96), .A (n_41_94), .B (n_35_97), .C1 (n_31_99), .C2 (n_25_102) );
AOI211_X1 g_42_94 (.ZN (n_42_94), .A (n_43_95), .B (n_37_96), .C1 (n_33_98), .C2 (n_27_101) );
AOI211_X1 g_40_95 (.ZN (n_40_95), .A (n_41_96), .B (n_39_95), .C1 (n_35_97), .C2 (n_29_100) );
AOI211_X1 g_38_96 (.ZN (n_38_96), .A (n_42_94), .B (n_41_94), .C1 (n_37_96), .C2 (n_31_99) );
AOI211_X1 g_36_97 (.ZN (n_36_97), .A (n_40_95), .B (n_43_95), .C1 (n_39_95), .C2 (n_33_98) );
AOI211_X1 g_34_98 (.ZN (n_34_98), .A (n_38_96), .B (n_41_96), .C1 (n_41_94), .C2 (n_35_97) );
AOI211_X1 g_33_100 (.ZN (n_33_100), .A (n_36_97), .B (n_42_94), .C1 (n_43_95), .C2 (n_37_96) );
AOI211_X1 g_32_98 (.ZN (n_32_98), .A (n_34_98), .B (n_40_95), .C1 (n_41_96), .C2 (n_39_95) );
AOI211_X1 g_34_97 (.ZN (n_34_97), .A (n_33_100), .B (n_38_96), .C1 (n_42_94), .C2 (n_41_94) );
AOI211_X1 g_36_96 (.ZN (n_36_96), .A (n_32_98), .B (n_36_97), .C1 (n_40_95), .C2 (n_43_95) );
AOI211_X1 g_38_95 (.ZN (n_38_95), .A (n_34_97), .B (n_34_98), .C1 (n_38_96), .C2 (n_41_96) );
AOI211_X1 g_40_94 (.ZN (n_40_94), .A (n_36_96), .B (n_33_100), .C1 (n_36_97), .C2 (n_42_94) );
AOI211_X1 g_39_96 (.ZN (n_39_96), .A (n_38_95), .B (n_32_98), .C1 (n_34_98), .C2 (n_40_95) );
AOI211_X1 g_37_97 (.ZN (n_37_97), .A (n_40_94), .B (n_34_97), .C1 (n_33_100), .C2 (n_38_96) );
AOI211_X1 g_35_98 (.ZN (n_35_98), .A (n_39_96), .B (n_36_96), .C1 (n_32_98), .C2 (n_36_97) );
AOI211_X1 g_33_99 (.ZN (n_33_99), .A (n_37_97), .B (n_38_95), .C1 (n_34_97), .C2 (n_34_98) );
AOI211_X1 g_31_100 (.ZN (n_31_100), .A (n_35_98), .B (n_40_94), .C1 (n_36_96), .C2 (n_33_100) );
AOI211_X1 g_29_101 (.ZN (n_29_101), .A (n_33_99), .B (n_39_96), .C1 (n_38_95), .C2 (n_32_98) );
AOI211_X1 g_30_99 (.ZN (n_30_99), .A (n_31_100), .B (n_37_97), .C1 (n_40_94), .C2 (n_34_97) );
AOI211_X1 g_28_100 (.ZN (n_28_100), .A (n_29_101), .B (n_35_98), .C1 (n_39_96), .C2 (n_36_96) );
AOI211_X1 g_26_101 (.ZN (n_26_101), .A (n_30_99), .B (n_33_99), .C1 (n_37_97), .C2 (n_38_95) );
AOI211_X1 g_24_102 (.ZN (n_24_102), .A (n_28_100), .B (n_31_100), .C1 (n_35_98), .C2 (n_40_94) );
AOI211_X1 g_22_103 (.ZN (n_22_103), .A (n_26_101), .B (n_29_101), .C1 (n_33_99), .C2 (n_39_96) );
AOI211_X1 g_20_104 (.ZN (n_20_104), .A (n_24_102), .B (n_30_99), .C1 (n_31_100), .C2 (n_37_97) );
AOI211_X1 g_18_105 (.ZN (n_18_105), .A (n_22_103), .B (n_28_100), .C1 (n_29_101), .C2 (n_35_98) );
AOI211_X1 g_17_107 (.ZN (n_17_107), .A (n_20_104), .B (n_26_101), .C1 (n_30_99), .C2 (n_33_99) );
AOI211_X1 g_15_106 (.ZN (n_15_106), .A (n_18_105), .B (n_24_102), .C1 (n_28_100), .C2 (n_31_100) );
AOI211_X1 g_17_105 (.ZN (n_17_105), .A (n_17_107), .B (n_22_103), .C1 (n_26_101), .C2 (n_29_101) );
AOI211_X1 g_19_104 (.ZN (n_19_104), .A (n_15_106), .B (n_20_104), .C1 (n_24_102), .C2 (n_30_99) );
AOI211_X1 g_18_106 (.ZN (n_18_106), .A (n_17_105), .B (n_18_105), .C1 (n_22_103), .C2 (n_28_100) );
AOI211_X1 g_20_105 (.ZN (n_20_105), .A (n_19_104), .B (n_17_107), .C1 (n_20_104), .C2 (n_26_101) );
AOI211_X1 g_22_104 (.ZN (n_22_104), .A (n_18_106), .B (n_15_106), .C1 (n_18_105), .C2 (n_24_102) );
AOI211_X1 g_24_103 (.ZN (n_24_103), .A (n_20_105), .B (n_17_105), .C1 (n_17_107), .C2 (n_22_103) );
AOI211_X1 g_26_102 (.ZN (n_26_102), .A (n_22_104), .B (n_19_104), .C1 (n_15_106), .C2 (n_20_104) );
AOI211_X1 g_28_101 (.ZN (n_28_101), .A (n_24_103), .B (n_18_106), .C1 (n_17_105), .C2 (n_18_105) );
AOI211_X1 g_30_100 (.ZN (n_30_100), .A (n_26_102), .B (n_20_105), .C1 (n_19_104), .C2 (n_17_107) );
AOI211_X1 g_29_102 (.ZN (n_29_102), .A (n_28_101), .B (n_22_104), .C1 (n_18_106), .C2 (n_15_106) );
AOI211_X1 g_31_101 (.ZN (n_31_101), .A (n_30_100), .B (n_24_103), .C1 (n_20_105), .C2 (n_17_105) );
AOI211_X1 g_30_103 (.ZN (n_30_103), .A (n_29_102), .B (n_26_102), .C1 (n_22_104), .C2 (n_19_104) );
AOI211_X1 g_28_102 (.ZN (n_28_102), .A (n_31_101), .B (n_28_101), .C1 (n_24_103), .C2 (n_18_106) );
AOI211_X1 g_30_101 (.ZN (n_30_101), .A (n_30_103), .B (n_30_100), .C1 (n_26_102), .C2 (n_20_105) );
AOI211_X1 g_32_100 (.ZN (n_32_100), .A (n_28_102), .B (n_29_102), .C1 (n_28_101), .C2 (n_22_104) );
AOI211_X1 g_34_99 (.ZN (n_34_99), .A (n_30_101), .B (n_31_101), .C1 (n_30_100), .C2 (n_24_103) );
AOI211_X1 g_36_98 (.ZN (n_36_98), .A (n_32_100), .B (n_30_103), .C1 (n_29_102), .C2 (n_26_102) );
AOI211_X1 g_38_97 (.ZN (n_38_97), .A (n_34_99), .B (n_28_102), .C1 (n_31_101), .C2 (n_28_101) );
AOI211_X1 g_40_96 (.ZN (n_40_96), .A (n_36_98), .B (n_30_101), .C1 (n_30_103), .C2 (n_30_100) );
AOI211_X1 g_42_95 (.ZN (n_42_95), .A (n_38_97), .B (n_32_100), .C1 (n_28_102), .C2 (n_29_102) );
AOI211_X1 g_44_94 (.ZN (n_44_94), .A (n_40_96), .B (n_34_99), .C1 (n_30_101), .C2 (n_31_101) );
AOI211_X1 g_43_96 (.ZN (n_43_96), .A (n_42_95), .B (n_36_98), .C1 (n_32_100), .C2 (n_30_103) );
AOI211_X1 g_45_95 (.ZN (n_45_95), .A (n_44_94), .B (n_38_97), .C1 (n_34_99), .C2 (n_28_102) );
AOI211_X1 g_47_94 (.ZN (n_47_94), .A (n_43_96), .B (n_40_96), .C1 (n_36_98), .C2 (n_30_101) );
AOI211_X1 g_49_93 (.ZN (n_49_93), .A (n_45_95), .B (n_42_95), .C1 (n_38_97), .C2 (n_32_100) );
AOI211_X1 g_51_92 (.ZN (n_51_92), .A (n_47_94), .B (n_44_94), .C1 (n_40_96), .C2 (n_34_99) );
AOI211_X1 g_53_91 (.ZN (n_53_91), .A (n_49_93), .B (n_43_96), .C1 (n_42_95), .C2 (n_36_98) );
AOI211_X1 g_55_90 (.ZN (n_55_90), .A (n_51_92), .B (n_45_95), .C1 (n_44_94), .C2 (n_38_97) );
AOI211_X1 g_54_92 (.ZN (n_54_92), .A (n_53_91), .B (n_47_94), .C1 (n_43_96), .C2 (n_40_96) );
AOI211_X1 g_52_91 (.ZN (n_52_91), .A (n_55_90), .B (n_49_93), .C1 (n_45_95), .C2 (n_42_95) );
AOI211_X1 g_54_90 (.ZN (n_54_90), .A (n_54_92), .B (n_51_92), .C1 (n_47_94), .C2 (n_44_94) );
AOI211_X1 g_56_89 (.ZN (n_56_89), .A (n_52_91), .B (n_53_91), .C1 (n_49_93), .C2 (n_43_96) );
AOI211_X1 g_55_91 (.ZN (n_55_91), .A (n_54_90), .B (n_55_90), .C1 (n_51_92), .C2 (n_45_95) );
AOI211_X1 g_57_90 (.ZN (n_57_90), .A (n_56_89), .B (n_54_92), .C1 (n_53_91), .C2 (n_47_94) );
AOI211_X1 g_59_89 (.ZN (n_59_89), .A (n_55_91), .B (n_52_91), .C1 (n_55_90), .C2 (n_49_93) );
AOI211_X1 g_61_88 (.ZN (n_61_88), .A (n_57_90), .B (n_54_90), .C1 (n_54_92), .C2 (n_51_92) );
AOI211_X1 g_62_86 (.ZN (n_62_86), .A (n_59_89), .B (n_56_89), .C1 (n_52_91), .C2 (n_53_91) );
AOI211_X1 g_64_85 (.ZN (n_64_85), .A (n_61_88), .B (n_55_91), .C1 (n_54_90), .C2 (n_55_90) );
AOI211_X1 g_66_84 (.ZN (n_66_84), .A (n_62_86), .B (n_57_90), .C1 (n_56_89), .C2 (n_54_92) );
AOI211_X1 g_68_83 (.ZN (n_68_83), .A (n_64_85), .B (n_59_89), .C1 (n_55_91), .C2 (n_52_91) );
AOI211_X1 g_70_82 (.ZN (n_70_82), .A (n_66_84), .B (n_61_88), .C1 (n_57_90), .C2 (n_54_90) );
AOI211_X1 g_72_81 (.ZN (n_72_81), .A (n_68_83), .B (n_62_86), .C1 (n_59_89), .C2 (n_56_89) );
AOI211_X1 g_74_80 (.ZN (n_74_80), .A (n_70_82), .B (n_64_85), .C1 (n_61_88), .C2 (n_55_91) );
AOI211_X1 g_76_79 (.ZN (n_76_79), .A (n_72_81), .B (n_66_84), .C1 (n_62_86), .C2 (n_57_90) );
AOI211_X1 g_78_78 (.ZN (n_78_78), .A (n_74_80), .B (n_68_83), .C1 (n_64_85), .C2 (n_59_89) );
AOI211_X1 g_80_77 (.ZN (n_80_77), .A (n_76_79), .B (n_70_82), .C1 (n_66_84), .C2 (n_61_88) );
AOI211_X1 g_82_78 (.ZN (n_82_78), .A (n_78_78), .B (n_72_81), .C1 (n_68_83), .C2 (n_62_86) );
AOI211_X1 g_80_79 (.ZN (n_80_79), .A (n_80_77), .B (n_74_80), .C1 (n_70_82), .C2 (n_64_85) );
AOI211_X1 g_78_80 (.ZN (n_78_80), .A (n_82_78), .B (n_76_79), .C1 (n_72_81), .C2 (n_66_84) );
AOI211_X1 g_76_81 (.ZN (n_76_81), .A (n_80_79), .B (n_78_78), .C1 (n_74_80), .C2 (n_68_83) );
AOI211_X1 g_74_82 (.ZN (n_74_82), .A (n_78_80), .B (n_80_77), .C1 (n_76_79), .C2 (n_70_82) );
AOI211_X1 g_72_83 (.ZN (n_72_83), .A (n_76_81), .B (n_82_78), .C1 (n_78_78), .C2 (n_72_81) );
AOI211_X1 g_70_84 (.ZN (n_70_84), .A (n_74_82), .B (n_80_79), .C1 (n_80_77), .C2 (n_74_80) );
AOI211_X1 g_68_85 (.ZN (n_68_85), .A (n_72_83), .B (n_78_80), .C1 (n_82_78), .C2 (n_76_79) );
AOI211_X1 g_66_86 (.ZN (n_66_86), .A (n_70_84), .B (n_76_81), .C1 (n_80_79), .C2 (n_78_78) );
AOI211_X1 g_64_87 (.ZN (n_64_87), .A (n_68_85), .B (n_74_82), .C1 (n_78_80), .C2 (n_80_77) );
AOI211_X1 g_62_88 (.ZN (n_62_88), .A (n_66_86), .B (n_72_83), .C1 (n_76_81), .C2 (n_82_78) );
AOI211_X1 g_60_89 (.ZN (n_60_89), .A (n_64_87), .B (n_70_84), .C1 (n_74_82), .C2 (n_80_79) );
AOI211_X1 g_58_90 (.ZN (n_58_90), .A (n_62_88), .B (n_68_85), .C1 (n_72_83), .C2 (n_78_80) );
AOI211_X1 g_56_91 (.ZN (n_56_91), .A (n_60_89), .B (n_66_86), .C1 (n_70_84), .C2 (n_76_81) );
AOI211_X1 g_58_92 (.ZN (n_58_92), .A (n_58_90), .B (n_64_87), .C1 (n_68_85), .C2 (n_74_82) );
AOI211_X1 g_60_91 (.ZN (n_60_91), .A (n_56_91), .B (n_62_88), .C1 (n_66_86), .C2 (n_72_83) );
AOI211_X1 g_62_90 (.ZN (n_62_90), .A (n_58_92), .B (n_60_89), .C1 (n_64_87), .C2 (n_70_84) );
AOI211_X1 g_63_88 (.ZN (n_63_88), .A (n_60_91), .B (n_58_90), .C1 (n_62_88), .C2 (n_68_85) );
AOI211_X1 g_64_86 (.ZN (n_64_86), .A (n_62_90), .B (n_56_91), .C1 (n_60_89), .C2 (n_66_86) );
AOI211_X1 g_66_85 (.ZN (n_66_85), .A (n_63_88), .B (n_58_92), .C1 (n_58_90), .C2 (n_64_87) );
AOI211_X1 g_68_84 (.ZN (n_68_84), .A (n_64_86), .B (n_60_91), .C1 (n_56_91), .C2 (n_62_88) );
AOI211_X1 g_70_83 (.ZN (n_70_83), .A (n_66_85), .B (n_62_90), .C1 (n_58_92), .C2 (n_60_89) );
AOI211_X1 g_72_82 (.ZN (n_72_82), .A (n_68_84), .B (n_63_88), .C1 (n_60_91), .C2 (n_58_90) );
AOI211_X1 g_74_81 (.ZN (n_74_81), .A (n_70_83), .B (n_64_86), .C1 (n_62_90), .C2 (n_56_91) );
AOI211_X1 g_76_80 (.ZN (n_76_80), .A (n_72_82), .B (n_66_85), .C1 (n_63_88), .C2 (n_58_92) );
AOI211_X1 g_78_79 (.ZN (n_78_79), .A (n_74_81), .B (n_68_84), .C1 (n_64_86), .C2 (n_60_91) );
AOI211_X1 g_80_78 (.ZN (n_80_78), .A (n_76_80), .B (n_70_83), .C1 (n_66_85), .C2 (n_62_90) );
AOI211_X1 g_82_77 (.ZN (n_82_77), .A (n_78_79), .B (n_72_82), .C1 (n_68_84), .C2 (n_63_88) );
AOI211_X1 g_84_76 (.ZN (n_84_76), .A (n_80_78), .B (n_74_81), .C1 (n_70_83), .C2 (n_64_86) );
AOI211_X1 g_83_78 (.ZN (n_83_78), .A (n_82_77), .B (n_76_80), .C1 (n_72_82), .C2 (n_66_85) );
AOI211_X1 g_85_77 (.ZN (n_85_77), .A (n_84_76), .B (n_78_79), .C1 (n_74_81), .C2 (n_68_84) );
AOI211_X1 g_87_76 (.ZN (n_87_76), .A (n_83_78), .B (n_80_78), .C1 (n_76_80), .C2 (n_70_83) );
AOI211_X1 g_89_75 (.ZN (n_89_75), .A (n_85_77), .B (n_82_77), .C1 (n_78_79), .C2 (n_72_82) );
AOI211_X1 g_91_74 (.ZN (n_91_74), .A (n_87_76), .B (n_84_76), .C1 (n_80_78), .C2 (n_74_81) );
AOI211_X1 g_93_73 (.ZN (n_93_73), .A (n_89_75), .B (n_83_78), .C1 (n_82_77), .C2 (n_76_80) );
AOI211_X1 g_95_72 (.ZN (n_95_72), .A (n_91_74), .B (n_85_77), .C1 (n_84_76), .C2 (n_78_79) );
AOI211_X1 g_97_71 (.ZN (n_97_71), .A (n_93_73), .B (n_87_76), .C1 (n_83_78), .C2 (n_80_78) );
AOI211_X1 g_99_70 (.ZN (n_99_70), .A (n_95_72), .B (n_89_75), .C1 (n_85_77), .C2 (n_82_77) );
AOI211_X1 g_101_69 (.ZN (n_101_69), .A (n_97_71), .B (n_91_74), .C1 (n_87_76), .C2 (n_84_76) );
AOI211_X1 g_103_68 (.ZN (n_103_68), .A (n_99_70), .B (n_93_73), .C1 (n_89_75), .C2 (n_83_78) );
AOI211_X1 g_105_67 (.ZN (n_105_67), .A (n_101_69), .B (n_95_72), .C1 (n_91_74), .C2 (n_85_77) );
AOI211_X1 g_107_66 (.ZN (n_107_66), .A (n_103_68), .B (n_97_71), .C1 (n_93_73), .C2 (n_87_76) );
AOI211_X1 g_109_65 (.ZN (n_109_65), .A (n_105_67), .B (n_99_70), .C1 (n_95_72), .C2 (n_89_75) );
AOI211_X1 g_108_67 (.ZN (n_108_67), .A (n_107_66), .B (n_101_69), .C1 (n_97_71), .C2 (n_91_74) );
AOI211_X1 g_110_66 (.ZN (n_110_66), .A (n_109_65), .B (n_103_68), .C1 (n_99_70), .C2 (n_93_73) );
AOI211_X1 g_112_65 (.ZN (n_112_65), .A (n_108_67), .B (n_105_67), .C1 (n_101_69), .C2 (n_95_72) );
AOI211_X1 g_114_64 (.ZN (n_114_64), .A (n_110_66), .B (n_107_66), .C1 (n_103_68), .C2 (n_97_71) );
AOI211_X1 g_116_63 (.ZN (n_116_63), .A (n_112_65), .B (n_109_65), .C1 (n_105_67), .C2 (n_99_70) );
AOI211_X1 g_118_62 (.ZN (n_118_62), .A (n_114_64), .B (n_108_67), .C1 (n_107_66), .C2 (n_101_69) );
AOI211_X1 g_120_61 (.ZN (n_120_61), .A (n_116_63), .B (n_110_66), .C1 (n_109_65), .C2 (n_103_68) );
AOI211_X1 g_122_60 (.ZN (n_122_60), .A (n_118_62), .B (n_112_65), .C1 (n_108_67), .C2 (n_105_67) );
AOI211_X1 g_124_59 (.ZN (n_124_59), .A (n_120_61), .B (n_114_64), .C1 (n_110_66), .C2 (n_107_66) );
AOI211_X1 g_126_58 (.ZN (n_126_58), .A (n_122_60), .B (n_116_63), .C1 (n_112_65), .C2 (n_109_65) );
AOI211_X1 g_128_57 (.ZN (n_128_57), .A (n_124_59), .B (n_118_62), .C1 (n_114_64), .C2 (n_108_67) );
AOI211_X1 g_130_56 (.ZN (n_130_56), .A (n_126_58), .B (n_120_61), .C1 (n_116_63), .C2 (n_110_66) );
AOI211_X1 g_129_58 (.ZN (n_129_58), .A (n_128_57), .B (n_122_60), .C1 (n_118_62), .C2 (n_112_65) );
AOI211_X1 g_127_57 (.ZN (n_127_57), .A (n_130_56), .B (n_124_59), .C1 (n_120_61), .C2 (n_114_64) );
AOI211_X1 g_129_56 (.ZN (n_129_56), .A (n_129_58), .B (n_126_58), .C1 (n_122_60), .C2 (n_116_63) );
AOI211_X1 g_131_55 (.ZN (n_131_55), .A (n_127_57), .B (n_128_57), .C1 (n_124_59), .C2 (n_118_62) );
AOI211_X1 g_133_54 (.ZN (n_133_54), .A (n_129_56), .B (n_130_56), .C1 (n_126_58), .C2 (n_120_61) );
AOI211_X1 g_135_53 (.ZN (n_135_53), .A (n_131_55), .B (n_129_58), .C1 (n_128_57), .C2 (n_122_60) );
AOI211_X1 g_137_52 (.ZN (n_137_52), .A (n_133_54), .B (n_127_57), .C1 (n_130_56), .C2 (n_124_59) );
AOI211_X1 g_139_51 (.ZN (n_139_51), .A (n_135_53), .B (n_129_56), .C1 (n_129_58), .C2 (n_126_58) );
AOI211_X1 g_141_50 (.ZN (n_141_50), .A (n_137_52), .B (n_131_55), .C1 (n_127_57), .C2 (n_128_57) );
AOI211_X1 g_143_49 (.ZN (n_143_49), .A (n_139_51), .B (n_133_54), .C1 (n_129_56), .C2 (n_130_56) );
AOI211_X1 g_145_48 (.ZN (n_145_48), .A (n_141_50), .B (n_135_53), .C1 (n_131_55), .C2 (n_129_58) );
AOI211_X1 g_147_49 (.ZN (n_147_49), .A (n_143_49), .B (n_137_52), .C1 (n_133_54), .C2 (n_127_57) );
AOI211_X1 g_145_50 (.ZN (n_145_50), .A (n_145_48), .B (n_139_51), .C1 (n_135_53), .C2 (n_129_56) );
AOI211_X1 g_143_51 (.ZN (n_143_51), .A (n_147_49), .B (n_141_50), .C1 (n_137_52), .C2 (n_131_55) );
AOI211_X1 g_141_52 (.ZN (n_141_52), .A (n_145_50), .B (n_143_49), .C1 (n_139_51), .C2 (n_133_54) );
AOI211_X1 g_139_53 (.ZN (n_139_53), .A (n_143_51), .B (n_145_48), .C1 (n_141_50), .C2 (n_135_53) );
AOI211_X1 g_137_54 (.ZN (n_137_54), .A (n_141_52), .B (n_147_49), .C1 (n_143_49), .C2 (n_137_52) );
AOI211_X1 g_135_55 (.ZN (n_135_55), .A (n_139_53), .B (n_145_50), .C1 (n_145_48), .C2 (n_139_51) );
AOI211_X1 g_133_56 (.ZN (n_133_56), .A (n_137_54), .B (n_143_51), .C1 (n_147_49), .C2 (n_141_50) );
AOI211_X1 g_131_57 (.ZN (n_131_57), .A (n_135_55), .B (n_141_52), .C1 (n_145_50), .C2 (n_143_49) );
AOI211_X1 g_130_59 (.ZN (n_130_59), .A (n_133_56), .B (n_139_53), .C1 (n_143_51), .C2 (n_145_48) );
AOI211_X1 g_128_58 (.ZN (n_128_58), .A (n_131_57), .B (n_137_54), .C1 (n_141_52), .C2 (n_147_49) );
AOI211_X1 g_130_57 (.ZN (n_130_57), .A (n_130_59), .B (n_135_55), .C1 (n_139_53), .C2 (n_145_50) );
AOI211_X1 g_132_56 (.ZN (n_132_56), .A (n_128_58), .B (n_133_56), .C1 (n_137_54), .C2 (n_143_51) );
AOI211_X1 g_134_55 (.ZN (n_134_55), .A (n_130_57), .B (n_131_57), .C1 (n_135_55), .C2 (n_141_52) );
AOI211_X1 g_136_54 (.ZN (n_136_54), .A (n_132_56), .B (n_130_59), .C1 (n_133_56), .C2 (n_139_53) );
AOI211_X1 g_138_53 (.ZN (n_138_53), .A (n_134_55), .B (n_128_58), .C1 (n_131_57), .C2 (n_137_54) );
AOI211_X1 g_140_52 (.ZN (n_140_52), .A (n_136_54), .B (n_130_57), .C1 (n_130_59), .C2 (n_135_55) );
AOI211_X1 g_142_51 (.ZN (n_142_51), .A (n_138_53), .B (n_132_56), .C1 (n_128_58), .C2 (n_133_56) );
AOI211_X1 g_144_50 (.ZN (n_144_50), .A (n_140_52), .B (n_134_55), .C1 (n_130_57), .C2 (n_131_57) );
AOI211_X1 g_146_51 (.ZN (n_146_51), .A (n_142_51), .B (n_136_54), .C1 (n_132_56), .C2 (n_130_59) );
AOI211_X1 g_144_52 (.ZN (n_144_52), .A (n_144_50), .B (n_138_53), .C1 (n_134_55), .C2 (n_128_58) );
AOI211_X1 g_142_53 (.ZN (n_142_53), .A (n_146_51), .B (n_140_52), .C1 (n_136_54), .C2 (n_130_57) );
AOI211_X1 g_140_54 (.ZN (n_140_54), .A (n_144_52), .B (n_142_51), .C1 (n_138_53), .C2 (n_132_56) );
AOI211_X1 g_138_55 (.ZN (n_138_55), .A (n_142_53), .B (n_144_50), .C1 (n_140_52), .C2 (n_134_55) );
AOI211_X1 g_136_56 (.ZN (n_136_56), .A (n_140_54), .B (n_146_51), .C1 (n_142_51), .C2 (n_136_54) );
AOI211_X1 g_134_57 (.ZN (n_134_57), .A (n_138_55), .B (n_144_52), .C1 (n_144_50), .C2 (n_138_53) );
AOI211_X1 g_132_58 (.ZN (n_132_58), .A (n_136_56), .B (n_142_53), .C1 (n_146_51), .C2 (n_140_52) );
AOI211_X1 g_131_60 (.ZN (n_131_60), .A (n_134_57), .B (n_140_54), .C1 (n_144_52), .C2 (n_142_51) );
AOI211_X1 g_130_58 (.ZN (n_130_58), .A (n_132_58), .B (n_138_55), .C1 (n_142_53), .C2 (n_144_50) );
AOI211_X1 g_132_57 (.ZN (n_132_57), .A (n_131_60), .B (n_136_56), .C1 (n_140_54), .C2 (n_146_51) );
AOI211_X1 g_134_56 (.ZN (n_134_56), .A (n_130_58), .B (n_134_57), .C1 (n_138_55), .C2 (n_144_52) );
AOI211_X1 g_136_55 (.ZN (n_136_55), .A (n_132_57), .B (n_132_58), .C1 (n_136_56), .C2 (n_142_53) );
AOI211_X1 g_138_54 (.ZN (n_138_54), .A (n_134_56), .B (n_131_60), .C1 (n_134_57), .C2 (n_140_54) );
AOI211_X1 g_140_53 (.ZN (n_140_53), .A (n_136_55), .B (n_130_58), .C1 (n_132_58), .C2 (n_138_55) );
AOI211_X1 g_142_52 (.ZN (n_142_52), .A (n_138_54), .B (n_132_57), .C1 (n_131_60), .C2 (n_136_56) );
AOI211_X1 g_144_51 (.ZN (n_144_51), .A (n_140_53), .B (n_134_56), .C1 (n_130_58), .C2 (n_134_57) );
AOI211_X1 g_146_50 (.ZN (n_146_50), .A (n_142_52), .B (n_136_55), .C1 (n_132_57), .C2 (n_132_58) );
AOI211_X1 g_147_52 (.ZN (n_147_52), .A (n_144_51), .B (n_138_54), .C1 (n_134_56), .C2 (n_131_60) );
AOI211_X1 g_149_53 (.ZN (n_149_53), .A (n_146_50), .B (n_140_53), .C1 (n_136_55), .C2 (n_130_58) );
AOI211_X1 g_148_51 (.ZN (n_148_51), .A (n_147_52), .B (n_142_52), .C1 (n_138_54), .C2 (n_132_57) );
AOI211_X1 g_146_52 (.ZN (n_146_52), .A (n_149_53), .B (n_144_51), .C1 (n_140_53), .C2 (n_134_56) );
AOI211_X1 g_147_54 (.ZN (n_147_54), .A (n_148_51), .B (n_146_50), .C1 (n_142_52), .C2 (n_136_55) );
AOI211_X1 g_145_53 (.ZN (n_145_53), .A (n_146_52), .B (n_147_52), .C1 (n_144_51), .C2 (n_138_54) );
AOI211_X1 g_143_52 (.ZN (n_143_52), .A (n_147_54), .B (n_149_53), .C1 (n_146_50), .C2 (n_140_53) );
AOI211_X1 g_141_53 (.ZN (n_141_53), .A (n_145_53), .B (n_148_51), .C1 (n_147_52), .C2 (n_142_52) );
AOI211_X1 g_139_54 (.ZN (n_139_54), .A (n_143_52), .B (n_146_52), .C1 (n_149_53), .C2 (n_144_51) );
AOI211_X1 g_137_55 (.ZN (n_137_55), .A (n_141_53), .B (n_147_54), .C1 (n_148_51), .C2 (n_146_50) );
AOI211_X1 g_135_56 (.ZN (n_135_56), .A (n_139_54), .B (n_145_53), .C1 (n_146_52), .C2 (n_147_52) );
AOI211_X1 g_133_57 (.ZN (n_133_57), .A (n_137_55), .B (n_143_52), .C1 (n_147_54), .C2 (n_149_53) );
AOI211_X1 g_131_58 (.ZN (n_131_58), .A (n_135_56), .B (n_141_53), .C1 (n_145_53), .C2 (n_148_51) );
AOI211_X1 g_129_59 (.ZN (n_129_59), .A (n_133_57), .B (n_139_54), .C1 (n_143_52), .C2 (n_146_52) );
AOI211_X1 g_127_60 (.ZN (n_127_60), .A (n_131_58), .B (n_137_55), .C1 (n_141_53), .C2 (n_147_54) );
AOI211_X1 g_125_61 (.ZN (n_125_61), .A (n_129_59), .B (n_135_56), .C1 (n_139_54), .C2 (n_145_53) );
AOI211_X1 g_126_59 (.ZN (n_126_59), .A (n_127_60), .B (n_133_57), .C1 (n_137_55), .C2 (n_143_52) );
AOI211_X1 g_128_60 (.ZN (n_128_60), .A (n_125_61), .B (n_131_58), .C1 (n_135_56), .C2 (n_141_53) );
AOI211_X1 g_126_61 (.ZN (n_126_61), .A (n_126_59), .B (n_129_59), .C1 (n_133_57), .C2 (n_139_54) );
AOI211_X1 g_127_59 (.ZN (n_127_59), .A (n_128_60), .B (n_127_60), .C1 (n_131_58), .C2 (n_137_55) );
AOI211_X1 g_125_58 (.ZN (n_125_58), .A (n_126_61), .B (n_125_61), .C1 (n_129_59), .C2 (n_135_56) );
AOI211_X1 g_124_60 (.ZN (n_124_60), .A (n_127_59), .B (n_126_59), .C1 (n_127_60), .C2 (n_133_57) );
AOI211_X1 g_123_62 (.ZN (n_123_62), .A (n_125_58), .B (n_128_60), .C1 (n_125_61), .C2 (n_131_58) );
AOI211_X1 g_121_63 (.ZN (n_121_63), .A (n_124_60), .B (n_126_61), .C1 (n_126_59), .C2 (n_129_59) );
AOI211_X1 g_122_61 (.ZN (n_122_61), .A (n_123_62), .B (n_127_59), .C1 (n_128_60), .C2 (n_127_60) );
AOI211_X1 g_123_59 (.ZN (n_123_59), .A (n_121_63), .B (n_125_58), .C1 (n_126_61), .C2 (n_125_61) );
AOI211_X1 g_121_60 (.ZN (n_121_60), .A (n_122_61), .B (n_124_60), .C1 (n_127_59), .C2 (n_126_59) );
AOI211_X1 g_119_61 (.ZN (n_119_61), .A (n_123_59), .B (n_123_62), .C1 (n_125_58), .C2 (n_128_60) );
AOI211_X1 g_117_62 (.ZN (n_117_62), .A (n_121_60), .B (n_121_63), .C1 (n_124_60), .C2 (n_126_61) );
AOI211_X1 g_115_63 (.ZN (n_115_63), .A (n_119_61), .B (n_122_61), .C1 (n_123_62), .C2 (n_127_59) );
AOI211_X1 g_113_64 (.ZN (n_113_64), .A (n_117_62), .B (n_123_59), .C1 (n_121_63), .C2 (n_125_58) );
AOI211_X1 g_111_65 (.ZN (n_111_65), .A (n_115_63), .B (n_121_60), .C1 (n_122_61), .C2 (n_124_60) );
AOI211_X1 g_109_66 (.ZN (n_109_66), .A (n_113_64), .B (n_119_61), .C1 (n_123_59), .C2 (n_123_62) );
AOI211_X1 g_107_67 (.ZN (n_107_67), .A (n_111_65), .B (n_117_62), .C1 (n_121_60), .C2 (n_121_63) );
AOI211_X1 g_105_68 (.ZN (n_105_68), .A (n_109_66), .B (n_115_63), .C1 (n_119_61), .C2 (n_122_61) );
AOI211_X1 g_103_69 (.ZN (n_103_69), .A (n_107_67), .B (n_113_64), .C1 (n_117_62), .C2 (n_123_59) );
AOI211_X1 g_101_70 (.ZN (n_101_70), .A (n_105_68), .B (n_111_65), .C1 (n_115_63), .C2 (n_121_60) );
AOI211_X1 g_99_71 (.ZN (n_99_71), .A (n_103_69), .B (n_109_66), .C1 (n_113_64), .C2 (n_119_61) );
AOI211_X1 g_97_72 (.ZN (n_97_72), .A (n_101_70), .B (n_107_67), .C1 (n_111_65), .C2 (n_117_62) );
AOI211_X1 g_95_71 (.ZN (n_95_71), .A (n_99_71), .B (n_105_68), .C1 (n_109_66), .C2 (n_115_63) );
AOI211_X1 g_93_72 (.ZN (n_93_72), .A (n_97_72), .B (n_103_69), .C1 (n_107_67), .C2 (n_113_64) );
AOI211_X1 g_91_73 (.ZN (n_91_73), .A (n_95_71), .B (n_101_70), .C1 (n_105_68), .C2 (n_111_65) );
AOI211_X1 g_89_74 (.ZN (n_89_74), .A (n_93_72), .B (n_99_71), .C1 (n_103_69), .C2 (n_109_66) );
AOI211_X1 g_88_76 (.ZN (n_88_76), .A (n_91_73), .B (n_97_72), .C1 (n_101_70), .C2 (n_107_67) );
AOI211_X1 g_90_75 (.ZN (n_90_75), .A (n_89_74), .B (n_95_71), .C1 (n_99_71), .C2 (n_105_68) );
AOI211_X1 g_92_74 (.ZN (n_92_74), .A (n_88_76), .B (n_93_72), .C1 (n_97_72), .C2 (n_103_69) );
AOI211_X1 g_94_73 (.ZN (n_94_73), .A (n_90_75), .B (n_91_73), .C1 (n_95_71), .C2 (n_101_70) );
AOI211_X1 g_93_75 (.ZN (n_93_75), .A (n_92_74), .B (n_89_74), .C1 (n_93_72), .C2 (n_99_71) );
AOI211_X1 g_95_74 (.ZN (n_95_74), .A (n_94_73), .B (n_88_76), .C1 (n_91_73), .C2 (n_97_72) );
AOI211_X1 g_97_73 (.ZN (n_97_73), .A (n_93_75), .B (n_90_75), .C1 (n_89_74), .C2 (n_95_71) );
AOI211_X1 g_99_72 (.ZN (n_99_72), .A (n_95_74), .B (n_92_74), .C1 (n_88_76), .C2 (n_93_72) );
AOI211_X1 g_101_71 (.ZN (n_101_71), .A (n_97_73), .B (n_94_73), .C1 (n_90_75), .C2 (n_91_73) );
AOI211_X1 g_103_70 (.ZN (n_103_70), .A (n_99_72), .B (n_93_75), .C1 (n_92_74), .C2 (n_89_74) );
AOI211_X1 g_105_69 (.ZN (n_105_69), .A (n_101_71), .B (n_95_74), .C1 (n_94_73), .C2 (n_88_76) );
AOI211_X1 g_107_68 (.ZN (n_107_68), .A (n_103_70), .B (n_97_73), .C1 (n_93_75), .C2 (n_90_75) );
AOI211_X1 g_109_67 (.ZN (n_109_67), .A (n_105_69), .B (n_99_72), .C1 (n_95_74), .C2 (n_92_74) );
AOI211_X1 g_108_69 (.ZN (n_108_69), .A (n_107_68), .B (n_101_71), .C1 (n_97_73), .C2 (n_94_73) );
AOI211_X1 g_106_68 (.ZN (n_106_68), .A (n_109_67), .B (n_103_70), .C1 (n_99_72), .C2 (n_93_75) );
AOI211_X1 g_104_69 (.ZN (n_104_69), .A (n_108_69), .B (n_105_69), .C1 (n_101_71), .C2 (n_95_74) );
AOI211_X1 g_102_70 (.ZN (n_102_70), .A (n_106_68), .B (n_107_68), .C1 (n_103_70), .C2 (n_97_73) );
AOI211_X1 g_100_71 (.ZN (n_100_71), .A (n_104_69), .B (n_109_67), .C1 (n_105_69), .C2 (n_99_72) );
AOI211_X1 g_98_72 (.ZN (n_98_72), .A (n_102_70), .B (n_108_69), .C1 (n_107_68), .C2 (n_101_71) );
AOI211_X1 g_96_73 (.ZN (n_96_73), .A (n_100_71), .B (n_106_68), .C1 (n_109_67), .C2 (n_103_70) );
AOI211_X1 g_94_74 (.ZN (n_94_74), .A (n_98_72), .B (n_104_69), .C1 (n_108_69), .C2 (n_105_69) );
AOI211_X1 g_92_75 (.ZN (n_92_75), .A (n_96_73), .B (n_102_70), .C1 (n_106_68), .C2 (n_107_68) );
AOI211_X1 g_90_76 (.ZN (n_90_76), .A (n_94_74), .B (n_100_71), .C1 (n_104_69), .C2 (n_109_67) );
AOI211_X1 g_88_77 (.ZN (n_88_77), .A (n_92_75), .B (n_98_72), .C1 (n_102_70), .C2 (n_108_69) );
AOI211_X1 g_86_78 (.ZN (n_86_78), .A (n_90_76), .B (n_96_73), .C1 (n_100_71), .C2 (n_106_68) );
AOI211_X1 g_85_76 (.ZN (n_85_76), .A (n_88_77), .B (n_94_74), .C1 (n_98_72), .C2 (n_104_69) );
AOI211_X1 g_83_77 (.ZN (n_83_77), .A (n_86_78), .B (n_92_75), .C1 (n_96_73), .C2 (n_102_70) );
AOI211_X1 g_81_78 (.ZN (n_81_78), .A (n_85_76), .B (n_90_76), .C1 (n_94_74), .C2 (n_100_71) );
AOI211_X1 g_79_79 (.ZN (n_79_79), .A (n_83_77), .B (n_88_77), .C1 (n_92_75), .C2 (n_98_72) );
AOI211_X1 g_77_80 (.ZN (n_77_80), .A (n_81_78), .B (n_86_78), .C1 (n_90_76), .C2 (n_96_73) );
AOI211_X1 g_75_81 (.ZN (n_75_81), .A (n_79_79), .B (n_85_76), .C1 (n_88_77), .C2 (n_94_74) );
AOI211_X1 g_73_82 (.ZN (n_73_82), .A (n_77_80), .B (n_83_77), .C1 (n_86_78), .C2 (n_92_75) );
AOI211_X1 g_71_83 (.ZN (n_71_83), .A (n_75_81), .B (n_81_78), .C1 (n_85_76), .C2 (n_90_76) );
AOI211_X1 g_69_84 (.ZN (n_69_84), .A (n_73_82), .B (n_79_79), .C1 (n_83_77), .C2 (n_88_77) );
AOI211_X1 g_67_85 (.ZN (n_67_85), .A (n_71_83), .B (n_77_80), .C1 (n_81_78), .C2 (n_86_78) );
AOI211_X1 g_65_86 (.ZN (n_65_86), .A (n_69_84), .B (n_75_81), .C1 (n_79_79), .C2 (n_85_76) );
AOI211_X1 g_63_87 (.ZN (n_63_87), .A (n_67_85), .B (n_73_82), .C1 (n_77_80), .C2 (n_83_77) );
AOI211_X1 g_64_89 (.ZN (n_64_89), .A (n_65_86), .B (n_71_83), .C1 (n_75_81), .C2 (n_81_78) );
AOI211_X1 g_65_87 (.ZN (n_65_87), .A (n_63_87), .B (n_69_84), .C1 (n_73_82), .C2 (n_79_79) );
AOI211_X1 g_67_86 (.ZN (n_67_86), .A (n_64_89), .B (n_67_85), .C1 (n_71_83), .C2 (n_77_80) );
AOI211_X1 g_69_85 (.ZN (n_69_85), .A (n_65_87), .B (n_65_86), .C1 (n_69_84), .C2 (n_75_81) );
AOI211_X1 g_71_84 (.ZN (n_71_84), .A (n_67_86), .B (n_63_87), .C1 (n_67_85), .C2 (n_73_82) );
AOI211_X1 g_73_83 (.ZN (n_73_83), .A (n_69_85), .B (n_64_89), .C1 (n_65_86), .C2 (n_71_83) );
AOI211_X1 g_75_82 (.ZN (n_75_82), .A (n_71_84), .B (n_65_87), .C1 (n_63_87), .C2 (n_69_84) );
AOI211_X1 g_77_81 (.ZN (n_77_81), .A (n_73_83), .B (n_67_86), .C1 (n_64_89), .C2 (n_67_85) );
AOI211_X1 g_79_80 (.ZN (n_79_80), .A (n_75_82), .B (n_69_85), .C1 (n_65_87), .C2 (n_65_86) );
AOI211_X1 g_81_79 (.ZN (n_81_79), .A (n_77_81), .B (n_71_84), .C1 (n_67_86), .C2 (n_63_87) );
AOI211_X1 g_80_81 (.ZN (n_80_81), .A (n_79_80), .B (n_73_83), .C1 (n_69_85), .C2 (n_64_89) );
AOI211_X1 g_82_80 (.ZN (n_82_80), .A (n_81_79), .B (n_75_82), .C1 (n_71_84), .C2 (n_65_87) );
AOI211_X1 g_84_79 (.ZN (n_84_79), .A (n_80_81), .B (n_77_81), .C1 (n_73_83), .C2 (n_67_86) );
AOI211_X1 g_83_81 (.ZN (n_83_81), .A (n_82_80), .B (n_79_80), .C1 (n_75_82), .C2 (n_69_85) );
AOI211_X1 g_82_79 (.ZN (n_82_79), .A (n_84_79), .B (n_81_79), .C1 (n_77_81), .C2 (n_71_84) );
AOI211_X1 g_84_78 (.ZN (n_84_78), .A (n_83_81), .B (n_80_81), .C1 (n_79_80), .C2 (n_73_83) );
AOI211_X1 g_86_77 (.ZN (n_86_77), .A (n_82_79), .B (n_82_80), .C1 (n_81_79), .C2 (n_75_82) );
AOI211_X1 g_85_79 (.ZN (n_85_79), .A (n_84_78), .B (n_84_79), .C1 (n_80_81), .C2 (n_77_81) );
AOI211_X1 g_87_78 (.ZN (n_87_78), .A (n_86_77), .B (n_83_81), .C1 (n_82_80), .C2 (n_79_80) );
AOI211_X1 g_89_77 (.ZN (n_89_77), .A (n_85_79), .B (n_82_79), .C1 (n_84_79), .C2 (n_81_79) );
AOI211_X1 g_91_76 (.ZN (n_91_76), .A (n_87_78), .B (n_84_78), .C1 (n_83_81), .C2 (n_80_81) );
AOI211_X1 g_90_78 (.ZN (n_90_78), .A (n_89_77), .B (n_86_77), .C1 (n_82_79), .C2 (n_82_80) );
AOI211_X1 g_89_76 (.ZN (n_89_76), .A (n_91_76), .B (n_85_79), .C1 (n_84_78), .C2 (n_84_79) );
AOI211_X1 g_91_75 (.ZN (n_91_75), .A (n_90_78), .B (n_87_78), .C1 (n_86_77), .C2 (n_83_81) );
AOI211_X1 g_93_74 (.ZN (n_93_74), .A (n_89_76), .B (n_89_77), .C1 (n_85_79), .C2 (n_82_79) );
AOI211_X1 g_95_73 (.ZN (n_95_73), .A (n_91_75), .B (n_91_76), .C1 (n_87_78), .C2 (n_84_78) );
AOI211_X1 g_94_75 (.ZN (n_94_75), .A (n_93_74), .B (n_90_78), .C1 (n_89_77), .C2 (n_86_77) );
AOI211_X1 g_96_74 (.ZN (n_96_74), .A (n_95_73), .B (n_89_76), .C1 (n_91_76), .C2 (n_85_79) );
AOI211_X1 g_98_73 (.ZN (n_98_73), .A (n_94_75), .B (n_91_75), .C1 (n_90_78), .C2 (n_87_78) );
AOI211_X1 g_100_72 (.ZN (n_100_72), .A (n_96_74), .B (n_93_74), .C1 (n_89_76), .C2 (n_89_77) );
AOI211_X1 g_102_71 (.ZN (n_102_71), .A (n_98_73), .B (n_95_73), .C1 (n_91_75), .C2 (n_91_76) );
AOI211_X1 g_104_70 (.ZN (n_104_70), .A (n_100_72), .B (n_94_75), .C1 (n_93_74), .C2 (n_90_78) );
AOI211_X1 g_106_69 (.ZN (n_106_69), .A (n_102_71), .B (n_96_74), .C1 (n_95_73), .C2 (n_89_76) );
AOI211_X1 g_108_68 (.ZN (n_108_68), .A (n_104_70), .B (n_98_73), .C1 (n_94_75), .C2 (n_91_75) );
AOI211_X1 g_110_67 (.ZN (n_110_67), .A (n_106_69), .B (n_100_72), .C1 (n_96_74), .C2 (n_93_74) );
AOI211_X1 g_112_66 (.ZN (n_112_66), .A (n_108_68), .B (n_102_71), .C1 (n_98_73), .C2 (n_95_73) );
AOI211_X1 g_114_65 (.ZN (n_114_65), .A (n_110_67), .B (n_104_70), .C1 (n_100_72), .C2 (n_94_75) );
AOI211_X1 g_116_64 (.ZN (n_116_64), .A (n_112_66), .B (n_106_69), .C1 (n_102_71), .C2 (n_96_74) );
AOI211_X1 g_118_63 (.ZN (n_118_63), .A (n_114_65), .B (n_108_68), .C1 (n_104_70), .C2 (n_98_73) );
AOI211_X1 g_120_62 (.ZN (n_120_62), .A (n_116_64), .B (n_110_67), .C1 (n_106_69), .C2 (n_100_72) );
AOI211_X1 g_119_64 (.ZN (n_119_64), .A (n_118_63), .B (n_112_66), .C1 (n_108_68), .C2 (n_102_71) );
AOI211_X1 g_117_65 (.ZN (n_117_65), .A (n_120_62), .B (n_114_65), .C1 (n_110_67), .C2 (n_104_70) );
AOI211_X1 g_115_66 (.ZN (n_115_66), .A (n_119_64), .B (n_116_64), .C1 (n_112_66), .C2 (n_106_69) );
AOI211_X1 g_113_67 (.ZN (n_113_67), .A (n_117_65), .B (n_118_63), .C1 (n_114_65), .C2 (n_108_68) );
AOI211_X1 g_111_68 (.ZN (n_111_68), .A (n_115_66), .B (n_120_62), .C1 (n_116_64), .C2 (n_110_67) );
AOI211_X1 g_109_69 (.ZN (n_109_69), .A (n_113_67), .B (n_119_64), .C1 (n_118_63), .C2 (n_112_66) );
AOI211_X1 g_107_70 (.ZN (n_107_70), .A (n_111_68), .B (n_117_65), .C1 (n_120_62), .C2 (n_114_65) );
AOI211_X1 g_105_71 (.ZN (n_105_71), .A (n_109_69), .B (n_115_66), .C1 (n_119_64), .C2 (n_116_64) );
AOI211_X1 g_103_72 (.ZN (n_103_72), .A (n_107_70), .B (n_113_67), .C1 (n_117_65), .C2 (n_118_63) );
AOI211_X1 g_101_73 (.ZN (n_101_73), .A (n_105_71), .B (n_111_68), .C1 (n_115_66), .C2 (n_120_62) );
AOI211_X1 g_99_74 (.ZN (n_99_74), .A (n_103_72), .B (n_109_69), .C1 (n_113_67), .C2 (n_119_64) );
AOI211_X1 g_97_75 (.ZN (n_97_75), .A (n_101_73), .B (n_107_70), .C1 (n_111_68), .C2 (n_117_65) );
AOI211_X1 g_95_76 (.ZN (n_95_76), .A (n_99_74), .B (n_105_71), .C1 (n_109_69), .C2 (n_115_66) );
AOI211_X1 g_93_77 (.ZN (n_93_77), .A (n_97_75), .B (n_103_72), .C1 (n_107_70), .C2 (n_113_67) );
AOI211_X1 g_91_78 (.ZN (n_91_78), .A (n_95_76), .B (n_101_73), .C1 (n_105_71), .C2 (n_111_68) );
AOI211_X1 g_92_76 (.ZN (n_92_76), .A (n_93_77), .B (n_99_74), .C1 (n_103_72), .C2 (n_109_69) );
AOI211_X1 g_90_77 (.ZN (n_90_77), .A (n_91_78), .B (n_97_75), .C1 (n_101_73), .C2 (n_107_70) );
AOI211_X1 g_88_78 (.ZN (n_88_78), .A (n_92_76), .B (n_95_76), .C1 (n_99_74), .C2 (n_105_71) );
AOI211_X1 g_86_79 (.ZN (n_86_79), .A (n_90_77), .B (n_93_77), .C1 (n_97_75), .C2 (n_103_72) );
AOI211_X1 g_87_77 (.ZN (n_87_77), .A (n_88_78), .B (n_91_78), .C1 (n_95_76), .C2 (n_101_73) );
AOI211_X1 g_85_78 (.ZN (n_85_78), .A (n_86_79), .B (n_92_76), .C1 (n_93_77), .C2 (n_99_74) );
AOI211_X1 g_83_79 (.ZN (n_83_79), .A (n_87_77), .B (n_90_77), .C1 (n_91_78), .C2 (n_97_75) );
AOI211_X1 g_81_80 (.ZN (n_81_80), .A (n_85_78), .B (n_88_78), .C1 (n_92_76), .C2 (n_95_76) );
AOI211_X1 g_79_81 (.ZN (n_79_81), .A (n_83_79), .B (n_86_79), .C1 (n_90_77), .C2 (n_93_77) );
AOI211_X1 g_77_82 (.ZN (n_77_82), .A (n_81_80), .B (n_87_77), .C1 (n_88_78), .C2 (n_91_78) );
AOI211_X1 g_75_83 (.ZN (n_75_83), .A (n_79_81), .B (n_85_78), .C1 (n_86_79), .C2 (n_92_76) );
AOI211_X1 g_73_84 (.ZN (n_73_84), .A (n_77_82), .B (n_83_79), .C1 (n_87_77), .C2 (n_90_77) );
AOI211_X1 g_71_85 (.ZN (n_71_85), .A (n_75_83), .B (n_81_80), .C1 (n_85_78), .C2 (n_88_78) );
AOI211_X1 g_69_86 (.ZN (n_69_86), .A (n_73_84), .B (n_79_81), .C1 (n_83_79), .C2 (n_86_79) );
AOI211_X1 g_67_87 (.ZN (n_67_87), .A (n_71_85), .B (n_77_82), .C1 (n_81_80), .C2 (n_87_77) );
AOI211_X1 g_65_88 (.ZN (n_65_88), .A (n_69_86), .B (n_75_83), .C1 (n_79_81), .C2 (n_85_78) );
AOI211_X1 g_63_89 (.ZN (n_63_89), .A (n_67_87), .B (n_73_84), .C1 (n_77_82), .C2 (n_83_79) );
AOI211_X1 g_62_87 (.ZN (n_62_87), .A (n_65_88), .B (n_71_85), .C1 (n_75_83), .C2 (n_81_80) );
AOI211_X1 g_61_89 (.ZN (n_61_89), .A (n_63_89), .B (n_69_86), .C1 (n_73_84), .C2 (n_79_81) );
AOI211_X1 g_59_90 (.ZN (n_59_90), .A (n_62_87), .B (n_67_87), .C1 (n_71_85), .C2 (n_77_82) );
AOI211_X1 g_60_88 (.ZN (n_60_88), .A (n_61_89), .B (n_65_88), .C1 (n_69_86), .C2 (n_75_83) );
AOI211_X1 g_58_89 (.ZN (n_58_89), .A (n_59_90), .B (n_63_89), .C1 (n_67_87), .C2 (n_73_84) );
AOI211_X1 g_56_90 (.ZN (n_56_90), .A (n_60_88), .B (n_62_87), .C1 (n_65_88), .C2 (n_71_85) );
AOI211_X1 g_54_91 (.ZN (n_54_91), .A (n_58_89), .B (n_61_89), .C1 (n_63_89), .C2 (n_69_86) );
AOI211_X1 g_52_92 (.ZN (n_52_92), .A (n_56_90), .B (n_59_90), .C1 (n_62_87), .C2 (n_67_87) );
AOI211_X1 g_50_93 (.ZN (n_50_93), .A (n_54_91), .B (n_60_88), .C1 (n_61_89), .C2 (n_65_88) );
AOI211_X1 g_48_94 (.ZN (n_48_94), .A (n_52_92), .B (n_58_89), .C1 (n_59_90), .C2 (n_63_89) );
AOI211_X1 g_46_95 (.ZN (n_46_95), .A (n_50_93), .B (n_56_90), .C1 (n_60_88), .C2 (n_62_87) );
AOI211_X1 g_44_96 (.ZN (n_44_96), .A (n_48_94), .B (n_54_91), .C1 (n_58_89), .C2 (n_61_89) );
AOI211_X1 g_42_97 (.ZN (n_42_97), .A (n_46_95), .B (n_52_92), .C1 (n_56_90), .C2 (n_59_90) );
AOI211_X1 g_40_98 (.ZN (n_40_98), .A (n_44_96), .B (n_50_93), .C1 (n_54_91), .C2 (n_60_88) );
AOI211_X1 g_38_99 (.ZN (n_38_99), .A (n_42_97), .B (n_48_94), .C1 (n_52_92), .C2 (n_58_89) );
AOI211_X1 g_39_97 (.ZN (n_39_97), .A (n_40_98), .B (n_46_95), .C1 (n_50_93), .C2 (n_56_90) );
AOI211_X1 g_37_98 (.ZN (n_37_98), .A (n_38_99), .B (n_44_96), .C1 (n_48_94), .C2 (n_54_91) );
AOI211_X1 g_35_99 (.ZN (n_35_99), .A (n_39_97), .B (n_42_97), .C1 (n_46_95), .C2 (n_52_92) );
AOI211_X1 g_34_101 (.ZN (n_34_101), .A (n_37_98), .B (n_40_98), .C1 (n_44_96), .C2 (n_50_93) );
AOI211_X1 g_36_100 (.ZN (n_36_100), .A (n_35_99), .B (n_38_99), .C1 (n_42_97), .C2 (n_48_94) );
AOI211_X1 g_35_102 (.ZN (n_35_102), .A (n_34_101), .B (n_39_97), .C1 (n_40_98), .C2 (n_46_95) );
AOI211_X1 g_34_100 (.ZN (n_34_100), .A (n_36_100), .B (n_37_98), .C1 (n_38_99), .C2 (n_44_96) );
AOI211_X1 g_36_99 (.ZN (n_36_99), .A (n_35_102), .B (n_35_99), .C1 (n_39_97), .C2 (n_42_97) );
AOI211_X1 g_38_98 (.ZN (n_38_98), .A (n_34_100), .B (n_34_101), .C1 (n_37_98), .C2 (n_40_98) );
AOI211_X1 g_40_97 (.ZN (n_40_97), .A (n_36_99), .B (n_36_100), .C1 (n_35_99), .C2 (n_38_99) );
AOI211_X1 g_42_96 (.ZN (n_42_96), .A (n_38_98), .B (n_35_102), .C1 (n_34_101), .C2 (n_39_97) );
AOI211_X1 g_44_95 (.ZN (n_44_95), .A (n_40_97), .B (n_34_100), .C1 (n_36_100), .C2 (n_37_98) );
AOI211_X1 g_46_94 (.ZN (n_46_94), .A (n_42_96), .B (n_36_99), .C1 (n_35_102), .C2 (n_35_99) );
AOI211_X1 g_48_93 (.ZN (n_48_93), .A (n_44_95), .B (n_38_98), .C1 (n_34_100), .C2 (n_34_101) );
AOI211_X1 g_50_92 (.ZN (n_50_92), .A (n_46_94), .B (n_40_97), .C1 (n_36_99), .C2 (n_36_100) );
AOI211_X1 g_52_93 (.ZN (n_52_93), .A (n_48_93), .B (n_42_96), .C1 (n_38_98), .C2 (n_35_102) );
AOI211_X1 g_50_94 (.ZN (n_50_94), .A (n_50_92), .B (n_44_95), .C1 (n_40_97), .C2 (n_34_100) );
AOI211_X1 g_48_95 (.ZN (n_48_95), .A (n_52_93), .B (n_46_94), .C1 (n_42_96), .C2 (n_36_99) );
AOI211_X1 g_46_96 (.ZN (n_46_96), .A (n_50_94), .B (n_48_93), .C1 (n_44_95), .C2 (n_38_98) );
AOI211_X1 g_44_97 (.ZN (n_44_97), .A (n_48_95), .B (n_50_92), .C1 (n_46_94), .C2 (n_40_97) );
AOI211_X1 g_42_98 (.ZN (n_42_98), .A (n_46_96), .B (n_52_93), .C1 (n_48_93), .C2 (n_42_96) );
AOI211_X1 g_40_99 (.ZN (n_40_99), .A (n_44_97), .B (n_50_94), .C1 (n_50_92), .C2 (n_44_95) );
AOI211_X1 g_41_97 (.ZN (n_41_97), .A (n_42_98), .B (n_48_95), .C1 (n_52_93), .C2 (n_46_94) );
AOI211_X1 g_39_98 (.ZN (n_39_98), .A (n_40_99), .B (n_46_96), .C1 (n_50_94), .C2 (n_48_93) );
AOI211_X1 g_37_99 (.ZN (n_37_99), .A (n_41_97), .B (n_44_97), .C1 (n_48_95), .C2 (n_50_92) );
AOI211_X1 g_35_100 (.ZN (n_35_100), .A (n_39_98), .B (n_42_98), .C1 (n_46_96), .C2 (n_52_93) );
AOI211_X1 g_33_101 (.ZN (n_33_101), .A (n_37_99), .B (n_40_99), .C1 (n_44_97), .C2 (n_50_94) );
AOI211_X1 g_31_102 (.ZN (n_31_102), .A (n_35_100), .B (n_41_97), .C1 (n_42_98), .C2 (n_48_95) );
AOI211_X1 g_29_103 (.ZN (n_29_103), .A (n_33_101), .B (n_39_98), .C1 (n_40_99), .C2 (n_46_96) );
AOI211_X1 g_27_102 (.ZN (n_27_102), .A (n_31_102), .B (n_37_99), .C1 (n_41_97), .C2 (n_44_97) );
AOI211_X1 g_25_103 (.ZN (n_25_103), .A (n_29_103), .B (n_35_100), .C1 (n_39_98), .C2 (n_42_98) );
AOI211_X1 g_23_104 (.ZN (n_23_104), .A (n_27_102), .B (n_33_101), .C1 (n_37_99), .C2 (n_40_99) );
AOI211_X1 g_21_105 (.ZN (n_21_105), .A (n_25_103), .B (n_31_102), .C1 (n_35_100), .C2 (n_41_97) );
AOI211_X1 g_19_106 (.ZN (n_19_106), .A (n_23_104), .B (n_29_103), .C1 (n_33_101), .C2 (n_39_98) );
AOI211_X1 g_18_108 (.ZN (n_18_108), .A (n_21_105), .B (n_27_102), .C1 (n_31_102), .C2 (n_37_99) );
AOI211_X1 g_16_107 (.ZN (n_16_107), .A (n_19_106), .B (n_25_103), .C1 (n_29_103), .C2 (n_35_100) );
AOI211_X1 g_14_108 (.ZN (n_14_108), .A (n_18_108), .B (n_23_104), .C1 (n_27_102), .C2 (n_33_101) );
AOI211_X1 g_16_109 (.ZN (n_16_109), .A (n_16_107), .B (n_21_105), .C1 (n_25_103), .C2 (n_31_102) );
AOI211_X1 g_14_110 (.ZN (n_14_110), .A (n_14_108), .B (n_19_106), .C1 (n_23_104), .C2 (n_29_103) );
AOI211_X1 g_15_108 (.ZN (n_15_108), .A (n_16_109), .B (n_18_108), .C1 (n_21_105), .C2 (n_27_102) );
AOI211_X1 g_13_107 (.ZN (n_13_107), .A (n_14_110), .B (n_16_107), .C1 (n_19_106), .C2 (n_25_103) );
AOI211_X1 g_11_108 (.ZN (n_11_108), .A (n_15_108), .B (n_14_108), .C1 (n_18_108), .C2 (n_23_104) );
AOI211_X1 g_13_109 (.ZN (n_13_109), .A (n_13_107), .B (n_16_109), .C1 (n_16_107), .C2 (n_21_105) );
AOI211_X1 g_11_110 (.ZN (n_11_110), .A (n_11_108), .B (n_14_110), .C1 (n_14_108), .C2 (n_19_106) );
AOI211_X1 g_9_111 (.ZN (n_9_111), .A (n_13_109), .B (n_15_108), .C1 (n_16_109), .C2 (n_18_108) );
AOI211_X1 g_7_112 (.ZN (n_7_112), .A (n_11_110), .B (n_13_107), .C1 (n_14_110), .C2 (n_16_107) );
AOI211_X1 g_5_113 (.ZN (n_5_113), .A (n_9_111), .B (n_11_108), .C1 (n_15_108), .C2 (n_14_108) );
AOI211_X1 g_3_112 (.ZN (n_3_112), .A (n_7_112), .B (n_13_109), .C1 (n_13_107), .C2 (n_16_109) );
AOI211_X1 g_4_114 (.ZN (n_4_114), .A (n_5_113), .B (n_11_110), .C1 (n_11_108), .C2 (n_14_110) );
AOI211_X1 g_6_113 (.ZN (n_6_113), .A (n_3_112), .B (n_9_111), .C1 (n_13_109), .C2 (n_15_108) );
AOI211_X1 g_8_112 (.ZN (n_8_112), .A (n_4_114), .B (n_7_112), .C1 (n_11_110), .C2 (n_13_107) );
AOI211_X1 g_10_111 (.ZN (n_10_111), .A (n_6_113), .B (n_5_113), .C1 (n_9_111), .C2 (n_11_108) );
AOI211_X1 g_12_110 (.ZN (n_12_110), .A (n_8_112), .B (n_3_112), .C1 (n_7_112), .C2 (n_13_109) );
AOI211_X1 g_14_109 (.ZN (n_14_109), .A (n_10_111), .B (n_4_114), .C1 (n_5_113), .C2 (n_11_110) );
AOI211_X1 g_16_108 (.ZN (n_16_108), .A (n_12_110), .B (n_6_113), .C1 (n_3_112), .C2 (n_9_111) );
AOI211_X1 g_18_107 (.ZN (n_18_107), .A (n_14_109), .B (n_8_112), .C1 (n_4_114), .C2 (n_7_112) );
AOI211_X1 g_20_106 (.ZN (n_20_106), .A (n_16_108), .B (n_10_111), .C1 (n_6_113), .C2 (n_5_113) );
AOI211_X1 g_22_105 (.ZN (n_22_105), .A (n_18_107), .B (n_12_110), .C1 (n_8_112), .C2 (n_3_112) );
AOI211_X1 g_24_104 (.ZN (n_24_104), .A (n_20_106), .B (n_14_109), .C1 (n_10_111), .C2 (n_4_114) );
AOI211_X1 g_26_103 (.ZN (n_26_103), .A (n_22_105), .B (n_16_108), .C1 (n_12_110), .C2 (n_6_113) );
AOI211_X1 g_28_104 (.ZN (n_28_104), .A (n_24_104), .B (n_18_107), .C1 (n_14_109), .C2 (n_8_112) );
AOI211_X1 g_26_105 (.ZN (n_26_105), .A (n_26_103), .B (n_20_106), .C1 (n_16_108), .C2 (n_10_111) );
AOI211_X1 g_27_103 (.ZN (n_27_103), .A (n_28_104), .B (n_22_105), .C1 (n_18_107), .C2 (n_12_110) );
AOI211_X1 g_25_104 (.ZN (n_25_104), .A (n_26_105), .B (n_24_104), .C1 (n_20_106), .C2 (n_14_109) );
AOI211_X1 g_23_105 (.ZN (n_23_105), .A (n_27_103), .B (n_26_103), .C1 (n_22_105), .C2 (n_16_108) );
AOI211_X1 g_21_106 (.ZN (n_21_106), .A (n_25_104), .B (n_28_104), .C1 (n_24_104), .C2 (n_18_107) );
AOI211_X1 g_19_107 (.ZN (n_19_107), .A (n_23_105), .B (n_26_105), .C1 (n_26_103), .C2 (n_20_106) );
AOI211_X1 g_17_108 (.ZN (n_17_108), .A (n_21_106), .B (n_27_103), .C1 (n_28_104), .C2 (n_22_105) );
AOI211_X1 g_15_109 (.ZN (n_15_109), .A (n_19_107), .B (n_25_104), .C1 (n_26_105), .C2 (n_24_104) );
AOI211_X1 g_13_110 (.ZN (n_13_110), .A (n_17_108), .B (n_23_105), .C1 (n_27_103), .C2 (n_26_103) );
AOI211_X1 g_11_111 (.ZN (n_11_111), .A (n_15_109), .B (n_21_106), .C1 (n_25_104), .C2 (n_28_104) );
AOI211_X1 g_12_109 (.ZN (n_12_109), .A (n_13_110), .B (n_19_107), .C1 (n_23_105), .C2 (n_26_105) );
AOI211_X1 g_10_110 (.ZN (n_10_110), .A (n_11_111), .B (n_17_108), .C1 (n_21_106), .C2 (n_27_103) );
AOI211_X1 g_8_111 (.ZN (n_8_111), .A (n_12_109), .B (n_15_109), .C1 (n_19_107), .C2 (n_25_104) );
AOI211_X1 g_7_113 (.ZN (n_7_113), .A (n_10_110), .B (n_13_110), .C1 (n_17_108), .C2 (n_23_105) );
AOI211_X1 g_9_112 (.ZN (n_9_112), .A (n_8_111), .B (n_11_111), .C1 (n_15_109), .C2 (n_21_106) );
AOI211_X1 g_8_114 (.ZN (n_8_114), .A (n_7_113), .B (n_12_109), .C1 (n_13_110), .C2 (n_19_107) );
AOI211_X1 g_6_115 (.ZN (n_6_115), .A (n_9_112), .B (n_10_110), .C1 (n_11_111), .C2 (n_17_108) );
AOI211_X1 g_5_117 (.ZN (n_5_117), .A (n_8_114), .B (n_8_111), .C1 (n_12_109), .C2 (n_15_109) );
AOI211_X1 g_4_115 (.ZN (n_4_115), .A (n_6_115), .B (n_7_113), .C1 (n_10_110), .C2 (n_13_110) );
AOI211_X1 g_3_117 (.ZN (n_3_117), .A (n_5_117), .B (n_9_112), .C1 (n_8_111), .C2 (n_11_111) );
AOI211_X1 g_5_116 (.ZN (n_5_116), .A (n_4_115), .B (n_8_114), .C1 (n_7_113), .C2 (n_12_109) );
AOI211_X1 g_6_114 (.ZN (n_6_114), .A (n_3_117), .B (n_6_115), .C1 (n_9_112), .C2 (n_10_110) );
AOI211_X1 g_8_113 (.ZN (n_8_113), .A (n_5_116), .B (n_5_117), .C1 (n_8_114), .C2 (n_8_111) );
AOI211_X1 g_10_112 (.ZN (n_10_112), .A (n_6_114), .B (n_4_115), .C1 (n_6_115), .C2 (n_7_113) );
AOI211_X1 g_12_111 (.ZN (n_12_111), .A (n_8_113), .B (n_3_117), .C1 (n_5_117), .C2 (n_9_112) );
AOI211_X1 g_11_113 (.ZN (n_11_113), .A (n_10_112), .B (n_5_116), .C1 (n_4_115), .C2 (n_8_114) );
AOI211_X1 g_13_112 (.ZN (n_13_112), .A (n_12_111), .B (n_6_114), .C1 (n_3_117), .C2 (n_6_115) );
AOI211_X1 g_15_111 (.ZN (n_15_111), .A (n_11_113), .B (n_8_113), .C1 (n_5_116), .C2 (n_5_117) );
AOI211_X1 g_17_110 (.ZN (n_17_110), .A (n_13_112), .B (n_10_112), .C1 (n_6_114), .C2 (n_4_115) );
AOI211_X1 g_19_109 (.ZN (n_19_109), .A (n_15_111), .B (n_12_111), .C1 (n_8_113), .C2 (n_3_117) );
AOI211_X1 g_20_107 (.ZN (n_20_107), .A (n_17_110), .B (n_11_113), .C1 (n_10_112), .C2 (n_5_116) );
AOI211_X1 g_22_106 (.ZN (n_22_106), .A (n_19_109), .B (n_13_112), .C1 (n_12_111), .C2 (n_6_114) );
AOI211_X1 g_24_105 (.ZN (n_24_105), .A (n_20_107), .B (n_15_111), .C1 (n_11_113), .C2 (n_8_113) );
AOI211_X1 g_26_104 (.ZN (n_26_104), .A (n_22_106), .B (n_17_110), .C1 (n_13_112), .C2 (n_10_112) );
AOI211_X1 g_28_103 (.ZN (n_28_103), .A (n_24_105), .B (n_19_109), .C1 (n_15_111), .C2 (n_12_111) );
AOI211_X1 g_30_102 (.ZN (n_30_102), .A (n_26_104), .B (n_20_107), .C1 (n_17_110), .C2 (n_11_113) );
AOI211_X1 g_32_101 (.ZN (n_32_101), .A (n_28_103), .B (n_22_106), .C1 (n_19_109), .C2 (n_13_112) );
AOI211_X1 g_33_103 (.ZN (n_33_103), .A (n_30_102), .B (n_24_105), .C1 (n_20_107), .C2 (n_15_111) );
AOI211_X1 g_31_104 (.ZN (n_31_104), .A (n_32_101), .B (n_26_104), .C1 (n_22_106), .C2 (n_17_110) );
AOI211_X1 g_32_102 (.ZN (n_32_102), .A (n_33_103), .B (n_28_103), .C1 (n_24_105), .C2 (n_19_109) );
AOI211_X1 g_34_103 (.ZN (n_34_103), .A (n_31_104), .B (n_30_102), .C1 (n_26_104), .C2 (n_20_107) );
AOI211_X1 g_35_101 (.ZN (n_35_101), .A (n_32_102), .B (n_32_101), .C1 (n_28_103), .C2 (n_22_106) );
AOI211_X1 g_37_100 (.ZN (n_37_100), .A (n_34_103), .B (n_33_103), .C1 (n_30_102), .C2 (n_24_105) );
AOI211_X1 g_39_99 (.ZN (n_39_99), .A (n_35_101), .B (n_31_104), .C1 (n_32_101), .C2 (n_26_104) );
AOI211_X1 g_41_98 (.ZN (n_41_98), .A (n_37_100), .B (n_32_102), .C1 (n_33_103), .C2 (n_28_103) );
AOI211_X1 g_43_97 (.ZN (n_43_97), .A (n_39_99), .B (n_34_103), .C1 (n_31_104), .C2 (n_30_102) );
AOI211_X1 g_45_96 (.ZN (n_45_96), .A (n_41_98), .B (n_35_101), .C1 (n_32_102), .C2 (n_32_101) );
AOI211_X1 g_47_95 (.ZN (n_47_95), .A (n_43_97), .B (n_37_100), .C1 (n_34_103), .C2 (n_33_103) );
AOI211_X1 g_49_94 (.ZN (n_49_94), .A (n_45_96), .B (n_39_99), .C1 (n_35_101), .C2 (n_31_104) );
AOI211_X1 g_51_93 (.ZN (n_51_93), .A (n_47_95), .B (n_41_98), .C1 (n_37_100), .C2 (n_32_102) );
AOI211_X1 g_53_92 (.ZN (n_53_92), .A (n_49_94), .B (n_43_97), .C1 (n_39_99), .C2 (n_34_103) );
AOI211_X1 g_52_94 (.ZN (n_52_94), .A (n_51_93), .B (n_45_96), .C1 (n_41_98), .C2 (n_35_101) );
AOI211_X1 g_54_93 (.ZN (n_54_93), .A (n_53_92), .B (n_47_95), .C1 (n_43_97), .C2 (n_37_100) );
AOI211_X1 g_56_92 (.ZN (n_56_92), .A (n_52_94), .B (n_49_94), .C1 (n_45_96), .C2 (n_39_99) );
AOI211_X1 g_58_91 (.ZN (n_58_91), .A (n_54_93), .B (n_51_93), .C1 (n_47_95), .C2 (n_41_98) );
AOI211_X1 g_60_90 (.ZN (n_60_90), .A (n_56_92), .B (n_53_92), .C1 (n_49_94), .C2 (n_43_97) );
AOI211_X1 g_62_89 (.ZN (n_62_89), .A (n_58_91), .B (n_52_94), .C1 (n_51_93), .C2 (n_45_96) );
AOI211_X1 g_64_88 (.ZN (n_64_88), .A (n_60_90), .B (n_54_93), .C1 (n_53_92), .C2 (n_47_95) );
AOI211_X1 g_66_87 (.ZN (n_66_87), .A (n_62_89), .B (n_56_92), .C1 (n_52_94), .C2 (n_49_94) );
AOI211_X1 g_68_86 (.ZN (n_68_86), .A (n_64_88), .B (n_58_91), .C1 (n_54_93), .C2 (n_51_93) );
AOI211_X1 g_70_85 (.ZN (n_70_85), .A (n_66_87), .B (n_60_90), .C1 (n_56_92), .C2 (n_53_92) );
AOI211_X1 g_72_84 (.ZN (n_72_84), .A (n_68_86), .B (n_62_89), .C1 (n_58_91), .C2 (n_52_94) );
AOI211_X1 g_74_83 (.ZN (n_74_83), .A (n_70_85), .B (n_64_88), .C1 (n_60_90), .C2 (n_54_93) );
AOI211_X1 g_76_82 (.ZN (n_76_82), .A (n_72_84), .B (n_66_87), .C1 (n_62_89), .C2 (n_56_92) );
AOI211_X1 g_78_81 (.ZN (n_78_81), .A (n_74_83), .B (n_68_86), .C1 (n_64_88), .C2 (n_58_91) );
AOI211_X1 g_80_80 (.ZN (n_80_80), .A (n_76_82), .B (n_70_85), .C1 (n_66_87), .C2 (n_60_90) );
AOI211_X1 g_81_82 (.ZN (n_81_82), .A (n_78_81), .B (n_72_84), .C1 (n_68_86), .C2 (n_62_89) );
AOI211_X1 g_79_83 (.ZN (n_79_83), .A (n_80_80), .B (n_74_83), .C1 (n_70_85), .C2 (n_64_88) );
AOI211_X1 g_77_84 (.ZN (n_77_84), .A (n_81_82), .B (n_76_82), .C1 (n_72_84), .C2 (n_66_87) );
AOI211_X1 g_78_82 (.ZN (n_78_82), .A (n_79_83), .B (n_78_81), .C1 (n_74_83), .C2 (n_68_86) );
AOI211_X1 g_76_83 (.ZN (n_76_83), .A (n_77_84), .B (n_80_80), .C1 (n_76_82), .C2 (n_70_85) );
AOI211_X1 g_74_84 (.ZN (n_74_84), .A (n_78_82), .B (n_81_82), .C1 (n_78_81), .C2 (n_72_84) );
AOI211_X1 g_72_85 (.ZN (n_72_85), .A (n_76_83), .B (n_79_83), .C1 (n_80_80), .C2 (n_74_83) );
AOI211_X1 g_70_86 (.ZN (n_70_86), .A (n_74_84), .B (n_77_84), .C1 (n_81_82), .C2 (n_76_82) );
AOI211_X1 g_68_87 (.ZN (n_68_87), .A (n_72_85), .B (n_78_82), .C1 (n_79_83), .C2 (n_78_81) );
AOI211_X1 g_66_88 (.ZN (n_66_88), .A (n_70_86), .B (n_76_83), .C1 (n_77_84), .C2 (n_80_80) );
AOI211_X1 g_65_90 (.ZN (n_65_90), .A (n_68_87), .B (n_74_84), .C1 (n_78_82), .C2 (n_81_82) );
AOI211_X1 g_67_89 (.ZN (n_67_89), .A (n_66_88), .B (n_72_85), .C1 (n_76_83), .C2 (n_79_83) );
AOI211_X1 g_69_88 (.ZN (n_69_88), .A (n_65_90), .B (n_70_86), .C1 (n_74_84), .C2 (n_77_84) );
AOI211_X1 g_71_87 (.ZN (n_71_87), .A (n_67_89), .B (n_68_87), .C1 (n_72_85), .C2 (n_78_82) );
AOI211_X1 g_73_86 (.ZN (n_73_86), .A (n_69_88), .B (n_66_88), .C1 (n_70_86), .C2 (n_76_83) );
AOI211_X1 g_75_85 (.ZN (n_75_85), .A (n_71_87), .B (n_65_90), .C1 (n_68_87), .C2 (n_74_84) );
AOI211_X1 g_74_87 (.ZN (n_74_87), .A (n_73_86), .B (n_67_89), .C1 (n_66_88), .C2 (n_72_85) );
AOI211_X1 g_73_85 (.ZN (n_73_85), .A (n_75_85), .B (n_69_88), .C1 (n_65_90), .C2 (n_70_86) );
AOI211_X1 g_75_84 (.ZN (n_75_84), .A (n_74_87), .B (n_71_87), .C1 (n_67_89), .C2 (n_68_87) );
AOI211_X1 g_77_83 (.ZN (n_77_83), .A (n_73_85), .B (n_73_86), .C1 (n_69_88), .C2 (n_66_88) );
AOI211_X1 g_79_82 (.ZN (n_79_82), .A (n_75_84), .B (n_75_85), .C1 (n_71_87), .C2 (n_65_90) );
AOI211_X1 g_81_81 (.ZN (n_81_81), .A (n_77_83), .B (n_74_87), .C1 (n_73_86), .C2 (n_67_89) );
AOI211_X1 g_83_80 (.ZN (n_83_80), .A (n_79_82), .B (n_73_85), .C1 (n_75_85), .C2 (n_69_88) );
AOI211_X1 g_82_82 (.ZN (n_82_82), .A (n_81_81), .B (n_75_84), .C1 (n_74_87), .C2 (n_71_87) );
AOI211_X1 g_84_81 (.ZN (n_84_81), .A (n_83_80), .B (n_77_83), .C1 (n_73_85), .C2 (n_73_86) );
AOI211_X1 g_86_80 (.ZN (n_86_80), .A (n_82_82), .B (n_79_82), .C1 (n_75_84), .C2 (n_75_85) );
AOI211_X1 g_88_79 (.ZN (n_88_79), .A (n_84_81), .B (n_81_81), .C1 (n_77_83), .C2 (n_74_87) );
AOI211_X1 g_87_81 (.ZN (n_87_81), .A (n_86_80), .B (n_83_80), .C1 (n_79_82), .C2 (n_73_85) );
AOI211_X1 g_85_80 (.ZN (n_85_80), .A (n_88_79), .B (n_82_82), .C1 (n_81_81), .C2 (n_75_84) );
AOI211_X1 g_87_79 (.ZN (n_87_79), .A (n_87_81), .B (n_84_81), .C1 (n_83_80), .C2 (n_77_83) );
AOI211_X1 g_89_78 (.ZN (n_89_78), .A (n_85_80), .B (n_86_80), .C1 (n_82_82), .C2 (n_79_82) );
AOI211_X1 g_91_77 (.ZN (n_91_77), .A (n_87_79), .B (n_88_79), .C1 (n_84_81), .C2 (n_81_81) );
AOI211_X1 g_93_76 (.ZN (n_93_76), .A (n_89_78), .B (n_87_81), .C1 (n_86_80), .C2 (n_83_80) );
AOI211_X1 g_95_75 (.ZN (n_95_75), .A (n_91_77), .B (n_85_80), .C1 (n_88_79), .C2 (n_82_82) );
AOI211_X1 g_97_74 (.ZN (n_97_74), .A (n_93_76), .B (n_87_79), .C1 (n_87_81), .C2 (n_84_81) );
AOI211_X1 g_99_73 (.ZN (n_99_73), .A (n_95_75), .B (n_89_78), .C1 (n_85_80), .C2 (n_86_80) );
AOI211_X1 g_101_72 (.ZN (n_101_72), .A (n_97_74), .B (n_91_77), .C1 (n_87_79), .C2 (n_88_79) );
AOI211_X1 g_103_71 (.ZN (n_103_71), .A (n_99_73), .B (n_93_76), .C1 (n_89_78), .C2 (n_87_81) );
AOI211_X1 g_105_70 (.ZN (n_105_70), .A (n_101_72), .B (n_95_75), .C1 (n_91_77), .C2 (n_85_80) );
AOI211_X1 g_107_69 (.ZN (n_107_69), .A (n_103_71), .B (n_97_74), .C1 (n_93_76), .C2 (n_87_79) );
AOI211_X1 g_109_68 (.ZN (n_109_68), .A (n_105_70), .B (n_99_73), .C1 (n_95_75), .C2 (n_89_78) );
AOI211_X1 g_111_67 (.ZN (n_111_67), .A (n_107_69), .B (n_101_72), .C1 (n_97_74), .C2 (n_91_77) );
AOI211_X1 g_113_66 (.ZN (n_113_66), .A (n_109_68), .B (n_103_71), .C1 (n_99_73), .C2 (n_93_76) );
AOI211_X1 g_115_65 (.ZN (n_115_65), .A (n_111_67), .B (n_105_70), .C1 (n_101_72), .C2 (n_95_75) );
AOI211_X1 g_117_64 (.ZN (n_117_64), .A (n_113_66), .B (n_107_69), .C1 (n_103_71), .C2 (n_97_74) );
AOI211_X1 g_119_63 (.ZN (n_119_63), .A (n_115_65), .B (n_109_68), .C1 (n_105_70), .C2 (n_99_73) );
AOI211_X1 g_121_62 (.ZN (n_121_62), .A (n_117_64), .B (n_111_67), .C1 (n_107_69), .C2 (n_101_72) );
AOI211_X1 g_123_61 (.ZN (n_123_61), .A (n_119_63), .B (n_113_66), .C1 (n_109_68), .C2 (n_103_71) );
AOI211_X1 g_125_60 (.ZN (n_125_60), .A (n_121_62), .B (n_115_65), .C1 (n_111_67), .C2 (n_105_70) );
AOI211_X1 g_124_62 (.ZN (n_124_62), .A (n_123_61), .B (n_117_64), .C1 (n_113_66), .C2 (n_107_69) );
AOI211_X1 g_122_63 (.ZN (n_122_63), .A (n_125_60), .B (n_119_63), .C1 (n_115_65), .C2 (n_109_68) );
AOI211_X1 g_120_64 (.ZN (n_120_64), .A (n_124_62), .B (n_121_62), .C1 (n_117_64), .C2 (n_111_67) );
AOI211_X1 g_118_65 (.ZN (n_118_65), .A (n_122_63), .B (n_123_61), .C1 (n_119_63), .C2 (n_113_66) );
AOI211_X1 g_116_66 (.ZN (n_116_66), .A (n_120_64), .B (n_125_60), .C1 (n_121_62), .C2 (n_115_65) );
AOI211_X1 g_114_67 (.ZN (n_114_67), .A (n_118_65), .B (n_124_62), .C1 (n_123_61), .C2 (n_117_64) );
AOI211_X1 g_112_68 (.ZN (n_112_68), .A (n_116_66), .B (n_122_63), .C1 (n_125_60), .C2 (n_119_63) );
AOI211_X1 g_110_69 (.ZN (n_110_69), .A (n_114_67), .B (n_120_64), .C1 (n_124_62), .C2 (n_121_62) );
AOI211_X1 g_108_70 (.ZN (n_108_70), .A (n_112_68), .B (n_118_65), .C1 (n_122_63), .C2 (n_123_61) );
AOI211_X1 g_106_71 (.ZN (n_106_71), .A (n_110_69), .B (n_116_66), .C1 (n_120_64), .C2 (n_125_60) );
AOI211_X1 g_104_72 (.ZN (n_104_72), .A (n_108_70), .B (n_114_67), .C1 (n_118_65), .C2 (n_124_62) );
AOI211_X1 g_102_73 (.ZN (n_102_73), .A (n_106_71), .B (n_112_68), .C1 (n_116_66), .C2 (n_122_63) );
AOI211_X1 g_100_74 (.ZN (n_100_74), .A (n_104_72), .B (n_110_69), .C1 (n_114_67), .C2 (n_120_64) );
AOI211_X1 g_98_75 (.ZN (n_98_75), .A (n_102_73), .B (n_108_70), .C1 (n_112_68), .C2 (n_118_65) );
AOI211_X1 g_96_76 (.ZN (n_96_76), .A (n_100_74), .B (n_106_71), .C1 (n_110_69), .C2 (n_116_66) );
AOI211_X1 g_94_77 (.ZN (n_94_77), .A (n_98_75), .B (n_104_72), .C1 (n_108_70), .C2 (n_114_67) );
AOI211_X1 g_92_78 (.ZN (n_92_78), .A (n_96_76), .B (n_102_73), .C1 (n_106_71), .C2 (n_112_68) );
AOI211_X1 g_90_79 (.ZN (n_90_79), .A (n_94_77), .B (n_100_74), .C1 (n_104_72), .C2 (n_110_69) );
AOI211_X1 g_88_80 (.ZN (n_88_80), .A (n_92_78), .B (n_98_75), .C1 (n_102_73), .C2 (n_108_70) );
AOI211_X1 g_86_81 (.ZN (n_86_81), .A (n_90_79), .B (n_96_76), .C1 (n_100_74), .C2 (n_106_71) );
AOI211_X1 g_84_80 (.ZN (n_84_80), .A (n_88_80), .B (n_94_77), .C1 (n_98_75), .C2 (n_104_72) );
AOI211_X1 g_82_81 (.ZN (n_82_81), .A (n_86_81), .B (n_92_78), .C1 (n_96_76), .C2 (n_102_73) );
AOI211_X1 g_80_82 (.ZN (n_80_82), .A (n_84_80), .B (n_90_79), .C1 (n_94_77), .C2 (n_100_74) );
AOI211_X1 g_78_83 (.ZN (n_78_83), .A (n_82_81), .B (n_88_80), .C1 (n_92_78), .C2 (n_98_75) );
AOI211_X1 g_76_84 (.ZN (n_76_84), .A (n_80_82), .B (n_86_81), .C1 (n_90_79), .C2 (n_96_76) );
AOI211_X1 g_74_85 (.ZN (n_74_85), .A (n_78_83), .B (n_84_80), .C1 (n_88_80), .C2 (n_94_77) );
AOI211_X1 g_72_86 (.ZN (n_72_86), .A (n_76_84), .B (n_82_81), .C1 (n_86_81), .C2 (n_92_78) );
AOI211_X1 g_70_87 (.ZN (n_70_87), .A (n_74_85), .B (n_80_82), .C1 (n_84_80), .C2 (n_90_79) );
AOI211_X1 g_68_88 (.ZN (n_68_88), .A (n_72_86), .B (n_78_83), .C1 (n_82_81), .C2 (n_88_80) );
AOI211_X1 g_66_89 (.ZN (n_66_89), .A (n_70_87), .B (n_76_84), .C1 (n_80_82), .C2 (n_86_81) );
AOI211_X1 g_64_90 (.ZN (n_64_90), .A (n_68_88), .B (n_74_85), .C1 (n_78_83), .C2 (n_84_80) );
AOI211_X1 g_62_91 (.ZN (n_62_91), .A (n_66_89), .B (n_72_86), .C1 (n_76_84), .C2 (n_82_81) );
AOI211_X1 g_60_92 (.ZN (n_60_92), .A (n_64_90), .B (n_70_87), .C1 (n_74_85), .C2 (n_80_82) );
AOI211_X1 g_61_90 (.ZN (n_61_90), .A (n_62_91), .B (n_68_88), .C1 (n_72_86), .C2 (n_78_83) );
AOI211_X1 g_59_91 (.ZN (n_59_91), .A (n_60_92), .B (n_66_89), .C1 (n_70_87), .C2 (n_76_84) );
AOI211_X1 g_57_92 (.ZN (n_57_92), .A (n_61_90), .B (n_64_90), .C1 (n_68_88), .C2 (n_74_85) );
AOI211_X1 g_55_93 (.ZN (n_55_93), .A (n_59_91), .B (n_62_91), .C1 (n_66_89), .C2 (n_72_86) );
AOI211_X1 g_53_94 (.ZN (n_53_94), .A (n_57_92), .B (n_60_92), .C1 (n_64_90), .C2 (n_70_87) );
AOI211_X1 g_51_95 (.ZN (n_51_95), .A (n_55_93), .B (n_61_90), .C1 (n_62_91), .C2 (n_68_88) );
AOI211_X1 g_49_96 (.ZN (n_49_96), .A (n_53_94), .B (n_59_91), .C1 (n_60_92), .C2 (n_66_89) );
AOI211_X1 g_47_97 (.ZN (n_47_97), .A (n_51_95), .B (n_57_92), .C1 (n_61_90), .C2 (n_64_90) );
AOI211_X1 g_45_98 (.ZN (n_45_98), .A (n_49_96), .B (n_55_93), .C1 (n_59_91), .C2 (n_62_91) );
AOI211_X1 g_43_99 (.ZN (n_43_99), .A (n_47_97), .B (n_53_94), .C1 (n_57_92), .C2 (n_60_92) );
AOI211_X1 g_41_100 (.ZN (n_41_100), .A (n_45_98), .B (n_51_95), .C1 (n_55_93), .C2 (n_61_90) );
AOI211_X1 g_39_101 (.ZN (n_39_101), .A (n_43_99), .B (n_49_96), .C1 (n_53_94), .C2 (n_59_91) );
AOI211_X1 g_37_102 (.ZN (n_37_102), .A (n_41_100), .B (n_47_97), .C1 (n_51_95), .C2 (n_57_92) );
AOI211_X1 g_38_100 (.ZN (n_38_100), .A (n_39_101), .B (n_45_98), .C1 (n_49_96), .C2 (n_55_93) );
AOI211_X1 g_36_101 (.ZN (n_36_101), .A (n_37_102), .B (n_43_99), .C1 (n_47_97), .C2 (n_53_94) );
AOI211_X1 g_34_102 (.ZN (n_34_102), .A (n_38_100), .B (n_41_100), .C1 (n_45_98), .C2 (n_51_95) );
AOI211_X1 g_32_103 (.ZN (n_32_103), .A (n_36_101), .B (n_39_101), .C1 (n_43_99), .C2 (n_49_96) );
AOI211_X1 g_30_104 (.ZN (n_30_104), .A (n_34_102), .B (n_37_102), .C1 (n_41_100), .C2 (n_47_97) );
AOI211_X1 g_28_105 (.ZN (n_28_105), .A (n_32_103), .B (n_38_100), .C1 (n_39_101), .C2 (n_45_98) );
AOI211_X1 g_26_106 (.ZN (n_26_106), .A (n_30_104), .B (n_36_101), .C1 (n_37_102), .C2 (n_43_99) );
AOI211_X1 g_27_104 (.ZN (n_27_104), .A (n_28_105), .B (n_34_102), .C1 (n_38_100), .C2 (n_41_100) );
AOI211_X1 g_25_105 (.ZN (n_25_105), .A (n_26_106), .B (n_32_103), .C1 (n_36_101), .C2 (n_39_101) );
AOI211_X1 g_23_106 (.ZN (n_23_106), .A (n_27_104), .B (n_30_104), .C1 (n_34_102), .C2 (n_37_102) );
AOI211_X1 g_21_107 (.ZN (n_21_107), .A (n_25_105), .B (n_28_105), .C1 (n_32_103), .C2 (n_38_100) );
AOI211_X1 g_19_108 (.ZN (n_19_108), .A (n_23_106), .B (n_26_106), .C1 (n_30_104), .C2 (n_36_101) );
AOI211_X1 g_17_109 (.ZN (n_17_109), .A (n_21_107), .B (n_27_104), .C1 (n_28_105), .C2 (n_34_102) );
AOI211_X1 g_15_110 (.ZN (n_15_110), .A (n_19_108), .B (n_25_105), .C1 (n_26_106), .C2 (n_32_103) );
AOI211_X1 g_13_111 (.ZN (n_13_111), .A (n_17_109), .B (n_23_106), .C1 (n_27_104), .C2 (n_30_104) );
AOI211_X1 g_11_112 (.ZN (n_11_112), .A (n_15_110), .B (n_21_107), .C1 (n_25_105), .C2 (n_28_105) );
AOI211_X1 g_9_113 (.ZN (n_9_113), .A (n_13_111), .B (n_19_108), .C1 (n_23_106), .C2 (n_26_106) );
AOI211_X1 g_7_114 (.ZN (n_7_114), .A (n_11_112), .B (n_17_109), .C1 (n_21_107), .C2 (n_27_104) );
AOI211_X1 g_5_115 (.ZN (n_5_115), .A (n_9_113), .B (n_15_110), .C1 (n_19_108), .C2 (n_25_105) );
AOI211_X1 g_3_116 (.ZN (n_3_116), .A (n_7_114), .B (n_13_111), .C1 (n_17_109), .C2 (n_23_106) );
AOI211_X1 g_2_118 (.ZN (n_2_118), .A (n_5_115), .B (n_11_112), .C1 (n_15_110), .C2 (n_21_107) );
AOI211_X1 g_1_120 (.ZN (n_1_120), .A (n_3_116), .B (n_9_113), .C1 (n_13_111), .C2 (n_19_108) );
AOI211_X1 g_3_119 (.ZN (n_3_119), .A (n_2_118), .B (n_7_114), .C1 (n_11_112), .C2 (n_17_109) );
AOI211_X1 g_4_117 (.ZN (n_4_117), .A (n_1_120), .B (n_5_115), .C1 (n_9_113), .C2 (n_15_110) );
AOI211_X1 g_6_116 (.ZN (n_6_116), .A (n_3_119), .B (n_3_116), .C1 (n_7_114), .C2 (n_13_111) );
AOI211_X1 g_5_118 (.ZN (n_5_118), .A (n_4_117), .B (n_2_118), .C1 (n_5_115), .C2 (n_11_112) );
AOI211_X1 g_7_117 (.ZN (n_7_117), .A (n_6_116), .B (n_1_120), .C1 (n_3_116), .C2 (n_9_113) );
AOI211_X1 g_8_115 (.ZN (n_8_115), .A (n_5_118), .B (n_3_119), .C1 (n_2_118), .C2 (n_7_114) );
AOI211_X1 g_10_114 (.ZN (n_10_114), .A (n_7_117), .B (n_4_117), .C1 (n_1_120), .C2 (n_5_115) );
AOI211_X1 g_12_113 (.ZN (n_12_113), .A (n_8_115), .B (n_6_116), .C1 (n_3_119), .C2 (n_3_116) );
AOI211_X1 g_14_112 (.ZN (n_14_112), .A (n_10_114), .B (n_5_118), .C1 (n_4_117), .C2 (n_2_118) );
AOI211_X1 g_16_111 (.ZN (n_16_111), .A (n_12_113), .B (n_7_117), .C1 (n_6_116), .C2 (n_1_120) );
AOI211_X1 g_18_110 (.ZN (n_18_110), .A (n_14_112), .B (n_8_115), .C1 (n_5_118), .C2 (n_3_119) );
AOI211_X1 g_20_109 (.ZN (n_20_109), .A (n_16_111), .B (n_10_114), .C1 (n_7_117), .C2 (n_4_117) );
AOI211_X1 g_22_108 (.ZN (n_22_108), .A (n_18_110), .B (n_12_113), .C1 (n_8_115), .C2 (n_6_116) );
AOI211_X1 g_24_107 (.ZN (n_24_107), .A (n_20_109), .B (n_14_112), .C1 (n_10_114), .C2 (n_5_118) );
AOI211_X1 g_23_109 (.ZN (n_23_109), .A (n_22_108), .B (n_16_111), .C1 (n_12_113), .C2 (n_7_117) );
AOI211_X1 g_21_108 (.ZN (n_21_108), .A (n_24_107), .B (n_18_110), .C1 (n_14_112), .C2 (n_8_115) );
AOI211_X1 g_23_107 (.ZN (n_23_107), .A (n_23_109), .B (n_20_109), .C1 (n_16_111), .C2 (n_10_114) );
AOI211_X1 g_25_106 (.ZN (n_25_106), .A (n_21_108), .B (n_22_108), .C1 (n_18_110), .C2 (n_12_113) );
AOI211_X1 g_27_105 (.ZN (n_27_105), .A (n_23_107), .B (n_24_107), .C1 (n_20_109), .C2 (n_14_112) );
AOI211_X1 g_29_104 (.ZN (n_29_104), .A (n_25_106), .B (n_23_109), .C1 (n_22_108), .C2 (n_16_111) );
AOI211_X1 g_31_103 (.ZN (n_31_103), .A (n_27_105), .B (n_21_108), .C1 (n_24_107), .C2 (n_18_110) );
AOI211_X1 g_33_102 (.ZN (n_33_102), .A (n_29_104), .B (n_23_107), .C1 (n_23_109), .C2 (n_20_109) );
AOI211_X1 g_32_104 (.ZN (n_32_104), .A (n_31_103), .B (n_25_106), .C1 (n_21_108), .C2 (n_22_108) );
AOI211_X1 g_30_105 (.ZN (n_30_105), .A (n_33_102), .B (n_27_105), .C1 (n_23_107), .C2 (n_24_107) );
AOI211_X1 g_28_106 (.ZN (n_28_106), .A (n_32_104), .B (n_29_104), .C1 (n_25_106), .C2 (n_23_109) );
AOI211_X1 g_26_107 (.ZN (n_26_107), .A (n_30_105), .B (n_31_103), .C1 (n_27_105), .C2 (n_21_108) );
AOI211_X1 g_24_106 (.ZN (n_24_106), .A (n_28_106), .B (n_33_102), .C1 (n_29_104), .C2 (n_23_107) );
AOI211_X1 g_22_107 (.ZN (n_22_107), .A (n_26_107), .B (n_32_104), .C1 (n_31_103), .C2 (n_25_106) );
AOI211_X1 g_20_108 (.ZN (n_20_108), .A (n_24_106), .B (n_30_105), .C1 (n_33_102), .C2 (n_27_105) );
AOI211_X1 g_18_109 (.ZN (n_18_109), .A (n_22_107), .B (n_28_106), .C1 (n_32_104), .C2 (n_29_104) );
AOI211_X1 g_16_110 (.ZN (n_16_110), .A (n_20_108), .B (n_26_107), .C1 (n_30_105), .C2 (n_31_103) );
AOI211_X1 g_14_111 (.ZN (n_14_111), .A (n_18_109), .B (n_24_106), .C1 (n_28_106), .C2 (n_33_102) );
AOI211_X1 g_12_112 (.ZN (n_12_112), .A (n_16_110), .B (n_22_107), .C1 (n_26_107), .C2 (n_32_104) );
AOI211_X1 g_10_113 (.ZN (n_10_113), .A (n_14_111), .B (n_20_108), .C1 (n_24_106), .C2 (n_30_105) );
AOI211_X1 g_9_115 (.ZN (n_9_115), .A (n_12_112), .B (n_18_109), .C1 (n_22_107), .C2 (n_28_106) );
AOI211_X1 g_7_116 (.ZN (n_7_116), .A (n_10_113), .B (n_16_110), .C1 (n_20_108), .C2 (n_26_107) );
AOI211_X1 g_6_118 (.ZN (n_6_118), .A (n_9_115), .B (n_14_111), .C1 (n_18_109), .C2 (n_24_106) );
AOI211_X1 g_4_119 (.ZN (n_4_119), .A (n_7_116), .B (n_12_112), .C1 (n_16_110), .C2 (n_22_107) );
AOI211_X1 g_3_121 (.ZN (n_3_121), .A (n_6_118), .B (n_10_113), .C1 (n_14_111), .C2 (n_20_108) );
AOI211_X1 g_5_120 (.ZN (n_5_120), .A (n_4_119), .B (n_9_115), .C1 (n_12_112), .C2 (n_18_109) );
AOI211_X1 g_4_118 (.ZN (n_4_118), .A (n_3_121), .B (n_7_116), .C1 (n_10_113), .C2 (n_16_110) );
AOI211_X1 g_3_120 (.ZN (n_3_120), .A (n_5_120), .B (n_6_118), .C1 (n_9_115), .C2 (n_14_111) );
AOI211_X1 g_2_122 (.ZN (n_2_122), .A (n_4_118), .B (n_4_119), .C1 (n_7_116), .C2 (n_12_112) );
AOI211_X1 g_1_124 (.ZN (n_1_124), .A (n_3_120), .B (n_3_121), .C1 (n_6_118), .C2 (n_10_113) );
AOI211_X1 g_3_123 (.ZN (n_3_123), .A (n_2_122), .B (n_5_120), .C1 (n_4_119), .C2 (n_9_115) );
AOI211_X1 g_5_122 (.ZN (n_5_122), .A (n_1_124), .B (n_4_118), .C1 (n_3_121), .C2 (n_7_116) );
AOI211_X1 g_6_120 (.ZN (n_6_120), .A (n_3_123), .B (n_3_120), .C1 (n_5_120), .C2 (n_6_118) );
AOI211_X1 g_4_121 (.ZN (n_4_121), .A (n_5_122), .B (n_2_122), .C1 (n_4_118), .C2 (n_4_119) );
AOI211_X1 g_5_119 (.ZN (n_5_119), .A (n_6_120), .B (n_1_124), .C1 (n_3_120), .C2 (n_3_121) );
AOI211_X1 g_7_118 (.ZN (n_7_118), .A (n_4_121), .B (n_3_123), .C1 (n_2_122), .C2 (n_5_120) );
AOI211_X1 g_9_117 (.ZN (n_9_117), .A (n_5_119), .B (n_5_122), .C1 (n_1_124), .C2 (n_4_118) );
AOI211_X1 g_10_115 (.ZN (n_10_115), .A (n_7_118), .B (n_6_120), .C1 (n_3_123), .C2 (n_3_120) );
AOI211_X1 g_12_114 (.ZN (n_12_114), .A (n_9_117), .B (n_4_121), .C1 (n_5_122), .C2 (n_2_122) );
AOI211_X1 g_14_113 (.ZN (n_14_113), .A (n_10_115), .B (n_5_119), .C1 (n_6_120), .C2 (n_1_124) );
AOI211_X1 g_16_112 (.ZN (n_16_112), .A (n_12_114), .B (n_7_118), .C1 (n_4_121), .C2 (n_3_123) );
AOI211_X1 g_18_111 (.ZN (n_18_111), .A (n_14_113), .B (n_9_117), .C1 (n_5_119), .C2 (n_5_122) );
AOI211_X1 g_20_110 (.ZN (n_20_110), .A (n_16_112), .B (n_10_115), .C1 (n_7_118), .C2 (n_6_120) );
AOI211_X1 g_22_109 (.ZN (n_22_109), .A (n_18_111), .B (n_12_114), .C1 (n_9_117), .C2 (n_4_121) );
AOI211_X1 g_24_108 (.ZN (n_24_108), .A (n_20_110), .B (n_14_113), .C1 (n_10_115), .C2 (n_5_119) );
AOI211_X1 g_23_110 (.ZN (n_23_110), .A (n_22_109), .B (n_16_112), .C1 (n_12_114), .C2 (n_7_118) );
AOI211_X1 g_21_109 (.ZN (n_21_109), .A (n_24_108), .B (n_18_111), .C1 (n_14_113), .C2 (n_9_117) );
AOI211_X1 g_23_108 (.ZN (n_23_108), .A (n_23_110), .B (n_20_110), .C1 (n_16_112), .C2 (n_10_115) );
AOI211_X1 g_25_107 (.ZN (n_25_107), .A (n_21_109), .B (n_22_109), .C1 (n_18_111), .C2 (n_12_114) );
AOI211_X1 g_27_106 (.ZN (n_27_106), .A (n_23_108), .B (n_24_108), .C1 (n_20_110), .C2 (n_14_113) );
AOI211_X1 g_29_105 (.ZN (n_29_105), .A (n_25_107), .B (n_23_110), .C1 (n_22_109), .C2 (n_16_112) );
AOI211_X1 g_28_107 (.ZN (n_28_107), .A (n_27_106), .B (n_21_109), .C1 (n_24_108), .C2 (n_18_111) );
AOI211_X1 g_30_106 (.ZN (n_30_106), .A (n_29_105), .B (n_23_108), .C1 (n_23_110), .C2 (n_20_110) );
AOI211_X1 g_32_105 (.ZN (n_32_105), .A (n_28_107), .B (n_25_107), .C1 (n_21_109), .C2 (n_22_109) );
AOI211_X1 g_34_104 (.ZN (n_34_104), .A (n_30_106), .B (n_27_106), .C1 (n_23_108), .C2 (n_24_108) );
AOI211_X1 g_36_103 (.ZN (n_36_103), .A (n_32_105), .B (n_29_105), .C1 (n_25_107), .C2 (n_23_110) );
AOI211_X1 g_37_101 (.ZN (n_37_101), .A (n_34_104), .B (n_28_107), .C1 (n_27_106), .C2 (n_21_109) );
AOI211_X1 g_39_100 (.ZN (n_39_100), .A (n_36_103), .B (n_30_106), .C1 (n_29_105), .C2 (n_23_108) );
AOI211_X1 g_41_99 (.ZN (n_41_99), .A (n_37_101), .B (n_32_105), .C1 (n_28_107), .C2 (n_25_107) );
AOI211_X1 g_43_98 (.ZN (n_43_98), .A (n_39_100), .B (n_34_104), .C1 (n_30_106), .C2 (n_27_106) );
AOI211_X1 g_45_97 (.ZN (n_45_97), .A (n_41_99), .B (n_36_103), .C1 (n_32_105), .C2 (n_29_105) );
AOI211_X1 g_47_96 (.ZN (n_47_96), .A (n_43_98), .B (n_37_101), .C1 (n_34_104), .C2 (n_28_107) );
AOI211_X1 g_49_95 (.ZN (n_49_95), .A (n_45_97), .B (n_39_100), .C1 (n_36_103), .C2 (n_30_106) );
AOI211_X1 g_51_94 (.ZN (n_51_94), .A (n_47_96), .B (n_41_99), .C1 (n_37_101), .C2 (n_32_105) );
AOI211_X1 g_53_93 (.ZN (n_53_93), .A (n_49_95), .B (n_43_98), .C1 (n_39_100), .C2 (n_34_104) );
AOI211_X1 g_55_92 (.ZN (n_55_92), .A (n_51_94), .B (n_45_97), .C1 (n_41_99), .C2 (n_36_103) );
AOI211_X1 g_57_91 (.ZN (n_57_91), .A (n_53_93), .B (n_47_96), .C1 (n_43_98), .C2 (n_37_101) );
AOI211_X1 g_56_93 (.ZN (n_56_93), .A (n_55_92), .B (n_49_95), .C1 (n_45_97), .C2 (n_39_100) );
AOI211_X1 g_54_94 (.ZN (n_54_94), .A (n_57_91), .B (n_51_94), .C1 (n_47_96), .C2 (n_41_99) );
AOI211_X1 g_52_95 (.ZN (n_52_95), .A (n_56_93), .B (n_53_93), .C1 (n_49_95), .C2 (n_43_98) );
AOI211_X1 g_50_96 (.ZN (n_50_96), .A (n_54_94), .B (n_55_92), .C1 (n_51_94), .C2 (n_45_97) );
AOI211_X1 g_48_97 (.ZN (n_48_97), .A (n_52_95), .B (n_57_91), .C1 (n_53_93), .C2 (n_47_96) );
AOI211_X1 g_46_98 (.ZN (n_46_98), .A (n_50_96), .B (n_56_93), .C1 (n_55_92), .C2 (n_49_95) );
AOI211_X1 g_44_99 (.ZN (n_44_99), .A (n_48_97), .B (n_54_94), .C1 (n_57_91), .C2 (n_51_94) );
AOI211_X1 g_42_100 (.ZN (n_42_100), .A (n_46_98), .B (n_52_95), .C1 (n_56_93), .C2 (n_53_93) );
AOI211_X1 g_40_101 (.ZN (n_40_101), .A (n_44_99), .B (n_50_96), .C1 (n_54_94), .C2 (n_55_92) );
AOI211_X1 g_38_102 (.ZN (n_38_102), .A (n_42_100), .B (n_48_97), .C1 (n_52_95), .C2 (n_57_91) );
AOI211_X1 g_40_103 (.ZN (n_40_103), .A (n_40_101), .B (n_46_98), .C1 (n_50_96), .C2 (n_56_93) );
AOI211_X1 g_42_102 (.ZN (n_42_102), .A (n_38_102), .B (n_44_99), .C1 (n_48_97), .C2 (n_54_94) );
AOI211_X1 g_44_101 (.ZN (n_44_101), .A (n_40_103), .B (n_42_100), .C1 (n_46_98), .C2 (n_52_95) );
AOI211_X1 g_46_100 (.ZN (n_46_100), .A (n_42_102), .B (n_40_101), .C1 (n_44_99), .C2 (n_50_96) );
AOI211_X1 g_48_99 (.ZN (n_48_99), .A (n_44_101), .B (n_38_102), .C1 (n_42_100), .C2 (n_48_97) );
AOI211_X1 g_50_98 (.ZN (n_50_98), .A (n_46_100), .B (n_40_103), .C1 (n_40_101), .C2 (n_46_98) );
AOI211_X1 g_51_96 (.ZN (n_51_96), .A (n_48_99), .B (n_42_102), .C1 (n_38_102), .C2 (n_44_99) );
AOI211_X1 g_53_95 (.ZN (n_53_95), .A (n_50_98), .B (n_44_101), .C1 (n_40_103), .C2 (n_42_100) );
AOI211_X1 g_55_94 (.ZN (n_55_94), .A (n_51_96), .B (n_46_100), .C1 (n_42_102), .C2 (n_40_101) );
AOI211_X1 g_57_93 (.ZN (n_57_93), .A (n_53_95), .B (n_48_99), .C1 (n_44_101), .C2 (n_38_102) );
AOI211_X1 g_59_92 (.ZN (n_59_92), .A (n_55_94), .B (n_50_98), .C1 (n_46_100), .C2 (n_40_103) );
AOI211_X1 g_61_91 (.ZN (n_61_91), .A (n_57_93), .B (n_51_96), .C1 (n_48_99), .C2 (n_42_102) );
AOI211_X1 g_63_90 (.ZN (n_63_90), .A (n_59_92), .B (n_53_95), .C1 (n_50_98), .C2 (n_44_101) );
AOI211_X1 g_65_89 (.ZN (n_65_89), .A (n_61_91), .B (n_55_94), .C1 (n_51_96), .C2 (n_46_100) );
AOI211_X1 g_67_88 (.ZN (n_67_88), .A (n_63_90), .B (n_57_93), .C1 (n_53_95), .C2 (n_48_99) );
AOI211_X1 g_69_87 (.ZN (n_69_87), .A (n_65_89), .B (n_59_92), .C1 (n_55_94), .C2 (n_50_98) );
AOI211_X1 g_71_86 (.ZN (n_71_86), .A (n_67_88), .B (n_61_91), .C1 (n_57_93), .C2 (n_51_96) );
AOI211_X1 g_72_88 (.ZN (n_72_88), .A (n_69_87), .B (n_63_90), .C1 (n_59_92), .C2 (n_53_95) );
AOI211_X1 g_70_89 (.ZN (n_70_89), .A (n_71_86), .B (n_65_89), .C1 (n_61_91), .C2 (n_55_94) );
AOI211_X1 g_68_90 (.ZN (n_68_90), .A (n_72_88), .B (n_67_88), .C1 (n_63_90), .C2 (n_57_93) );
AOI211_X1 g_66_91 (.ZN (n_66_91), .A (n_70_89), .B (n_69_87), .C1 (n_65_89), .C2 (n_59_92) );
AOI211_X1 g_64_92 (.ZN (n_64_92), .A (n_68_90), .B (n_71_86), .C1 (n_67_88), .C2 (n_61_91) );
AOI211_X1 g_62_93 (.ZN (n_62_93), .A (n_66_91), .B (n_72_88), .C1 (n_69_87), .C2 (n_63_90) );
AOI211_X1 g_63_91 (.ZN (n_63_91), .A (n_64_92), .B (n_70_89), .C1 (n_71_86), .C2 (n_65_89) );
AOI211_X1 g_61_92 (.ZN (n_61_92), .A (n_62_93), .B (n_68_90), .C1 (n_72_88), .C2 (n_67_88) );
AOI211_X1 g_59_93 (.ZN (n_59_93), .A (n_63_91), .B (n_66_91), .C1 (n_70_89), .C2 (n_69_87) );
AOI211_X1 g_57_94 (.ZN (n_57_94), .A (n_61_92), .B (n_64_92), .C1 (n_68_90), .C2 (n_71_86) );
AOI211_X1 g_55_95 (.ZN (n_55_95), .A (n_59_93), .B (n_62_93), .C1 (n_66_91), .C2 (n_72_88) );
AOI211_X1 g_53_96 (.ZN (n_53_96), .A (n_57_94), .B (n_63_91), .C1 (n_64_92), .C2 (n_70_89) );
AOI211_X1 g_51_97 (.ZN (n_51_97), .A (n_55_95), .B (n_61_92), .C1 (n_62_93), .C2 (n_68_90) );
AOI211_X1 g_50_95 (.ZN (n_50_95), .A (n_53_96), .B (n_59_93), .C1 (n_63_91), .C2 (n_66_91) );
AOI211_X1 g_49_97 (.ZN (n_49_97), .A (n_51_97), .B (n_57_94), .C1 (n_61_92), .C2 (n_64_92) );
AOI211_X1 g_47_98 (.ZN (n_47_98), .A (n_50_95), .B (n_55_95), .C1 (n_59_93), .C2 (n_62_93) );
AOI211_X1 g_48_96 (.ZN (n_48_96), .A (n_49_97), .B (n_53_96), .C1 (n_57_94), .C2 (n_63_91) );
AOI211_X1 g_46_97 (.ZN (n_46_97), .A (n_47_98), .B (n_51_97), .C1 (n_55_95), .C2 (n_61_92) );
AOI211_X1 g_45_99 (.ZN (n_45_99), .A (n_48_96), .B (n_50_95), .C1 (n_53_96), .C2 (n_59_93) );
AOI211_X1 g_43_100 (.ZN (n_43_100), .A (n_46_97), .B (n_49_97), .C1 (n_51_97), .C2 (n_57_94) );
AOI211_X1 g_44_98 (.ZN (n_44_98), .A (n_45_99), .B (n_47_98), .C1 (n_50_95), .C2 (n_55_95) );
AOI211_X1 g_42_99 (.ZN (n_42_99), .A (n_43_100), .B (n_48_96), .C1 (n_49_97), .C2 (n_53_96) );
AOI211_X1 g_41_101 (.ZN (n_41_101), .A (n_44_98), .B (n_46_97), .C1 (n_47_98), .C2 (n_51_97) );
AOI211_X1 g_39_102 (.ZN (n_39_102), .A (n_42_99), .B (n_45_99), .C1 (n_48_96), .C2 (n_50_95) );
AOI211_X1 g_40_100 (.ZN (n_40_100), .A (n_41_101), .B (n_43_100), .C1 (n_46_97), .C2 (n_49_97) );
AOI211_X1 g_38_101 (.ZN (n_38_101), .A (n_39_102), .B (n_44_98), .C1 (n_45_99), .C2 (n_47_98) );
AOI211_X1 g_36_102 (.ZN (n_36_102), .A (n_40_100), .B (n_42_99), .C1 (n_43_100), .C2 (n_48_96) );
AOI211_X1 g_35_104 (.ZN (n_35_104), .A (n_38_101), .B (n_41_101), .C1 (n_44_98), .C2 (n_46_97) );
AOI211_X1 g_37_103 (.ZN (n_37_103), .A (n_36_102), .B (n_39_102), .C1 (n_42_99), .C2 (n_45_99) );
AOI211_X1 g_36_105 (.ZN (n_36_105), .A (n_35_104), .B (n_40_100), .C1 (n_41_101), .C2 (n_43_100) );
AOI211_X1 g_38_104 (.ZN (n_38_104), .A (n_37_103), .B (n_38_101), .C1 (n_39_102), .C2 (n_44_98) );
AOI211_X1 g_37_106 (.ZN (n_37_106), .A (n_36_105), .B (n_36_102), .C1 (n_40_100), .C2 (n_42_99) );
AOI211_X1 g_36_104 (.ZN (n_36_104), .A (n_38_104), .B (n_35_104), .C1 (n_38_101), .C2 (n_41_101) );
AOI211_X1 g_38_103 (.ZN (n_38_103), .A (n_37_106), .B (n_37_103), .C1 (n_36_102), .C2 (n_39_102) );
AOI211_X1 g_40_102 (.ZN (n_40_102), .A (n_36_104), .B (n_36_105), .C1 (n_35_104), .C2 (n_40_100) );
AOI211_X1 g_42_101 (.ZN (n_42_101), .A (n_38_103), .B (n_38_104), .C1 (n_37_103), .C2 (n_38_101) );
AOI211_X1 g_44_100 (.ZN (n_44_100), .A (n_40_102), .B (n_37_106), .C1 (n_36_105), .C2 (n_36_102) );
AOI211_X1 g_46_99 (.ZN (n_46_99), .A (n_42_101), .B (n_36_104), .C1 (n_38_104), .C2 (n_35_104) );
AOI211_X1 g_48_98 (.ZN (n_48_98), .A (n_44_100), .B (n_38_103), .C1 (n_37_106), .C2 (n_37_103) );
AOI211_X1 g_50_97 (.ZN (n_50_97), .A (n_46_99), .B (n_40_102), .C1 (n_36_104), .C2 (n_36_105) );
AOI211_X1 g_52_96 (.ZN (n_52_96), .A (n_48_98), .B (n_42_101), .C1 (n_38_103), .C2 (n_38_104) );
AOI211_X1 g_54_95 (.ZN (n_54_95), .A (n_50_97), .B (n_44_100), .C1 (n_40_102), .C2 (n_37_106) );
AOI211_X1 g_56_94 (.ZN (n_56_94), .A (n_52_96), .B (n_46_99), .C1 (n_42_101), .C2 (n_36_104) );
AOI211_X1 g_58_93 (.ZN (n_58_93), .A (n_54_95), .B (n_48_98), .C1 (n_44_100), .C2 (n_38_103) );
AOI211_X1 g_60_94 (.ZN (n_60_94), .A (n_56_94), .B (n_50_97), .C1 (n_46_99), .C2 (n_40_102) );
AOI211_X1 g_58_95 (.ZN (n_58_95), .A (n_58_93), .B (n_52_96), .C1 (n_48_98), .C2 (n_42_101) );
AOI211_X1 g_56_96 (.ZN (n_56_96), .A (n_60_94), .B (n_54_95), .C1 (n_50_97), .C2 (n_44_100) );
AOI211_X1 g_54_97 (.ZN (n_54_97), .A (n_58_95), .B (n_56_94), .C1 (n_52_96), .C2 (n_46_99) );
AOI211_X1 g_52_98 (.ZN (n_52_98), .A (n_56_96), .B (n_58_93), .C1 (n_54_95), .C2 (n_48_98) );
AOI211_X1 g_50_99 (.ZN (n_50_99), .A (n_54_97), .B (n_60_94), .C1 (n_56_94), .C2 (n_50_97) );
AOI211_X1 g_48_100 (.ZN (n_48_100), .A (n_52_98), .B (n_58_95), .C1 (n_58_93), .C2 (n_52_96) );
AOI211_X1 g_49_98 (.ZN (n_49_98), .A (n_50_99), .B (n_56_96), .C1 (n_60_94), .C2 (n_54_95) );
AOI211_X1 g_47_99 (.ZN (n_47_99), .A (n_48_100), .B (n_54_97), .C1 (n_58_95), .C2 (n_56_94) );
AOI211_X1 g_45_100 (.ZN (n_45_100), .A (n_49_98), .B (n_52_98), .C1 (n_56_96), .C2 (n_58_93) );
AOI211_X1 g_43_101 (.ZN (n_43_101), .A (n_47_99), .B (n_50_99), .C1 (n_54_97), .C2 (n_60_94) );
AOI211_X1 g_41_102 (.ZN (n_41_102), .A (n_45_100), .B (n_48_100), .C1 (n_52_98), .C2 (n_58_95) );
AOI211_X1 g_39_103 (.ZN (n_39_103), .A (n_43_101), .B (n_49_98), .C1 (n_50_99), .C2 (n_56_96) );
AOI211_X1 g_37_104 (.ZN (n_37_104), .A (n_41_102), .B (n_47_99), .C1 (n_48_100), .C2 (n_54_97) );
AOI211_X1 g_35_103 (.ZN (n_35_103), .A (n_39_103), .B (n_45_100), .C1 (n_49_98), .C2 (n_52_98) );
AOI211_X1 g_33_104 (.ZN (n_33_104), .A (n_37_104), .B (n_43_101), .C1 (n_47_99), .C2 (n_50_99) );
AOI211_X1 g_35_105 (.ZN (n_35_105), .A (n_35_103), .B (n_41_102), .C1 (n_45_100), .C2 (n_48_100) );
AOI211_X1 g_33_106 (.ZN (n_33_106), .A (n_33_104), .B (n_39_103), .C1 (n_43_101), .C2 (n_49_98) );
AOI211_X1 g_31_105 (.ZN (n_31_105), .A (n_35_105), .B (n_37_104), .C1 (n_41_102), .C2 (n_47_99) );
AOI211_X1 g_29_106 (.ZN (n_29_106), .A (n_33_106), .B (n_35_103), .C1 (n_39_103), .C2 (n_45_100) );
AOI211_X1 g_27_107 (.ZN (n_27_107), .A (n_31_105), .B (n_33_104), .C1 (n_37_104), .C2 (n_43_101) );
AOI211_X1 g_25_108 (.ZN (n_25_108), .A (n_29_106), .B (n_35_105), .C1 (n_35_103), .C2 (n_41_102) );
AOI211_X1 g_24_110 (.ZN (n_24_110), .A (n_27_107), .B (n_33_106), .C1 (n_33_104), .C2 (n_39_103) );
AOI211_X1 g_26_109 (.ZN (n_26_109), .A (n_25_108), .B (n_31_105), .C1 (n_35_105), .C2 (n_37_104) );
AOI211_X1 g_28_108 (.ZN (n_28_108), .A (n_24_110), .B (n_29_106), .C1 (n_33_106), .C2 (n_35_103) );
AOI211_X1 g_30_107 (.ZN (n_30_107), .A (n_26_109), .B (n_27_107), .C1 (n_31_105), .C2 (n_33_104) );
AOI211_X1 g_32_106 (.ZN (n_32_106), .A (n_28_108), .B (n_25_108), .C1 (n_29_106), .C2 (n_35_105) );
AOI211_X1 g_34_105 (.ZN (n_34_105), .A (n_30_107), .B (n_24_110), .C1 (n_27_107), .C2 (n_33_106) );
AOI211_X1 g_35_107 (.ZN (n_35_107), .A (n_32_106), .B (n_26_109), .C1 (n_25_108), .C2 (n_31_105) );
AOI211_X1 g_33_108 (.ZN (n_33_108), .A (n_34_105), .B (n_28_108), .C1 (n_24_110), .C2 (n_29_106) );
AOI211_X1 g_34_106 (.ZN (n_34_106), .A (n_35_107), .B (n_30_107), .C1 (n_26_109), .C2 (n_27_107) );
AOI211_X1 g_32_107 (.ZN (n_32_107), .A (n_33_108), .B (n_32_106), .C1 (n_28_108), .C2 (n_25_108) );
AOI211_X1 g_33_105 (.ZN (n_33_105), .A (n_34_106), .B (n_34_105), .C1 (n_30_107), .C2 (n_24_110) );
AOI211_X1 g_31_106 (.ZN (n_31_106), .A (n_32_107), .B (n_35_107), .C1 (n_32_106), .C2 (n_26_109) );
AOI211_X1 g_29_107 (.ZN (n_29_107), .A (n_33_105), .B (n_33_108), .C1 (n_34_105), .C2 (n_28_108) );
AOI211_X1 g_27_108 (.ZN (n_27_108), .A (n_31_106), .B (n_34_106), .C1 (n_35_107), .C2 (n_30_107) );
AOI211_X1 g_25_109 (.ZN (n_25_109), .A (n_29_107), .B (n_32_107), .C1 (n_33_108), .C2 (n_32_106) );
AOI211_X1 g_24_111 (.ZN (n_24_111), .A (n_27_108), .B (n_33_105), .C1 (n_34_106), .C2 (n_34_105) );
AOI211_X1 g_22_110 (.ZN (n_22_110), .A (n_25_109), .B (n_31_106), .C1 (n_32_107), .C2 (n_35_107) );
AOI211_X1 g_24_109 (.ZN (n_24_109), .A (n_24_111), .B (n_29_107), .C1 (n_33_105), .C2 (n_33_108) );
AOI211_X1 g_26_108 (.ZN (n_26_108), .A (n_22_110), .B (n_27_108), .C1 (n_31_106), .C2 (n_34_106) );
AOI211_X1 g_25_110 (.ZN (n_25_110), .A (n_24_109), .B (n_25_109), .C1 (n_29_107), .C2 (n_32_107) );
AOI211_X1 g_27_109 (.ZN (n_27_109), .A (n_26_108), .B (n_24_111), .C1 (n_27_108), .C2 (n_33_105) );
AOI211_X1 g_29_108 (.ZN (n_29_108), .A (n_25_110), .B (n_22_110), .C1 (n_25_109), .C2 (n_31_106) );
AOI211_X1 g_31_107 (.ZN (n_31_107), .A (n_27_109), .B (n_24_109), .C1 (n_24_111), .C2 (n_29_107) );
AOI211_X1 g_30_109 (.ZN (n_30_109), .A (n_29_108), .B (n_26_108), .C1 (n_22_110), .C2 (n_27_108) );
AOI211_X1 g_32_108 (.ZN (n_32_108), .A (n_31_107), .B (n_25_110), .C1 (n_24_109), .C2 (n_25_109) );
AOI211_X1 g_34_107 (.ZN (n_34_107), .A (n_30_109), .B (n_27_109), .C1 (n_26_108), .C2 (n_24_111) );
AOI211_X1 g_36_106 (.ZN (n_36_106), .A (n_32_108), .B (n_29_108), .C1 (n_25_110), .C2 (n_22_110) );
AOI211_X1 g_38_105 (.ZN (n_38_105), .A (n_34_107), .B (n_31_107), .C1 (n_27_109), .C2 (n_24_109) );
AOI211_X1 g_40_104 (.ZN (n_40_104), .A (n_36_106), .B (n_30_109), .C1 (n_29_108), .C2 (n_26_108) );
AOI211_X1 g_42_103 (.ZN (n_42_103), .A (n_38_105), .B (n_32_108), .C1 (n_31_107), .C2 (n_25_110) );
AOI211_X1 g_44_102 (.ZN (n_44_102), .A (n_40_104), .B (n_34_107), .C1 (n_30_109), .C2 (n_27_109) );
AOI211_X1 g_46_101 (.ZN (n_46_101), .A (n_42_103), .B (n_36_106), .C1 (n_32_108), .C2 (n_29_108) );
AOI211_X1 g_45_103 (.ZN (n_45_103), .A (n_44_102), .B (n_38_105), .C1 (n_34_107), .C2 (n_31_107) );
AOI211_X1 g_43_102 (.ZN (n_43_102), .A (n_46_101), .B (n_40_104), .C1 (n_36_106), .C2 (n_30_109) );
AOI211_X1 g_45_101 (.ZN (n_45_101), .A (n_45_103), .B (n_42_103), .C1 (n_38_105), .C2 (n_32_108) );
AOI211_X1 g_47_100 (.ZN (n_47_100), .A (n_43_102), .B (n_44_102), .C1 (n_40_104), .C2 (n_34_107) );
AOI211_X1 g_49_99 (.ZN (n_49_99), .A (n_45_101), .B (n_46_101), .C1 (n_42_103), .C2 (n_36_106) );
AOI211_X1 g_51_98 (.ZN (n_51_98), .A (n_47_100), .B (n_45_103), .C1 (n_44_102), .C2 (n_38_105) );
AOI211_X1 g_53_97 (.ZN (n_53_97), .A (n_49_99), .B (n_43_102), .C1 (n_46_101), .C2 (n_40_104) );
AOI211_X1 g_55_96 (.ZN (n_55_96), .A (n_51_98), .B (n_45_101), .C1 (n_45_103), .C2 (n_42_103) );
AOI211_X1 g_57_95 (.ZN (n_57_95), .A (n_53_97), .B (n_47_100), .C1 (n_43_102), .C2 (n_44_102) );
AOI211_X1 g_59_94 (.ZN (n_59_94), .A (n_55_96), .B (n_49_99), .C1 (n_45_101), .C2 (n_46_101) );
AOI211_X1 g_61_93 (.ZN (n_61_93), .A (n_57_95), .B (n_51_98), .C1 (n_47_100), .C2 (n_45_103) );
AOI211_X1 g_63_92 (.ZN (n_63_92), .A (n_59_94), .B (n_53_97), .C1 (n_49_99), .C2 (n_43_102) );
AOI211_X1 g_65_91 (.ZN (n_65_91), .A (n_61_93), .B (n_55_96), .C1 (n_51_98), .C2 (n_45_101) );
AOI211_X1 g_67_90 (.ZN (n_67_90), .A (n_63_92), .B (n_57_95), .C1 (n_53_97), .C2 (n_47_100) );
AOI211_X1 g_69_89 (.ZN (n_69_89), .A (n_65_91), .B (n_59_94), .C1 (n_55_96), .C2 (n_49_99) );
AOI211_X1 g_71_88 (.ZN (n_71_88), .A (n_67_90), .B (n_61_93), .C1 (n_57_95), .C2 (n_51_98) );
AOI211_X1 g_73_87 (.ZN (n_73_87), .A (n_69_89), .B (n_63_92), .C1 (n_59_94), .C2 (n_53_97) );
AOI211_X1 g_75_86 (.ZN (n_75_86), .A (n_71_88), .B (n_65_91), .C1 (n_61_93), .C2 (n_55_96) );
AOI211_X1 g_77_85 (.ZN (n_77_85), .A (n_73_87), .B (n_67_90), .C1 (n_63_92), .C2 (n_57_95) );
AOI211_X1 g_79_84 (.ZN (n_79_84), .A (n_75_86), .B (n_69_89), .C1 (n_65_91), .C2 (n_59_94) );
AOI211_X1 g_81_83 (.ZN (n_81_83), .A (n_77_85), .B (n_71_88), .C1 (n_67_90), .C2 (n_61_93) );
AOI211_X1 g_83_82 (.ZN (n_83_82), .A (n_79_84), .B (n_73_87), .C1 (n_69_89), .C2 (n_63_92) );
AOI211_X1 g_85_81 (.ZN (n_85_81), .A (n_81_83), .B (n_75_86), .C1 (n_71_88), .C2 (n_65_91) );
AOI211_X1 g_87_80 (.ZN (n_87_80), .A (n_83_82), .B (n_77_85), .C1 (n_73_87), .C2 (n_67_90) );
AOI211_X1 g_89_79 (.ZN (n_89_79), .A (n_85_81), .B (n_79_84), .C1 (n_75_86), .C2 (n_69_89) );
AOI211_X1 g_88_81 (.ZN (n_88_81), .A (n_87_80), .B (n_81_83), .C1 (n_77_85), .C2 (n_71_88) );
AOI211_X1 g_90_80 (.ZN (n_90_80), .A (n_89_79), .B (n_83_82), .C1 (n_79_84), .C2 (n_73_87) );
AOI211_X1 g_92_79 (.ZN (n_92_79), .A (n_88_81), .B (n_85_81), .C1 (n_81_83), .C2 (n_75_86) );
AOI211_X1 g_94_78 (.ZN (n_94_78), .A (n_90_80), .B (n_87_80), .C1 (n_83_82), .C2 (n_77_85) );
AOI211_X1 g_92_77 (.ZN (n_92_77), .A (n_92_79), .B (n_89_79), .C1 (n_85_81), .C2 (n_79_84) );
AOI211_X1 g_94_76 (.ZN (n_94_76), .A (n_94_78), .B (n_88_81), .C1 (n_87_80), .C2 (n_81_83) );
AOI211_X1 g_96_75 (.ZN (n_96_75), .A (n_92_77), .B (n_90_80), .C1 (n_89_79), .C2 (n_83_82) );
AOI211_X1 g_98_74 (.ZN (n_98_74), .A (n_94_76), .B (n_92_79), .C1 (n_88_81), .C2 (n_85_81) );
AOI211_X1 g_100_73 (.ZN (n_100_73), .A (n_96_75), .B (n_94_78), .C1 (n_90_80), .C2 (n_87_80) );
AOI211_X1 g_102_72 (.ZN (n_102_72), .A (n_98_74), .B (n_92_77), .C1 (n_92_79), .C2 (n_89_79) );
AOI211_X1 g_104_71 (.ZN (n_104_71), .A (n_100_73), .B (n_94_76), .C1 (n_94_78), .C2 (n_88_81) );
AOI211_X1 g_106_70 (.ZN (n_106_70), .A (n_102_72), .B (n_96_75), .C1 (n_92_77), .C2 (n_90_80) );
AOI211_X1 g_105_72 (.ZN (n_105_72), .A (n_104_71), .B (n_98_74), .C1 (n_94_76), .C2 (n_92_79) );
AOI211_X1 g_107_71 (.ZN (n_107_71), .A (n_106_70), .B (n_100_73), .C1 (n_96_75), .C2 (n_94_78) );
AOI211_X1 g_109_70 (.ZN (n_109_70), .A (n_105_72), .B (n_102_72), .C1 (n_98_74), .C2 (n_92_77) );
AOI211_X1 g_110_68 (.ZN (n_110_68), .A (n_107_71), .B (n_104_71), .C1 (n_100_73), .C2 (n_94_76) );
AOI211_X1 g_112_67 (.ZN (n_112_67), .A (n_109_70), .B (n_106_70), .C1 (n_102_72), .C2 (n_96_75) );
AOI211_X1 g_114_66 (.ZN (n_114_66), .A (n_110_68), .B (n_105_72), .C1 (n_104_71), .C2 (n_98_74) );
AOI211_X1 g_116_65 (.ZN (n_116_65), .A (n_112_67), .B (n_107_71), .C1 (n_106_70), .C2 (n_100_73) );
AOI211_X1 g_118_64 (.ZN (n_118_64), .A (n_114_66), .B (n_109_70), .C1 (n_105_72), .C2 (n_102_72) );
AOI211_X1 g_120_63 (.ZN (n_120_63), .A (n_116_65), .B (n_110_68), .C1 (n_107_71), .C2 (n_104_71) );
AOI211_X1 g_122_62 (.ZN (n_122_62), .A (n_118_64), .B (n_112_67), .C1 (n_109_70), .C2 (n_106_70) );
AOI211_X1 g_124_61 (.ZN (n_124_61), .A (n_120_63), .B (n_114_66), .C1 (n_110_68), .C2 (n_105_72) );
AOI211_X1 g_126_60 (.ZN (n_126_60), .A (n_122_62), .B (n_116_65), .C1 (n_112_67), .C2 (n_107_71) );
AOI211_X1 g_128_59 (.ZN (n_128_59), .A (n_124_61), .B (n_118_64), .C1 (n_114_66), .C2 (n_109_70) );
AOI211_X1 g_129_61 (.ZN (n_129_61), .A (n_126_60), .B (n_120_63), .C1 (n_116_65), .C2 (n_110_68) );
AOI211_X1 g_127_62 (.ZN (n_127_62), .A (n_128_59), .B (n_122_62), .C1 (n_118_64), .C2 (n_112_67) );
AOI211_X1 g_125_63 (.ZN (n_125_63), .A (n_129_61), .B (n_124_61), .C1 (n_120_63), .C2 (n_114_66) );
AOI211_X1 g_123_64 (.ZN (n_123_64), .A (n_127_62), .B (n_126_60), .C1 (n_122_62), .C2 (n_116_65) );
AOI211_X1 g_121_65 (.ZN (n_121_65), .A (n_125_63), .B (n_128_59), .C1 (n_124_61), .C2 (n_118_64) );
AOI211_X1 g_119_66 (.ZN (n_119_66), .A (n_123_64), .B (n_129_61), .C1 (n_126_60), .C2 (n_120_63) );
AOI211_X1 g_117_67 (.ZN (n_117_67), .A (n_121_65), .B (n_127_62), .C1 (n_128_59), .C2 (n_122_62) );
AOI211_X1 g_115_68 (.ZN (n_115_68), .A (n_119_66), .B (n_125_63), .C1 (n_129_61), .C2 (n_124_61) );
AOI211_X1 g_113_69 (.ZN (n_113_69), .A (n_117_67), .B (n_123_64), .C1 (n_127_62), .C2 (n_126_60) );
AOI211_X1 g_111_70 (.ZN (n_111_70), .A (n_115_68), .B (n_121_65), .C1 (n_125_63), .C2 (n_128_59) );
AOI211_X1 g_109_71 (.ZN (n_109_71), .A (n_113_69), .B (n_119_66), .C1 (n_123_64), .C2 (n_129_61) );
AOI211_X1 g_107_72 (.ZN (n_107_72), .A (n_111_70), .B (n_117_67), .C1 (n_121_65), .C2 (n_127_62) );
AOI211_X1 g_105_73 (.ZN (n_105_73), .A (n_109_71), .B (n_115_68), .C1 (n_119_66), .C2 (n_125_63) );
AOI211_X1 g_103_74 (.ZN (n_103_74), .A (n_107_72), .B (n_113_69), .C1 (n_117_67), .C2 (n_123_64) );
AOI211_X1 g_101_75 (.ZN (n_101_75), .A (n_105_73), .B (n_111_70), .C1 (n_115_68), .C2 (n_121_65) );
AOI211_X1 g_99_76 (.ZN (n_99_76), .A (n_103_74), .B (n_109_71), .C1 (n_113_69), .C2 (n_119_66) );
AOI211_X1 g_97_77 (.ZN (n_97_77), .A (n_101_75), .B (n_107_72), .C1 (n_111_70), .C2 (n_117_67) );
AOI211_X1 g_95_78 (.ZN (n_95_78), .A (n_99_76), .B (n_105_73), .C1 (n_109_71), .C2 (n_115_68) );
AOI211_X1 g_93_79 (.ZN (n_93_79), .A (n_97_77), .B (n_103_74), .C1 (n_107_72), .C2 (n_113_69) );
AOI211_X1 g_91_80 (.ZN (n_91_80), .A (n_95_78), .B (n_101_75), .C1 (n_105_73), .C2 (n_111_70) );
AOI211_X1 g_89_81 (.ZN (n_89_81), .A (n_93_79), .B (n_99_76), .C1 (n_103_74), .C2 (n_109_71) );
AOI211_X1 g_87_82 (.ZN (n_87_82), .A (n_91_80), .B (n_97_77), .C1 (n_101_75), .C2 (n_107_72) );
AOI211_X1 g_85_83 (.ZN (n_85_83), .A (n_89_81), .B (n_95_78), .C1 (n_99_76), .C2 (n_105_73) );
AOI211_X1 g_83_84 (.ZN (n_83_84), .A (n_87_82), .B (n_93_79), .C1 (n_97_77), .C2 (n_103_74) );
AOI211_X1 g_84_82 (.ZN (n_84_82), .A (n_85_83), .B (n_91_80), .C1 (n_95_78), .C2 (n_101_75) );
AOI211_X1 g_82_83 (.ZN (n_82_83), .A (n_83_84), .B (n_89_81), .C1 (n_93_79), .C2 (n_99_76) );
AOI211_X1 g_80_84 (.ZN (n_80_84), .A (n_84_82), .B (n_87_82), .C1 (n_91_80), .C2 (n_97_77) );
AOI211_X1 g_78_85 (.ZN (n_78_85), .A (n_82_83), .B (n_85_83), .C1 (n_89_81), .C2 (n_95_78) );
AOI211_X1 g_76_86 (.ZN (n_76_86), .A (n_80_84), .B (n_83_84), .C1 (n_87_82), .C2 (n_93_79) );
AOI211_X1 g_75_88 (.ZN (n_75_88), .A (n_78_85), .B (n_84_82), .C1 (n_85_83), .C2 (n_91_80) );
AOI211_X1 g_74_86 (.ZN (n_74_86), .A (n_76_86), .B (n_82_83), .C1 (n_83_84), .C2 (n_89_81) );
AOI211_X1 g_76_85 (.ZN (n_76_85), .A (n_75_88), .B (n_80_84), .C1 (n_84_82), .C2 (n_87_82) );
AOI211_X1 g_78_84 (.ZN (n_78_84), .A (n_74_86), .B (n_78_85), .C1 (n_82_83), .C2 (n_85_83) );
AOI211_X1 g_80_83 (.ZN (n_80_83), .A (n_76_85), .B (n_76_86), .C1 (n_80_84), .C2 (n_83_84) );
AOI211_X1 g_81_85 (.ZN (n_81_85), .A (n_78_84), .B (n_75_88), .C1 (n_78_85), .C2 (n_84_82) );
AOI211_X1 g_79_86 (.ZN (n_79_86), .A (n_80_83), .B (n_74_86), .C1 (n_76_86), .C2 (n_82_83) );
AOI211_X1 g_77_87 (.ZN (n_77_87), .A (n_81_85), .B (n_76_85), .C1 (n_75_88), .C2 (n_80_84) );
AOI211_X1 g_76_89 (.ZN (n_76_89), .A (n_79_86), .B (n_78_84), .C1 (n_74_86), .C2 (n_78_85) );
AOI211_X1 g_75_87 (.ZN (n_75_87), .A (n_77_87), .B (n_80_83), .C1 (n_76_85), .C2 (n_76_86) );
AOI211_X1 g_77_86 (.ZN (n_77_86), .A (n_76_89), .B (n_81_85), .C1 (n_78_84), .C2 (n_75_88) );
AOI211_X1 g_79_85 (.ZN (n_79_85), .A (n_75_87), .B (n_79_86), .C1 (n_80_83), .C2 (n_74_86) );
AOI211_X1 g_81_84 (.ZN (n_81_84), .A (n_77_86), .B (n_77_87), .C1 (n_81_85), .C2 (n_76_85) );
AOI211_X1 g_83_83 (.ZN (n_83_83), .A (n_79_85), .B (n_76_89), .C1 (n_79_86), .C2 (n_78_84) );
AOI211_X1 g_85_82 (.ZN (n_85_82), .A (n_81_84), .B (n_75_87), .C1 (n_77_87), .C2 (n_80_83) );
AOI211_X1 g_84_84 (.ZN (n_84_84), .A (n_83_83), .B (n_77_86), .C1 (n_76_89), .C2 (n_81_85) );
AOI211_X1 g_86_83 (.ZN (n_86_83), .A (n_85_82), .B (n_79_85), .C1 (n_75_87), .C2 (n_79_86) );
AOI211_X1 g_88_82 (.ZN (n_88_82), .A (n_84_84), .B (n_81_84), .C1 (n_77_86), .C2 (n_77_87) );
AOI211_X1 g_89_80 (.ZN (n_89_80), .A (n_86_83), .B (n_83_83), .C1 (n_79_85), .C2 (n_76_89) );
AOI211_X1 g_91_79 (.ZN (n_91_79), .A (n_88_82), .B (n_85_82), .C1 (n_81_84), .C2 (n_75_87) );
AOI211_X1 g_93_78 (.ZN (n_93_78), .A (n_89_80), .B (n_84_84), .C1 (n_83_83), .C2 (n_77_86) );
AOI211_X1 g_95_77 (.ZN (n_95_77), .A (n_91_79), .B (n_86_83), .C1 (n_85_82), .C2 (n_79_85) );
AOI211_X1 g_97_76 (.ZN (n_97_76), .A (n_93_78), .B (n_88_82), .C1 (n_84_84), .C2 (n_81_84) );
AOI211_X1 g_99_75 (.ZN (n_99_75), .A (n_95_77), .B (n_89_80), .C1 (n_86_83), .C2 (n_83_83) );
AOI211_X1 g_101_74 (.ZN (n_101_74), .A (n_97_76), .B (n_91_79), .C1 (n_88_82), .C2 (n_85_82) );
AOI211_X1 g_103_73 (.ZN (n_103_73), .A (n_99_75), .B (n_93_78), .C1 (n_89_80), .C2 (n_84_84) );
AOI211_X1 g_102_75 (.ZN (n_102_75), .A (n_101_74), .B (n_95_77), .C1 (n_91_79), .C2 (n_86_83) );
AOI211_X1 g_104_74 (.ZN (n_104_74), .A (n_103_73), .B (n_97_76), .C1 (n_93_78), .C2 (n_88_82) );
AOI211_X1 g_106_73 (.ZN (n_106_73), .A (n_102_75), .B (n_99_75), .C1 (n_95_77), .C2 (n_89_80) );
AOI211_X1 g_108_72 (.ZN (n_108_72), .A (n_104_74), .B (n_101_74), .C1 (n_97_76), .C2 (n_91_79) );
AOI211_X1 g_110_71 (.ZN (n_110_71), .A (n_106_73), .B (n_103_73), .C1 (n_99_75), .C2 (n_93_78) );
AOI211_X1 g_111_69 (.ZN (n_111_69), .A (n_108_72), .B (n_102_75), .C1 (n_101_74), .C2 (n_95_77) );
AOI211_X1 g_113_68 (.ZN (n_113_68), .A (n_110_71), .B (n_104_74), .C1 (n_103_73), .C2 (n_97_76) );
AOI211_X1 g_115_67 (.ZN (n_115_67), .A (n_111_69), .B (n_106_73), .C1 (n_102_75), .C2 (n_99_75) );
AOI211_X1 g_117_66 (.ZN (n_117_66), .A (n_113_68), .B (n_108_72), .C1 (n_104_74), .C2 (n_101_74) );
AOI211_X1 g_119_65 (.ZN (n_119_65), .A (n_115_67), .B (n_110_71), .C1 (n_106_73), .C2 (n_103_73) );
AOI211_X1 g_121_64 (.ZN (n_121_64), .A (n_117_66), .B (n_111_69), .C1 (n_108_72), .C2 (n_102_75) );
AOI211_X1 g_123_63 (.ZN (n_123_63), .A (n_119_65), .B (n_113_68), .C1 (n_110_71), .C2 (n_104_74) );
AOI211_X1 g_125_62 (.ZN (n_125_62), .A (n_121_64), .B (n_115_67), .C1 (n_111_69), .C2 (n_106_73) );
AOI211_X1 g_127_61 (.ZN (n_127_61), .A (n_123_63), .B (n_117_66), .C1 (n_113_68), .C2 (n_108_72) );
AOI211_X1 g_129_60 (.ZN (n_129_60), .A (n_125_62), .B (n_119_65), .C1 (n_115_67), .C2 (n_110_71) );
AOI211_X1 g_131_59 (.ZN (n_131_59), .A (n_127_61), .B (n_121_64), .C1 (n_117_66), .C2 (n_111_69) );
AOI211_X1 g_133_58 (.ZN (n_133_58), .A (n_129_60), .B (n_123_63), .C1 (n_119_65), .C2 (n_113_68) );
AOI211_X1 g_135_57 (.ZN (n_135_57), .A (n_131_59), .B (n_125_62), .C1 (n_121_64), .C2 (n_115_67) );
AOI211_X1 g_137_56 (.ZN (n_137_56), .A (n_133_58), .B (n_127_61), .C1 (n_123_63), .C2 (n_117_66) );
AOI211_X1 g_139_55 (.ZN (n_139_55), .A (n_135_57), .B (n_129_60), .C1 (n_125_62), .C2 (n_119_65) );
AOI211_X1 g_141_54 (.ZN (n_141_54), .A (n_137_56), .B (n_131_59), .C1 (n_127_61), .C2 (n_121_64) );
AOI211_X1 g_143_53 (.ZN (n_143_53), .A (n_139_55), .B (n_133_58), .C1 (n_129_60), .C2 (n_123_63) );
AOI211_X1 g_145_52 (.ZN (n_145_52), .A (n_141_54), .B (n_135_57), .C1 (n_131_59), .C2 (n_125_62) );
AOI211_X1 g_147_53 (.ZN (n_147_53), .A (n_143_53), .B (n_137_56), .C1 (n_133_58), .C2 (n_127_61) );
AOI211_X1 g_145_54 (.ZN (n_145_54), .A (n_145_52), .B (n_139_55), .C1 (n_135_57), .C2 (n_129_60) );
AOI211_X1 g_143_55 (.ZN (n_143_55), .A (n_147_53), .B (n_141_54), .C1 (n_137_56), .C2 (n_131_59) );
AOI211_X1 g_144_53 (.ZN (n_144_53), .A (n_145_54), .B (n_143_53), .C1 (n_139_55), .C2 (n_133_58) );
AOI211_X1 g_142_54 (.ZN (n_142_54), .A (n_143_55), .B (n_145_52), .C1 (n_141_54), .C2 (n_135_57) );
AOI211_X1 g_140_55 (.ZN (n_140_55), .A (n_144_53), .B (n_147_53), .C1 (n_143_53), .C2 (n_137_56) );
AOI211_X1 g_138_56 (.ZN (n_138_56), .A (n_142_54), .B (n_145_54), .C1 (n_145_52), .C2 (n_139_55) );
AOI211_X1 g_136_57 (.ZN (n_136_57), .A (n_140_55), .B (n_143_55), .C1 (n_147_53), .C2 (n_141_54) );
AOI211_X1 g_134_58 (.ZN (n_134_58), .A (n_138_56), .B (n_144_53), .C1 (n_145_54), .C2 (n_143_53) );
AOI211_X1 g_132_59 (.ZN (n_132_59), .A (n_136_57), .B (n_142_54), .C1 (n_143_55), .C2 (n_145_52) );
AOI211_X1 g_130_60 (.ZN (n_130_60), .A (n_134_58), .B (n_140_55), .C1 (n_144_53), .C2 (n_147_53) );
AOI211_X1 g_128_61 (.ZN (n_128_61), .A (n_132_59), .B (n_138_56), .C1 (n_142_54), .C2 (n_145_54) );
AOI211_X1 g_126_62 (.ZN (n_126_62), .A (n_130_60), .B (n_136_57), .C1 (n_140_55), .C2 (n_143_55) );
AOI211_X1 g_124_63 (.ZN (n_124_63), .A (n_128_61), .B (n_134_58), .C1 (n_138_56), .C2 (n_144_53) );
AOI211_X1 g_122_64 (.ZN (n_122_64), .A (n_126_62), .B (n_132_59), .C1 (n_136_57), .C2 (n_142_54) );
AOI211_X1 g_120_65 (.ZN (n_120_65), .A (n_124_63), .B (n_130_60), .C1 (n_134_58), .C2 (n_140_55) );
AOI211_X1 g_118_66 (.ZN (n_118_66), .A (n_122_64), .B (n_128_61), .C1 (n_132_59), .C2 (n_138_56) );
AOI211_X1 g_116_67 (.ZN (n_116_67), .A (n_120_65), .B (n_126_62), .C1 (n_130_60), .C2 (n_136_57) );
AOI211_X1 g_114_68 (.ZN (n_114_68), .A (n_118_66), .B (n_124_63), .C1 (n_128_61), .C2 (n_134_58) );
AOI211_X1 g_112_69 (.ZN (n_112_69), .A (n_116_67), .B (n_122_64), .C1 (n_126_62), .C2 (n_132_59) );
AOI211_X1 g_110_70 (.ZN (n_110_70), .A (n_114_68), .B (n_120_65), .C1 (n_124_63), .C2 (n_130_60) );
AOI211_X1 g_108_71 (.ZN (n_108_71), .A (n_112_69), .B (n_118_66), .C1 (n_122_64), .C2 (n_128_61) );
AOI211_X1 g_106_72 (.ZN (n_106_72), .A (n_110_70), .B (n_116_67), .C1 (n_120_65), .C2 (n_126_62) );
AOI211_X1 g_104_73 (.ZN (n_104_73), .A (n_108_71), .B (n_114_68), .C1 (n_118_66), .C2 (n_124_63) );
AOI211_X1 g_102_74 (.ZN (n_102_74), .A (n_106_72), .B (n_112_69), .C1 (n_116_67), .C2 (n_122_64) );
AOI211_X1 g_100_75 (.ZN (n_100_75), .A (n_104_73), .B (n_110_70), .C1 (n_114_68), .C2 (n_120_65) );
AOI211_X1 g_98_76 (.ZN (n_98_76), .A (n_102_74), .B (n_108_71), .C1 (n_112_69), .C2 (n_118_66) );
AOI211_X1 g_96_77 (.ZN (n_96_77), .A (n_100_75), .B (n_106_72), .C1 (n_110_70), .C2 (n_116_67) );
AOI211_X1 g_95_79 (.ZN (n_95_79), .A (n_98_76), .B (n_104_73), .C1 (n_108_71), .C2 (n_114_68) );
AOI211_X1 g_97_78 (.ZN (n_97_78), .A (n_96_77), .B (n_102_74), .C1 (n_106_72), .C2 (n_112_69) );
AOI211_X1 g_99_77 (.ZN (n_99_77), .A (n_95_79), .B (n_100_75), .C1 (n_104_73), .C2 (n_110_70) );
AOI211_X1 g_101_76 (.ZN (n_101_76), .A (n_97_78), .B (n_98_76), .C1 (n_102_74), .C2 (n_108_71) );
AOI211_X1 g_103_75 (.ZN (n_103_75), .A (n_99_77), .B (n_96_77), .C1 (n_100_75), .C2 (n_106_72) );
AOI211_X1 g_105_74 (.ZN (n_105_74), .A (n_101_76), .B (n_95_79), .C1 (n_98_76), .C2 (n_104_73) );
AOI211_X1 g_107_73 (.ZN (n_107_73), .A (n_103_75), .B (n_97_78), .C1 (n_96_77), .C2 (n_102_74) );
AOI211_X1 g_109_72 (.ZN (n_109_72), .A (n_105_74), .B (n_99_77), .C1 (n_95_79), .C2 (n_100_75) );
AOI211_X1 g_111_71 (.ZN (n_111_71), .A (n_107_73), .B (n_101_76), .C1 (n_97_78), .C2 (n_98_76) );
AOI211_X1 g_113_70 (.ZN (n_113_70), .A (n_109_72), .B (n_103_75), .C1 (n_99_77), .C2 (n_96_77) );
AOI211_X1 g_115_69 (.ZN (n_115_69), .A (n_111_71), .B (n_105_74), .C1 (n_101_76), .C2 (n_95_79) );
AOI211_X1 g_117_68 (.ZN (n_117_68), .A (n_113_70), .B (n_107_73), .C1 (n_103_75), .C2 (n_97_78) );
AOI211_X1 g_119_67 (.ZN (n_119_67), .A (n_115_69), .B (n_109_72), .C1 (n_105_74), .C2 (n_99_77) );
AOI211_X1 g_121_66 (.ZN (n_121_66), .A (n_117_68), .B (n_111_71), .C1 (n_107_73), .C2 (n_101_76) );
AOI211_X1 g_123_65 (.ZN (n_123_65), .A (n_119_67), .B (n_113_70), .C1 (n_109_72), .C2 (n_103_75) );
AOI211_X1 g_125_64 (.ZN (n_125_64), .A (n_121_66), .B (n_115_69), .C1 (n_111_71), .C2 (n_105_74) );
AOI211_X1 g_127_63 (.ZN (n_127_63), .A (n_123_65), .B (n_117_68), .C1 (n_113_70), .C2 (n_107_73) );
AOI211_X1 g_129_62 (.ZN (n_129_62), .A (n_125_64), .B (n_119_67), .C1 (n_115_69), .C2 (n_109_72) );
AOI211_X1 g_131_61 (.ZN (n_131_61), .A (n_127_63), .B (n_121_66), .C1 (n_117_68), .C2 (n_111_71) );
AOI211_X1 g_133_60 (.ZN (n_133_60), .A (n_129_62), .B (n_123_65), .C1 (n_119_67), .C2 (n_113_70) );
AOI211_X1 g_135_59 (.ZN (n_135_59), .A (n_131_61), .B (n_125_64), .C1 (n_121_66), .C2 (n_115_69) );
AOI211_X1 g_137_58 (.ZN (n_137_58), .A (n_133_60), .B (n_127_63), .C1 (n_123_65), .C2 (n_117_68) );
AOI211_X1 g_139_57 (.ZN (n_139_57), .A (n_135_59), .B (n_129_62), .C1 (n_125_64), .C2 (n_119_67) );
AOI211_X1 g_141_56 (.ZN (n_141_56), .A (n_137_58), .B (n_131_61), .C1 (n_127_63), .C2 (n_121_66) );
AOI211_X1 g_140_58 (.ZN (n_140_58), .A (n_139_57), .B (n_133_60), .C1 (n_129_62), .C2 (n_123_65) );
AOI211_X1 g_139_56 (.ZN (n_139_56), .A (n_141_56), .B (n_135_59), .C1 (n_131_61), .C2 (n_125_64) );
AOI211_X1 g_141_55 (.ZN (n_141_55), .A (n_140_58), .B (n_137_58), .C1 (n_133_60), .C2 (n_127_63) );
AOI211_X1 g_143_54 (.ZN (n_143_54), .A (n_139_56), .B (n_139_57), .C1 (n_135_59), .C2 (n_129_62) );
AOI211_X1 g_145_55 (.ZN (n_145_55), .A (n_141_55), .B (n_141_56), .C1 (n_137_58), .C2 (n_131_61) );
AOI211_X1 g_147_56 (.ZN (n_147_56), .A (n_143_54), .B (n_140_58), .C1 (n_139_57), .C2 (n_133_60) );
AOI211_X1 g_146_54 (.ZN (n_146_54), .A (n_145_55), .B (n_139_56), .C1 (n_141_56), .C2 (n_135_59) );
AOI211_X1 g_148_55 (.ZN (n_148_55), .A (n_147_56), .B (n_141_55), .C1 (n_140_58), .C2 (n_137_58) );
AOI211_X1 g_149_57 (.ZN (n_149_57), .A (n_146_54), .B (n_143_54), .C1 (n_139_56), .C2 (n_139_57) );
AOI211_X1 g_147_58 (.ZN (n_147_58), .A (n_148_55), .B (n_145_55), .C1 (n_141_55), .C2 (n_141_56) );
AOI211_X1 g_146_56 (.ZN (n_146_56), .A (n_149_57), .B (n_147_56), .C1 (n_143_54), .C2 (n_140_58) );
AOI211_X1 g_144_55 (.ZN (n_144_55), .A (n_147_58), .B (n_146_54), .C1 (n_145_55), .C2 (n_139_56) );
AOI211_X1 g_142_56 (.ZN (n_142_56), .A (n_146_56), .B (n_148_55), .C1 (n_147_56), .C2 (n_141_55) );
AOI211_X1 g_140_57 (.ZN (n_140_57), .A (n_144_55), .B (n_149_57), .C1 (n_146_54), .C2 (n_143_54) );
AOI211_X1 g_138_58 (.ZN (n_138_58), .A (n_142_56), .B (n_147_58), .C1 (n_148_55), .C2 (n_145_55) );
AOI211_X1 g_136_59 (.ZN (n_136_59), .A (n_140_57), .B (n_146_56), .C1 (n_149_57), .C2 (n_147_56) );
AOI211_X1 g_137_57 (.ZN (n_137_57), .A (n_138_58), .B (n_144_55), .C1 (n_147_58), .C2 (n_146_54) );
AOI211_X1 g_135_58 (.ZN (n_135_58), .A (n_136_59), .B (n_142_56), .C1 (n_146_56), .C2 (n_148_55) );
AOI211_X1 g_133_59 (.ZN (n_133_59), .A (n_137_57), .B (n_140_57), .C1 (n_144_55), .C2 (n_149_57) );
AOI211_X1 g_132_61 (.ZN (n_132_61), .A (n_135_58), .B (n_138_58), .C1 (n_142_56), .C2 (n_147_58) );
AOI211_X1 g_134_60 (.ZN (n_134_60), .A (n_133_59), .B (n_136_59), .C1 (n_140_57), .C2 (n_146_56) );
AOI211_X1 g_133_62 (.ZN (n_133_62), .A (n_132_61), .B (n_137_57), .C1 (n_138_58), .C2 (n_144_55) );
AOI211_X1 g_132_60 (.ZN (n_132_60), .A (n_134_60), .B (n_135_58), .C1 (n_136_59), .C2 (n_142_56) );
AOI211_X1 g_134_59 (.ZN (n_134_59), .A (n_133_62), .B (n_133_59), .C1 (n_137_57), .C2 (n_140_57) );
AOI211_X1 g_136_58 (.ZN (n_136_58), .A (n_132_60), .B (n_132_61), .C1 (n_135_58), .C2 (n_138_58) );
AOI211_X1 g_138_57 (.ZN (n_138_57), .A (n_134_59), .B (n_134_60), .C1 (n_133_59), .C2 (n_136_59) );
AOI211_X1 g_140_56 (.ZN (n_140_56), .A (n_136_58), .B (n_133_62), .C1 (n_132_61), .C2 (n_137_57) );
AOI211_X1 g_142_55 (.ZN (n_142_55), .A (n_138_57), .B (n_132_60), .C1 (n_134_60), .C2 (n_135_58) );
AOI211_X1 g_144_54 (.ZN (n_144_54), .A (n_140_56), .B (n_134_59), .C1 (n_133_62), .C2 (n_133_59) );
AOI211_X1 g_146_55 (.ZN (n_146_55), .A (n_142_55), .B (n_136_58), .C1 (n_132_60), .C2 (n_132_61) );
AOI211_X1 g_144_56 (.ZN (n_144_56), .A (n_144_54), .B (n_138_57), .C1 (n_134_59), .C2 (n_134_60) );
AOI211_X1 g_142_57 (.ZN (n_142_57), .A (n_146_55), .B (n_140_56), .C1 (n_136_58), .C2 (n_133_62) );
AOI211_X1 g_141_59 (.ZN (n_141_59), .A (n_144_56), .B (n_142_55), .C1 (n_138_57), .C2 (n_132_60) );
AOI211_X1 g_139_58 (.ZN (n_139_58), .A (n_142_57), .B (n_144_54), .C1 (n_140_56), .C2 (n_134_59) );
AOI211_X1 g_141_57 (.ZN (n_141_57), .A (n_141_59), .B (n_146_55), .C1 (n_142_55), .C2 (n_136_58) );
AOI211_X1 g_143_56 (.ZN (n_143_56), .A (n_139_58), .B (n_144_56), .C1 (n_144_54), .C2 (n_138_57) );
AOI211_X1 g_145_57 (.ZN (n_145_57), .A (n_141_57), .B (n_142_57), .C1 (n_146_55), .C2 (n_140_56) );
AOI211_X1 g_143_58 (.ZN (n_143_58), .A (n_143_56), .B (n_141_59), .C1 (n_144_56), .C2 (n_142_55) );
AOI211_X1 g_145_59 (.ZN (n_145_59), .A (n_145_57), .B (n_139_58), .C1 (n_142_57), .C2 (n_144_54) );
AOI211_X1 g_144_57 (.ZN (n_144_57), .A (n_143_58), .B (n_141_57), .C1 (n_141_59), .C2 (n_146_55) );
AOI211_X1 g_142_58 (.ZN (n_142_58), .A (n_145_59), .B (n_143_56), .C1 (n_139_58), .C2 (n_144_56) );
AOI211_X1 g_140_59 (.ZN (n_140_59), .A (n_144_57), .B (n_145_57), .C1 (n_141_57), .C2 (n_142_57) );
AOI211_X1 g_138_60 (.ZN (n_138_60), .A (n_142_58), .B (n_143_58), .C1 (n_143_56), .C2 (n_141_59) );
AOI211_X1 g_136_61 (.ZN (n_136_61), .A (n_140_59), .B (n_145_59), .C1 (n_145_57), .C2 (n_139_58) );
AOI211_X1 g_137_59 (.ZN (n_137_59), .A (n_138_60), .B (n_144_57), .C1 (n_143_58), .C2 (n_141_57) );
AOI211_X1 g_135_60 (.ZN (n_135_60), .A (n_136_61), .B (n_142_58), .C1 (n_145_59), .C2 (n_143_56) );
AOI211_X1 g_133_61 (.ZN (n_133_61), .A (n_137_59), .B (n_140_59), .C1 (n_144_57), .C2 (n_145_57) );
AOI211_X1 g_131_62 (.ZN (n_131_62), .A (n_135_60), .B (n_138_60), .C1 (n_142_58), .C2 (n_143_58) );
AOI211_X1 g_129_63 (.ZN (n_129_63), .A (n_133_61), .B (n_136_61), .C1 (n_140_59), .C2 (n_145_59) );
AOI211_X1 g_130_61 (.ZN (n_130_61), .A (n_131_62), .B (n_137_59), .C1 (n_138_60), .C2 (n_144_57) );
AOI211_X1 g_128_62 (.ZN (n_128_62), .A (n_129_63), .B (n_135_60), .C1 (n_136_61), .C2 (n_142_58) );
AOI211_X1 g_126_63 (.ZN (n_126_63), .A (n_130_61), .B (n_133_61), .C1 (n_137_59), .C2 (n_140_59) );
AOI211_X1 g_124_64 (.ZN (n_124_64), .A (n_128_62), .B (n_131_62), .C1 (n_135_60), .C2 (n_138_60) );
AOI211_X1 g_122_65 (.ZN (n_122_65), .A (n_126_63), .B (n_129_63), .C1 (n_133_61), .C2 (n_136_61) );
AOI211_X1 g_120_66 (.ZN (n_120_66), .A (n_124_64), .B (n_130_61), .C1 (n_131_62), .C2 (n_137_59) );
AOI211_X1 g_118_67 (.ZN (n_118_67), .A (n_122_65), .B (n_128_62), .C1 (n_129_63), .C2 (n_135_60) );
AOI211_X1 g_116_68 (.ZN (n_116_68), .A (n_120_66), .B (n_126_63), .C1 (n_130_61), .C2 (n_133_61) );
AOI211_X1 g_114_69 (.ZN (n_114_69), .A (n_118_67), .B (n_124_64), .C1 (n_128_62), .C2 (n_131_62) );
AOI211_X1 g_112_70 (.ZN (n_112_70), .A (n_116_68), .B (n_122_65), .C1 (n_126_63), .C2 (n_129_63) );
AOI211_X1 g_111_72 (.ZN (n_111_72), .A (n_114_69), .B (n_120_66), .C1 (n_124_64), .C2 (n_130_61) );
AOI211_X1 g_113_71 (.ZN (n_113_71), .A (n_112_70), .B (n_118_67), .C1 (n_122_65), .C2 (n_128_62) );
AOI211_X1 g_115_70 (.ZN (n_115_70), .A (n_111_72), .B (n_116_68), .C1 (n_120_66), .C2 (n_126_63) );
AOI211_X1 g_117_69 (.ZN (n_117_69), .A (n_113_71), .B (n_114_69), .C1 (n_118_67), .C2 (n_124_64) );
AOI211_X1 g_119_68 (.ZN (n_119_68), .A (n_115_70), .B (n_112_70), .C1 (n_116_68), .C2 (n_122_65) );
AOI211_X1 g_121_67 (.ZN (n_121_67), .A (n_117_69), .B (n_111_72), .C1 (n_114_69), .C2 (n_120_66) );
AOI211_X1 g_123_66 (.ZN (n_123_66), .A (n_119_68), .B (n_113_71), .C1 (n_112_70), .C2 (n_118_67) );
AOI211_X1 g_125_65 (.ZN (n_125_65), .A (n_121_67), .B (n_115_70), .C1 (n_111_72), .C2 (n_116_68) );
AOI211_X1 g_127_64 (.ZN (n_127_64), .A (n_123_66), .B (n_117_69), .C1 (n_113_71), .C2 (n_114_69) );
AOI211_X1 g_126_66 (.ZN (n_126_66), .A (n_125_65), .B (n_119_68), .C1 (n_115_70), .C2 (n_112_70) );
AOI211_X1 g_124_65 (.ZN (n_124_65), .A (n_127_64), .B (n_121_67), .C1 (n_117_69), .C2 (n_111_72) );
AOI211_X1 g_126_64 (.ZN (n_126_64), .A (n_126_66), .B (n_123_66), .C1 (n_119_68), .C2 (n_113_71) );
AOI211_X1 g_128_63 (.ZN (n_128_63), .A (n_124_65), .B (n_125_65), .C1 (n_121_67), .C2 (n_115_70) );
AOI211_X1 g_130_62 (.ZN (n_130_62), .A (n_126_64), .B (n_127_64), .C1 (n_123_66), .C2 (n_117_69) );
AOI211_X1 g_129_64 (.ZN (n_129_64), .A (n_128_63), .B (n_126_66), .C1 (n_125_65), .C2 (n_119_68) );
AOI211_X1 g_131_63 (.ZN (n_131_63), .A (n_130_62), .B (n_124_65), .C1 (n_127_64), .C2 (n_121_67) );
AOI211_X1 g_130_65 (.ZN (n_130_65), .A (n_129_64), .B (n_126_64), .C1 (n_126_66), .C2 (n_123_66) );
AOI211_X1 g_128_64 (.ZN (n_128_64), .A (n_131_63), .B (n_128_63), .C1 (n_124_65), .C2 (n_125_65) );
AOI211_X1 g_130_63 (.ZN (n_130_63), .A (n_130_65), .B (n_130_62), .C1 (n_126_64), .C2 (n_127_64) );
AOI211_X1 g_132_62 (.ZN (n_132_62), .A (n_128_64), .B (n_129_64), .C1 (n_128_63), .C2 (n_126_66) );
AOI211_X1 g_134_61 (.ZN (n_134_61), .A (n_130_63), .B (n_131_63), .C1 (n_130_62), .C2 (n_124_65) );
AOI211_X1 g_136_60 (.ZN (n_136_60), .A (n_132_62), .B (n_130_65), .C1 (n_129_64), .C2 (n_126_64) );
AOI211_X1 g_138_59 (.ZN (n_138_59), .A (n_134_61), .B (n_128_64), .C1 (n_131_63), .C2 (n_128_63) );
AOI211_X1 g_137_61 (.ZN (n_137_61), .A (n_136_60), .B (n_130_63), .C1 (n_130_65), .C2 (n_130_62) );
AOI211_X1 g_139_60 (.ZN (n_139_60), .A (n_138_59), .B (n_132_62), .C1 (n_128_64), .C2 (n_129_64) );
AOI211_X1 g_138_62 (.ZN (n_138_62), .A (n_137_61), .B (n_134_61), .C1 (n_130_63), .C2 (n_131_63) );
AOI211_X1 g_137_60 (.ZN (n_137_60), .A (n_139_60), .B (n_136_60), .C1 (n_132_62), .C2 (n_130_65) );
AOI211_X1 g_135_61 (.ZN (n_135_61), .A (n_138_62), .B (n_138_59), .C1 (n_134_61), .C2 (n_128_64) );
AOI211_X1 g_134_63 (.ZN (n_134_63), .A (n_137_60), .B (n_137_61), .C1 (n_136_60), .C2 (n_130_63) );
AOI211_X1 g_132_64 (.ZN (n_132_64), .A (n_135_61), .B (n_139_60), .C1 (n_138_59), .C2 (n_132_62) );
AOI211_X1 g_131_66 (.ZN (n_131_66), .A (n_134_63), .B (n_138_62), .C1 (n_137_61), .C2 (n_134_61) );
AOI211_X1 g_130_64 (.ZN (n_130_64), .A (n_132_64), .B (n_137_60), .C1 (n_139_60), .C2 (n_136_60) );
AOI211_X1 g_128_65 (.ZN (n_128_65), .A (n_131_66), .B (n_135_61), .C1 (n_138_62), .C2 (n_138_59) );
AOI211_X1 g_129_67 (.ZN (n_129_67), .A (n_130_64), .B (n_134_63), .C1 (n_137_60), .C2 (n_137_61) );
AOI211_X1 g_127_66 (.ZN (n_127_66), .A (n_128_65), .B (n_132_64), .C1 (n_135_61), .C2 (n_139_60) );
AOI211_X1 g_129_65 (.ZN (n_129_65), .A (n_129_67), .B (n_131_66), .C1 (n_134_63), .C2 (n_138_62) );
AOI211_X1 g_131_64 (.ZN (n_131_64), .A (n_127_66), .B (n_130_64), .C1 (n_132_64), .C2 (n_137_60) );
AOI211_X1 g_133_63 (.ZN (n_133_63), .A (n_129_65), .B (n_128_65), .C1 (n_131_66), .C2 (n_135_61) );
AOI211_X1 g_135_62 (.ZN (n_135_62), .A (n_131_64), .B (n_129_67), .C1 (n_130_64), .C2 (n_134_63) );
AOI211_X1 g_134_64 (.ZN (n_134_64), .A (n_133_63), .B (n_127_66), .C1 (n_128_65), .C2 (n_132_64) );
AOI211_X1 g_132_63 (.ZN (n_132_63), .A (n_135_62), .B (n_129_65), .C1 (n_129_67), .C2 (n_131_66) );
AOI211_X1 g_134_62 (.ZN (n_134_62), .A (n_134_64), .B (n_131_64), .C1 (n_127_66), .C2 (n_130_64) );
AOI211_X1 g_136_63 (.ZN (n_136_63), .A (n_132_63), .B (n_133_63), .C1 (n_129_65), .C2 (n_128_65) );
AOI211_X1 g_135_65 (.ZN (n_135_65), .A (n_134_62), .B (n_135_62), .C1 (n_131_64), .C2 (n_129_67) );
AOI211_X1 g_133_64 (.ZN (n_133_64), .A (n_136_63), .B (n_134_64), .C1 (n_133_63), .C2 (n_127_66) );
AOI211_X1 g_135_63 (.ZN (n_135_63), .A (n_135_65), .B (n_132_63), .C1 (n_135_62), .C2 (n_129_65) );
AOI211_X1 g_137_62 (.ZN (n_137_62), .A (n_133_64), .B (n_134_62), .C1 (n_134_64), .C2 (n_131_64) );
AOI211_X1 g_139_61 (.ZN (n_139_61), .A (n_135_63), .B (n_136_63), .C1 (n_132_63), .C2 (n_133_63) );
AOI211_X1 g_141_60 (.ZN (n_141_60), .A (n_137_62), .B (n_135_65), .C1 (n_134_62), .C2 (n_135_62) );
AOI211_X1 g_139_59 (.ZN (n_139_59), .A (n_139_61), .B (n_133_64), .C1 (n_136_63), .C2 (n_134_64) );
AOI211_X1 g_141_58 (.ZN (n_141_58), .A (n_141_60), .B (n_135_63), .C1 (n_135_65), .C2 (n_132_63) );
AOI211_X1 g_143_57 (.ZN (n_143_57), .A (n_139_59), .B (n_137_62), .C1 (n_133_64), .C2 (n_134_62) );
AOI211_X1 g_145_56 (.ZN (n_145_56), .A (n_141_58), .B (n_139_61), .C1 (n_135_63), .C2 (n_136_63) );
AOI211_X1 g_147_57 (.ZN (n_147_57), .A (n_143_57), .B (n_141_60), .C1 (n_137_62), .C2 (n_135_65) );
AOI211_X1 g_145_58 (.ZN (n_145_58), .A (n_145_56), .B (n_139_59), .C1 (n_139_61), .C2 (n_133_64) );
AOI211_X1 g_143_59 (.ZN (n_143_59), .A (n_147_57), .B (n_141_58), .C1 (n_141_60), .C2 (n_135_63) );
AOI211_X1 g_142_61 (.ZN (n_142_61), .A (n_145_58), .B (n_143_57), .C1 (n_139_59), .C2 (n_137_62) );
AOI211_X1 g_144_60 (.ZN (n_144_60), .A (n_143_59), .B (n_145_56), .C1 (n_141_58), .C2 (n_139_61) );
AOI211_X1 g_146_59 (.ZN (n_146_59), .A (n_142_61), .B (n_147_57), .C1 (n_143_57), .C2 (n_141_60) );
AOI211_X1 g_144_58 (.ZN (n_144_58), .A (n_144_60), .B (n_145_58), .C1 (n_145_56), .C2 (n_139_59) );
AOI211_X1 g_142_59 (.ZN (n_142_59), .A (n_146_59), .B (n_143_59), .C1 (n_147_57), .C2 (n_141_58) );
AOI211_X1 g_140_60 (.ZN (n_140_60), .A (n_144_58), .B (n_142_61), .C1 (n_145_58), .C2 (n_143_57) );
AOI211_X1 g_138_61 (.ZN (n_138_61), .A (n_142_59), .B (n_144_60), .C1 (n_143_59), .C2 (n_145_56) );
AOI211_X1 g_136_62 (.ZN (n_136_62), .A (n_140_60), .B (n_146_59), .C1 (n_142_61), .C2 (n_147_57) );
AOI211_X1 g_137_64 (.ZN (n_137_64), .A (n_138_61), .B (n_144_58), .C1 (n_144_60), .C2 (n_145_58) );
AOI211_X1 g_139_63 (.ZN (n_139_63), .A (n_136_62), .B (n_142_59), .C1 (n_146_59), .C2 (n_143_59) );
AOI211_X1 g_140_61 (.ZN (n_140_61), .A (n_137_64), .B (n_140_60), .C1 (n_144_58), .C2 (n_142_61) );
AOI211_X1 g_142_60 (.ZN (n_142_60), .A (n_139_63), .B (n_138_61), .C1 (n_142_59), .C2 (n_144_60) );
AOI211_X1 g_144_59 (.ZN (n_144_59), .A (n_140_61), .B (n_136_62), .C1 (n_140_60), .C2 (n_146_59) );
AOI211_X1 g_146_58 (.ZN (n_146_58), .A (n_142_60), .B (n_137_64), .C1 (n_138_61), .C2 (n_144_58) );
AOI211_X1 g_147_60 (.ZN (n_147_60), .A (n_144_59), .B (n_139_63), .C1 (n_136_62), .C2 (n_142_59) );
AOI211_X1 g_149_61 (.ZN (n_149_61), .A (n_146_58), .B (n_140_61), .C1 (n_137_64), .C2 (n_140_60) );
AOI211_X1 g_148_59 (.ZN (n_148_59), .A (n_147_60), .B (n_142_60), .C1 (n_139_63), .C2 (n_138_61) );
AOI211_X1 g_146_60 (.ZN (n_146_60), .A (n_149_61), .B (n_144_59), .C1 (n_140_61), .C2 (n_136_62) );
AOI211_X1 g_147_62 (.ZN (n_147_62), .A (n_148_59), .B (n_146_58), .C1 (n_142_60), .C2 (n_137_64) );
AOI211_X1 g_145_61 (.ZN (n_145_61), .A (n_146_60), .B (n_147_60), .C1 (n_144_59), .C2 (n_139_63) );
AOI211_X1 g_143_60 (.ZN (n_143_60), .A (n_147_62), .B (n_149_61), .C1 (n_146_58), .C2 (n_140_61) );
AOI211_X1 g_141_61 (.ZN (n_141_61), .A (n_145_61), .B (n_148_59), .C1 (n_147_60), .C2 (n_142_60) );
AOI211_X1 g_139_62 (.ZN (n_139_62), .A (n_143_60), .B (n_146_60), .C1 (n_149_61), .C2 (n_144_59) );
AOI211_X1 g_137_63 (.ZN (n_137_63), .A (n_141_61), .B (n_147_62), .C1 (n_148_59), .C2 (n_146_58) );
AOI211_X1 g_135_64 (.ZN (n_135_64), .A (n_139_62), .B (n_145_61), .C1 (n_146_60), .C2 (n_147_60) );
AOI211_X1 g_133_65 (.ZN (n_133_65), .A (n_137_63), .B (n_143_60), .C1 (n_147_62), .C2 (n_149_61) );
AOI211_X1 g_134_67 (.ZN (n_134_67), .A (n_135_64), .B (n_141_61), .C1 (n_145_61), .C2 (n_148_59) );
AOI211_X1 g_132_66 (.ZN (n_132_66), .A (n_133_65), .B (n_139_62), .C1 (n_143_60), .C2 (n_146_60) );
AOI211_X1 g_134_65 (.ZN (n_134_65), .A (n_134_67), .B (n_137_63), .C1 (n_141_61), .C2 (n_147_62) );
AOI211_X1 g_136_64 (.ZN (n_136_64), .A (n_132_66), .B (n_135_64), .C1 (n_139_62), .C2 (n_145_61) );
AOI211_X1 g_138_63 (.ZN (n_138_63), .A (n_134_65), .B (n_133_65), .C1 (n_137_63), .C2 (n_143_60) );
AOI211_X1 g_140_62 (.ZN (n_140_62), .A (n_136_64), .B (n_134_67), .C1 (n_135_64), .C2 (n_141_61) );
AOI211_X1 g_139_64 (.ZN (n_139_64), .A (n_138_63), .B (n_132_66), .C1 (n_133_65), .C2 (n_139_62) );
AOI211_X1 g_141_63 (.ZN (n_141_63), .A (n_140_62), .B (n_134_65), .C1 (n_134_67), .C2 (n_137_63) );
AOI211_X1 g_143_62 (.ZN (n_143_62), .A (n_139_64), .B (n_136_64), .C1 (n_132_66), .C2 (n_135_64) );
AOI211_X1 g_145_63 (.ZN (n_145_63), .A (n_141_63), .B (n_138_63), .C1 (n_134_65), .C2 (n_133_65) );
AOI211_X1 g_144_61 (.ZN (n_144_61), .A (n_143_62), .B (n_140_62), .C1 (n_136_64), .C2 (n_134_67) );
AOI211_X1 g_142_62 (.ZN (n_142_62), .A (n_145_63), .B (n_139_64), .C1 (n_138_63), .C2 (n_132_66) );
AOI211_X1 g_140_63 (.ZN (n_140_63), .A (n_144_61), .B (n_141_63), .C1 (n_140_62), .C2 (n_134_65) );
AOI211_X1 g_138_64 (.ZN (n_138_64), .A (n_142_62), .B (n_143_62), .C1 (n_139_64), .C2 (n_136_64) );
AOI211_X1 g_136_65 (.ZN (n_136_65), .A (n_140_63), .B (n_145_63), .C1 (n_141_63), .C2 (n_138_63) );
AOI211_X1 g_134_66 (.ZN (n_134_66), .A (n_138_64), .B (n_144_61), .C1 (n_143_62), .C2 (n_140_62) );
AOI211_X1 g_132_65 (.ZN (n_132_65), .A (n_136_65), .B (n_142_62), .C1 (n_145_63), .C2 (n_139_64) );
AOI211_X1 g_130_66 (.ZN (n_130_66), .A (n_134_66), .B (n_140_63), .C1 (n_144_61), .C2 (n_141_63) );
AOI211_X1 g_128_67 (.ZN (n_128_67), .A (n_132_65), .B (n_138_64), .C1 (n_142_62), .C2 (n_143_62) );
AOI211_X1 g_127_65 (.ZN (n_127_65), .A (n_130_66), .B (n_136_65), .C1 (n_140_63), .C2 (n_145_63) );
AOI211_X1 g_125_66 (.ZN (n_125_66), .A (n_128_67), .B (n_134_66), .C1 (n_138_64), .C2 (n_144_61) );
AOI211_X1 g_123_67 (.ZN (n_123_67), .A (n_127_65), .B (n_132_65), .C1 (n_136_65), .C2 (n_142_62) );
AOI211_X1 g_121_68 (.ZN (n_121_68), .A (n_125_66), .B (n_130_66), .C1 (n_134_66), .C2 (n_140_63) );
AOI211_X1 g_122_66 (.ZN (n_122_66), .A (n_123_67), .B (n_128_67), .C1 (n_132_65), .C2 (n_138_64) );
AOI211_X1 g_120_67 (.ZN (n_120_67), .A (n_121_68), .B (n_127_65), .C1 (n_130_66), .C2 (n_136_65) );
AOI211_X1 g_118_68 (.ZN (n_118_68), .A (n_122_66), .B (n_125_66), .C1 (n_128_67), .C2 (n_134_66) );
AOI211_X1 g_116_69 (.ZN (n_116_69), .A (n_120_67), .B (n_123_67), .C1 (n_127_65), .C2 (n_132_65) );
AOI211_X1 g_114_70 (.ZN (n_114_70), .A (n_118_68), .B (n_121_68), .C1 (n_125_66), .C2 (n_130_66) );
AOI211_X1 g_112_71 (.ZN (n_112_71), .A (n_116_69), .B (n_122_66), .C1 (n_123_67), .C2 (n_128_67) );
AOI211_X1 g_110_72 (.ZN (n_110_72), .A (n_114_70), .B (n_120_67), .C1 (n_121_68), .C2 (n_127_65) );
AOI211_X1 g_108_73 (.ZN (n_108_73), .A (n_112_71), .B (n_118_68), .C1 (n_122_66), .C2 (n_125_66) );
AOI211_X1 g_106_74 (.ZN (n_106_74), .A (n_110_72), .B (n_116_69), .C1 (n_120_67), .C2 (n_123_67) );
AOI211_X1 g_104_75 (.ZN (n_104_75), .A (n_108_73), .B (n_114_70), .C1 (n_118_68), .C2 (n_121_68) );
AOI211_X1 g_102_76 (.ZN (n_102_76), .A (n_106_74), .B (n_112_71), .C1 (n_116_69), .C2 (n_122_66) );
AOI211_X1 g_100_77 (.ZN (n_100_77), .A (n_104_75), .B (n_110_72), .C1 (n_114_70), .C2 (n_120_67) );
AOI211_X1 g_98_78 (.ZN (n_98_78), .A (n_102_76), .B (n_108_73), .C1 (n_112_71), .C2 (n_118_68) );
AOI211_X1 g_96_79 (.ZN (n_96_79), .A (n_100_77), .B (n_106_74), .C1 (n_110_72), .C2 (n_116_69) );
AOI211_X1 g_94_80 (.ZN (n_94_80), .A (n_98_78), .B (n_104_75), .C1 (n_108_73), .C2 (n_114_70) );
AOI211_X1 g_92_81 (.ZN (n_92_81), .A (n_96_79), .B (n_102_76), .C1 (n_106_74), .C2 (n_112_71) );
AOI211_X1 g_90_82 (.ZN (n_90_82), .A (n_94_80), .B (n_100_77), .C1 (n_104_75), .C2 (n_110_72) );
AOI211_X1 g_88_83 (.ZN (n_88_83), .A (n_92_81), .B (n_98_78), .C1 (n_102_76), .C2 (n_108_73) );
AOI211_X1 g_86_82 (.ZN (n_86_82), .A (n_90_82), .B (n_96_79), .C1 (n_100_77), .C2 (n_106_74) );
AOI211_X1 g_84_83 (.ZN (n_84_83), .A (n_88_83), .B (n_94_80), .C1 (n_98_78), .C2 (n_104_75) );
AOI211_X1 g_82_84 (.ZN (n_82_84), .A (n_86_82), .B (n_92_81), .C1 (n_96_79), .C2 (n_102_76) );
AOI211_X1 g_80_85 (.ZN (n_80_85), .A (n_84_83), .B (n_90_82), .C1 (n_94_80), .C2 (n_100_77) );
AOI211_X1 g_78_86 (.ZN (n_78_86), .A (n_82_84), .B (n_88_83), .C1 (n_92_81), .C2 (n_98_78) );
AOI211_X1 g_76_87 (.ZN (n_76_87), .A (n_80_85), .B (n_86_82), .C1 (n_90_82), .C2 (n_96_79) );
AOI211_X1 g_74_88 (.ZN (n_74_88), .A (n_78_86), .B (n_84_83), .C1 (n_88_83), .C2 (n_94_80) );
AOI211_X1 g_72_87 (.ZN (n_72_87), .A (n_76_87), .B (n_82_84), .C1 (n_86_82), .C2 (n_92_81) );
AOI211_X1 g_70_88 (.ZN (n_70_88), .A (n_74_88), .B (n_80_85), .C1 (n_84_83), .C2 (n_90_82) );
AOI211_X1 g_68_89 (.ZN (n_68_89), .A (n_72_87), .B (n_78_86), .C1 (n_82_84), .C2 (n_88_83) );
AOI211_X1 g_66_90 (.ZN (n_66_90), .A (n_70_88), .B (n_76_87), .C1 (n_80_85), .C2 (n_86_82) );
AOI211_X1 g_64_91 (.ZN (n_64_91), .A (n_68_89), .B (n_74_88), .C1 (n_78_86), .C2 (n_84_83) );
AOI211_X1 g_62_92 (.ZN (n_62_92), .A (n_66_90), .B (n_72_87), .C1 (n_76_87), .C2 (n_82_84) );
AOI211_X1 g_60_93 (.ZN (n_60_93), .A (n_64_91), .B (n_70_88), .C1 (n_74_88), .C2 (n_80_85) );
AOI211_X1 g_58_94 (.ZN (n_58_94), .A (n_62_92), .B (n_68_89), .C1 (n_72_87), .C2 (n_78_86) );
AOI211_X1 g_56_95 (.ZN (n_56_95), .A (n_60_93), .B (n_66_90), .C1 (n_70_88), .C2 (n_76_87) );
AOI211_X1 g_54_96 (.ZN (n_54_96), .A (n_58_94), .B (n_64_91), .C1 (n_68_89), .C2 (n_74_88) );
AOI211_X1 g_52_97 (.ZN (n_52_97), .A (n_56_95), .B (n_62_92), .C1 (n_66_90), .C2 (n_72_87) );
AOI211_X1 g_51_99 (.ZN (n_51_99), .A (n_54_96), .B (n_60_93), .C1 (n_64_91), .C2 (n_70_88) );
AOI211_X1 g_53_98 (.ZN (n_53_98), .A (n_52_97), .B (n_58_94), .C1 (n_62_92), .C2 (n_68_89) );
AOI211_X1 g_55_97 (.ZN (n_55_97), .A (n_51_99), .B (n_56_95), .C1 (n_60_93), .C2 (n_66_90) );
AOI211_X1 g_57_96 (.ZN (n_57_96), .A (n_53_98), .B (n_54_96), .C1 (n_58_94), .C2 (n_64_91) );
AOI211_X1 g_59_95 (.ZN (n_59_95), .A (n_55_97), .B (n_52_97), .C1 (n_56_95), .C2 (n_62_92) );
AOI211_X1 g_61_94 (.ZN (n_61_94), .A (n_57_96), .B (n_51_99), .C1 (n_54_96), .C2 (n_60_93) );
AOI211_X1 g_63_93 (.ZN (n_63_93), .A (n_59_95), .B (n_53_98), .C1 (n_52_97), .C2 (n_58_94) );
AOI211_X1 g_65_92 (.ZN (n_65_92), .A (n_61_94), .B (n_55_97), .C1 (n_51_99), .C2 (n_56_95) );
AOI211_X1 g_67_91 (.ZN (n_67_91), .A (n_63_93), .B (n_57_96), .C1 (n_53_98), .C2 (n_54_96) );
AOI211_X1 g_69_90 (.ZN (n_69_90), .A (n_65_92), .B (n_59_95), .C1 (n_55_97), .C2 (n_52_97) );
AOI211_X1 g_71_89 (.ZN (n_71_89), .A (n_67_91), .B (n_61_94), .C1 (n_57_96), .C2 (n_51_99) );
AOI211_X1 g_73_88 (.ZN (n_73_88), .A (n_69_90), .B (n_63_93), .C1 (n_59_95), .C2 (n_53_98) );
AOI211_X1 g_72_90 (.ZN (n_72_90), .A (n_71_89), .B (n_65_92), .C1 (n_61_94), .C2 (n_55_97) );
AOI211_X1 g_74_89 (.ZN (n_74_89), .A (n_73_88), .B (n_67_91), .C1 (n_63_93), .C2 (n_57_96) );
AOI211_X1 g_76_88 (.ZN (n_76_88), .A (n_72_90), .B (n_69_90), .C1 (n_65_92), .C2 (n_59_95) );
AOI211_X1 g_78_87 (.ZN (n_78_87), .A (n_74_89), .B (n_71_89), .C1 (n_67_91), .C2 (n_61_94) );
AOI211_X1 g_80_86 (.ZN (n_80_86), .A (n_76_88), .B (n_73_88), .C1 (n_69_90), .C2 (n_63_93) );
AOI211_X1 g_82_85 (.ZN (n_82_85), .A (n_78_87), .B (n_72_90), .C1 (n_71_89), .C2 (n_65_92) );
AOI211_X1 g_81_87 (.ZN (n_81_87), .A (n_80_86), .B (n_74_89), .C1 (n_73_88), .C2 (n_67_91) );
AOI211_X1 g_83_86 (.ZN (n_83_86), .A (n_82_85), .B (n_76_88), .C1 (n_72_90), .C2 (n_69_90) );
AOI211_X1 g_85_85 (.ZN (n_85_85), .A (n_81_87), .B (n_78_87), .C1 (n_74_89), .C2 (n_71_89) );
AOI211_X1 g_87_84 (.ZN (n_87_84), .A (n_83_86), .B (n_80_86), .C1 (n_76_88), .C2 (n_73_88) );
AOI211_X1 g_89_83 (.ZN (n_89_83), .A (n_85_85), .B (n_82_85), .C1 (n_78_87), .C2 (n_72_90) );
AOI211_X1 g_90_81 (.ZN (n_90_81), .A (n_87_84), .B (n_81_87), .C1 (n_80_86), .C2 (n_74_89) );
AOI211_X1 g_92_80 (.ZN (n_92_80), .A (n_89_83), .B (n_83_86), .C1 (n_82_85), .C2 (n_76_88) );
AOI211_X1 g_94_79 (.ZN (n_94_79), .A (n_90_81), .B (n_85_85), .C1 (n_81_87), .C2 (n_78_87) );
AOI211_X1 g_96_78 (.ZN (n_96_78), .A (n_92_80), .B (n_87_84), .C1 (n_83_86), .C2 (n_80_86) );
AOI211_X1 g_98_77 (.ZN (n_98_77), .A (n_94_79), .B (n_89_83), .C1 (n_85_85), .C2 (n_82_85) );
AOI211_X1 g_100_76 (.ZN (n_100_76), .A (n_96_78), .B (n_90_81), .C1 (n_87_84), .C2 (n_81_87) );
AOI211_X1 g_99_78 (.ZN (n_99_78), .A (n_98_77), .B (n_92_80), .C1 (n_89_83), .C2 (n_83_86) );
AOI211_X1 g_101_77 (.ZN (n_101_77), .A (n_100_76), .B (n_94_79), .C1 (n_90_81), .C2 (n_85_85) );
AOI211_X1 g_103_76 (.ZN (n_103_76), .A (n_99_78), .B (n_96_78), .C1 (n_92_80), .C2 (n_87_84) );
AOI211_X1 g_105_75 (.ZN (n_105_75), .A (n_101_77), .B (n_98_77), .C1 (n_94_79), .C2 (n_89_83) );
AOI211_X1 g_107_74 (.ZN (n_107_74), .A (n_103_76), .B (n_100_76), .C1 (n_96_78), .C2 (n_90_81) );
AOI211_X1 g_109_73 (.ZN (n_109_73), .A (n_105_75), .B (n_99_78), .C1 (n_98_77), .C2 (n_92_80) );
AOI211_X1 g_108_75 (.ZN (n_108_75), .A (n_107_74), .B (n_101_77), .C1 (n_100_76), .C2 (n_94_79) );
AOI211_X1 g_110_74 (.ZN (n_110_74), .A (n_109_73), .B (n_103_76), .C1 (n_99_78), .C2 (n_96_78) );
AOI211_X1 g_112_73 (.ZN (n_112_73), .A (n_108_75), .B (n_105_75), .C1 (n_101_77), .C2 (n_98_77) );
AOI211_X1 g_114_72 (.ZN (n_114_72), .A (n_110_74), .B (n_107_74), .C1 (n_103_76), .C2 (n_100_76) );
AOI211_X1 g_116_71 (.ZN (n_116_71), .A (n_112_73), .B (n_109_73), .C1 (n_105_75), .C2 (n_99_78) );
AOI211_X1 g_118_70 (.ZN (n_118_70), .A (n_114_72), .B (n_108_75), .C1 (n_107_74), .C2 (n_101_77) );
AOI211_X1 g_120_69 (.ZN (n_120_69), .A (n_116_71), .B (n_110_74), .C1 (n_109_73), .C2 (n_103_76) );
AOI211_X1 g_122_68 (.ZN (n_122_68), .A (n_118_70), .B (n_112_73), .C1 (n_108_75), .C2 (n_105_75) );
AOI211_X1 g_124_67 (.ZN (n_124_67), .A (n_120_69), .B (n_114_72), .C1 (n_110_74), .C2 (n_107_74) );
AOI211_X1 g_126_68 (.ZN (n_126_68), .A (n_122_68), .B (n_116_71), .C1 (n_112_73), .C2 (n_109_73) );
AOI211_X1 g_124_69 (.ZN (n_124_69), .A (n_124_67), .B (n_118_70), .C1 (n_114_72), .C2 (n_108_75) );
AOI211_X1 g_125_67 (.ZN (n_125_67), .A (n_126_68), .B (n_120_69), .C1 (n_116_71), .C2 (n_110_74) );
AOI211_X1 g_126_65 (.ZN (n_126_65), .A (n_124_69), .B (n_122_68), .C1 (n_118_70), .C2 (n_112_73) );
AOI211_X1 g_124_66 (.ZN (n_124_66), .A (n_125_67), .B (n_124_67), .C1 (n_120_69), .C2 (n_114_72) );
AOI211_X1 g_122_67 (.ZN (n_122_67), .A (n_126_65), .B (n_126_68), .C1 (n_122_68), .C2 (n_116_71) );
AOI211_X1 g_120_68 (.ZN (n_120_68), .A (n_124_66), .B (n_124_69), .C1 (n_124_67), .C2 (n_118_70) );
AOI211_X1 g_118_69 (.ZN (n_118_69), .A (n_122_67), .B (n_125_67), .C1 (n_126_68), .C2 (n_120_69) );
AOI211_X1 g_116_70 (.ZN (n_116_70), .A (n_120_68), .B (n_126_65), .C1 (n_124_69), .C2 (n_122_68) );
AOI211_X1 g_114_71 (.ZN (n_114_71), .A (n_118_69), .B (n_124_66), .C1 (n_125_67), .C2 (n_124_67) );
AOI211_X1 g_112_72 (.ZN (n_112_72), .A (n_116_70), .B (n_122_67), .C1 (n_126_65), .C2 (n_126_68) );
AOI211_X1 g_110_73 (.ZN (n_110_73), .A (n_114_71), .B (n_120_68), .C1 (n_124_66), .C2 (n_124_69) );
AOI211_X1 g_108_74 (.ZN (n_108_74), .A (n_112_72), .B (n_118_69), .C1 (n_122_67), .C2 (n_125_67) );
AOI211_X1 g_106_75 (.ZN (n_106_75), .A (n_110_73), .B (n_116_70), .C1 (n_120_68), .C2 (n_126_65) );
AOI211_X1 g_104_76 (.ZN (n_104_76), .A (n_108_74), .B (n_114_71), .C1 (n_118_69), .C2 (n_124_66) );
AOI211_X1 g_102_77 (.ZN (n_102_77), .A (n_106_75), .B (n_112_72), .C1 (n_116_70), .C2 (n_122_67) );
AOI211_X1 g_100_78 (.ZN (n_100_78), .A (n_104_76), .B (n_110_73), .C1 (n_114_71), .C2 (n_120_68) );
AOI211_X1 g_98_79 (.ZN (n_98_79), .A (n_102_77), .B (n_108_74), .C1 (n_112_72), .C2 (n_118_69) );
AOI211_X1 g_96_80 (.ZN (n_96_80), .A (n_100_78), .B (n_106_75), .C1 (n_110_73), .C2 (n_116_70) );
AOI211_X1 g_94_81 (.ZN (n_94_81), .A (n_98_79), .B (n_104_76), .C1 (n_108_74), .C2 (n_114_71) );
AOI211_X1 g_92_82 (.ZN (n_92_82), .A (n_96_80), .B (n_102_77), .C1 (n_106_75), .C2 (n_112_72) );
AOI211_X1 g_93_80 (.ZN (n_93_80), .A (n_94_81), .B (n_100_78), .C1 (n_104_76), .C2 (n_110_73) );
AOI211_X1 g_91_81 (.ZN (n_91_81), .A (n_92_82), .B (n_98_79), .C1 (n_102_77), .C2 (n_108_74) );
AOI211_X1 g_89_82 (.ZN (n_89_82), .A (n_93_80), .B (n_96_80), .C1 (n_100_78), .C2 (n_106_75) );
AOI211_X1 g_87_83 (.ZN (n_87_83), .A (n_91_81), .B (n_94_81), .C1 (n_98_79), .C2 (n_104_76) );
AOI211_X1 g_85_84 (.ZN (n_85_84), .A (n_89_82), .B (n_92_82), .C1 (n_96_80), .C2 (n_102_77) );
AOI211_X1 g_83_85 (.ZN (n_83_85), .A (n_87_83), .B (n_93_80), .C1 (n_94_81), .C2 (n_100_78) );
AOI211_X1 g_81_86 (.ZN (n_81_86), .A (n_85_84), .B (n_91_81), .C1 (n_92_82), .C2 (n_98_79) );
AOI211_X1 g_79_87 (.ZN (n_79_87), .A (n_83_85), .B (n_89_82), .C1 (n_93_80), .C2 (n_96_80) );
AOI211_X1 g_77_88 (.ZN (n_77_88), .A (n_81_86), .B (n_87_83), .C1 (n_91_81), .C2 (n_94_81) );
AOI211_X1 g_75_89 (.ZN (n_75_89), .A (n_79_87), .B (n_85_84), .C1 (n_89_82), .C2 (n_92_82) );
AOI211_X1 g_73_90 (.ZN (n_73_90), .A (n_77_88), .B (n_83_85), .C1 (n_87_83), .C2 (n_93_80) );
AOI211_X1 g_71_91 (.ZN (n_71_91), .A (n_75_89), .B (n_81_86), .C1 (n_85_84), .C2 (n_91_81) );
AOI211_X1 g_72_89 (.ZN (n_72_89), .A (n_73_90), .B (n_79_87), .C1 (n_83_85), .C2 (n_89_82) );
AOI211_X1 g_70_90 (.ZN (n_70_90), .A (n_71_91), .B (n_77_88), .C1 (n_81_86), .C2 (n_87_83) );
AOI211_X1 g_68_91 (.ZN (n_68_91), .A (n_72_89), .B (n_75_89), .C1 (n_79_87), .C2 (n_85_84) );
AOI211_X1 g_66_92 (.ZN (n_66_92), .A (n_70_90), .B (n_73_90), .C1 (n_77_88), .C2 (n_83_85) );
AOI211_X1 g_64_93 (.ZN (n_64_93), .A (n_68_91), .B (n_71_91), .C1 (n_75_89), .C2 (n_81_86) );
AOI211_X1 g_62_94 (.ZN (n_62_94), .A (n_66_92), .B (n_72_89), .C1 (n_73_90), .C2 (n_79_87) );
AOI211_X1 g_60_95 (.ZN (n_60_95), .A (n_64_93), .B (n_70_90), .C1 (n_71_91), .C2 (n_77_88) );
AOI211_X1 g_58_96 (.ZN (n_58_96), .A (n_62_94), .B (n_68_91), .C1 (n_72_89), .C2 (n_75_89) );
AOI211_X1 g_56_97 (.ZN (n_56_97), .A (n_60_95), .B (n_66_92), .C1 (n_70_90), .C2 (n_73_90) );
AOI211_X1 g_54_98 (.ZN (n_54_98), .A (n_58_96), .B (n_64_93), .C1 (n_68_91), .C2 (n_71_91) );
AOI211_X1 g_52_99 (.ZN (n_52_99), .A (n_56_97), .B (n_62_94), .C1 (n_66_92), .C2 (n_72_89) );
AOI211_X1 g_50_100 (.ZN (n_50_100), .A (n_54_98), .B (n_60_95), .C1 (n_64_93), .C2 (n_70_90) );
AOI211_X1 g_48_101 (.ZN (n_48_101), .A (n_52_99), .B (n_58_96), .C1 (n_62_94), .C2 (n_68_91) );
AOI211_X1 g_46_102 (.ZN (n_46_102), .A (n_50_100), .B (n_56_97), .C1 (n_60_95), .C2 (n_66_92) );
AOI211_X1 g_44_103 (.ZN (n_44_103), .A (n_48_101), .B (n_54_98), .C1 (n_58_96), .C2 (n_64_93) );
AOI211_X1 g_42_104 (.ZN (n_42_104), .A (n_46_102), .B (n_52_99), .C1 (n_56_97), .C2 (n_62_94) );
AOI211_X1 g_40_105 (.ZN (n_40_105), .A (n_44_103), .B (n_50_100), .C1 (n_54_98), .C2 (n_60_95) );
AOI211_X1 g_41_103 (.ZN (n_41_103), .A (n_42_104), .B (n_48_101), .C1 (n_52_99), .C2 (n_58_96) );
AOI211_X1 g_39_104 (.ZN (n_39_104), .A (n_40_105), .B (n_46_102), .C1 (n_50_100), .C2 (n_56_97) );
AOI211_X1 g_37_105 (.ZN (n_37_105), .A (n_41_103), .B (n_44_103), .C1 (n_48_101), .C2 (n_54_98) );
AOI211_X1 g_35_106 (.ZN (n_35_106), .A (n_39_104), .B (n_42_104), .C1 (n_46_102), .C2 (n_52_99) );
AOI211_X1 g_33_107 (.ZN (n_33_107), .A (n_37_105), .B (n_40_105), .C1 (n_44_103), .C2 (n_50_100) );
AOI211_X1 g_31_108 (.ZN (n_31_108), .A (n_35_106), .B (n_41_103), .C1 (n_42_104), .C2 (n_48_101) );
AOI211_X1 g_29_109 (.ZN (n_29_109), .A (n_33_107), .B (n_39_104), .C1 (n_40_105), .C2 (n_46_102) );
AOI211_X1 g_27_110 (.ZN (n_27_110), .A (n_31_108), .B (n_37_105), .C1 (n_41_103), .C2 (n_44_103) );
AOI211_X1 g_25_111 (.ZN (n_25_111), .A (n_29_109), .B (n_35_106), .C1 (n_39_104), .C2 (n_42_104) );
AOI211_X1 g_23_112 (.ZN (n_23_112), .A (n_27_110), .B (n_33_107), .C1 (n_37_105), .C2 (n_40_105) );
AOI211_X1 g_21_111 (.ZN (n_21_111), .A (n_25_111), .B (n_31_108), .C1 (n_35_106), .C2 (n_41_103) );
AOI211_X1 g_19_110 (.ZN (n_19_110), .A (n_23_112), .B (n_29_109), .C1 (n_33_107), .C2 (n_39_104) );
AOI211_X1 g_17_111 (.ZN (n_17_111), .A (n_21_111), .B (n_27_110), .C1 (n_31_108), .C2 (n_37_105) );
AOI211_X1 g_15_112 (.ZN (n_15_112), .A (n_19_110), .B (n_25_111), .C1 (n_29_109), .C2 (n_35_106) );
AOI211_X1 g_13_113 (.ZN (n_13_113), .A (n_17_111), .B (n_23_112), .C1 (n_27_110), .C2 (n_33_107) );
AOI211_X1 g_11_114 (.ZN (n_11_114), .A (n_15_112), .B (n_21_111), .C1 (n_25_111), .C2 (n_31_108) );
AOI211_X1 g_13_115 (.ZN (n_13_115), .A (n_13_113), .B (n_19_110), .C1 (n_23_112), .C2 (n_29_109) );
AOI211_X1 g_11_116 (.ZN (n_11_116), .A (n_11_114), .B (n_17_111), .C1 (n_21_111), .C2 (n_27_110) );
AOI211_X1 g_10_118 (.ZN (n_10_118), .A (n_13_115), .B (n_15_112), .C1 (n_19_110), .C2 (n_25_111) );
AOI211_X1 g_8_119 (.ZN (n_8_119), .A (n_11_116), .B (n_13_113), .C1 (n_17_111), .C2 (n_23_112) );
AOI211_X1 g_7_121 (.ZN (n_7_121), .A (n_10_118), .B (n_11_114), .C1 (n_15_112), .C2 (n_21_111) );
AOI211_X1 g_6_119 (.ZN (n_6_119), .A (n_8_119), .B (n_13_115), .C1 (n_13_113), .C2 (n_19_110) );
AOI211_X1 g_5_121 (.ZN (n_5_121), .A (n_7_121), .B (n_11_116), .C1 (n_11_114), .C2 (n_17_111) );
AOI211_X1 g_4_123 (.ZN (n_4_123), .A (n_6_119), .B (n_10_118), .C1 (n_13_115), .C2 (n_15_112) );
AOI211_X1 g_3_125 (.ZN (n_3_125), .A (n_5_121), .B (n_8_119), .C1 (n_11_116), .C2 (n_13_113) );
AOI211_X1 g_5_126 (.ZN (n_5_126), .A (n_4_123), .B (n_7_121), .C1 (n_10_118), .C2 (n_11_114) );
AOI211_X1 g_3_127 (.ZN (n_3_127), .A (n_3_125), .B (n_6_119), .C1 (n_8_119), .C2 (n_13_115) );
AOI211_X1 g_1_128 (.ZN (n_1_128), .A (n_5_126), .B (n_5_121), .C1 (n_7_121), .C2 (n_11_116) );
AOI211_X1 g_2_126 (.ZN (n_2_126), .A (n_3_127), .B (n_4_123), .C1 (n_6_119), .C2 (n_10_118) );
AOI211_X1 g_4_125 (.ZN (n_4_125), .A (n_1_128), .B (n_3_125), .C1 (n_5_121), .C2 (n_8_119) );
AOI211_X1 g_6_124 (.ZN (n_6_124), .A (n_2_126), .B (n_5_126), .C1 (n_4_123), .C2 (n_7_121) );
AOI211_X1 g_7_122 (.ZN (n_7_122), .A (n_4_125), .B (n_3_127), .C1 (n_3_125), .C2 (n_6_119) );
AOI211_X1 g_5_123 (.ZN (n_5_123), .A (n_6_124), .B (n_1_128), .C1 (n_5_126), .C2 (n_5_121) );
AOI211_X1 g_3_124 (.ZN (n_3_124), .A (n_7_122), .B (n_2_126), .C1 (n_3_127), .C2 (n_4_123) );
AOI211_X1 g_4_122 (.ZN (n_4_122), .A (n_5_123), .B (n_4_125), .C1 (n_1_128), .C2 (n_3_125) );
AOI211_X1 g_6_121 (.ZN (n_6_121), .A (n_3_124), .B (n_6_124), .C1 (n_2_126), .C2 (n_5_126) );
AOI211_X1 g_8_120 (.ZN (n_8_120), .A (n_4_122), .B (n_7_122), .C1 (n_4_125), .C2 (n_3_127) );
AOI211_X1 g_10_119 (.ZN (n_10_119), .A (n_6_121), .B (n_5_123), .C1 (n_6_124), .C2 (n_1_128) );
AOI211_X1 g_8_118 (.ZN (n_8_118), .A (n_8_120), .B (n_3_124), .C1 (n_7_122), .C2 (n_2_126) );
AOI211_X1 g_9_116 (.ZN (n_9_116), .A (n_10_119), .B (n_4_122), .C1 (n_5_123), .C2 (n_4_125) );
AOI211_X1 g_7_115 (.ZN (n_7_115), .A (n_8_118), .B (n_6_121), .C1 (n_3_124), .C2 (n_6_124) );
AOI211_X1 g_6_117 (.ZN (n_6_117), .A (n_9_116), .B (n_8_120), .C1 (n_4_122), .C2 (n_7_122) );
AOI211_X1 g_8_116 (.ZN (n_8_116), .A (n_7_115), .B (n_10_119), .C1 (n_6_121), .C2 (n_5_123) );
AOI211_X1 g_9_114 (.ZN (n_9_114), .A (n_6_117), .B (n_8_118), .C1 (n_8_120), .C2 (n_3_124) );
AOI211_X1 g_11_115 (.ZN (n_11_115), .A (n_8_116), .B (n_9_116), .C1 (n_10_119), .C2 (n_4_122) );
AOI211_X1 g_13_114 (.ZN (n_13_114), .A (n_9_114), .B (n_7_115), .C1 (n_8_118), .C2 (n_6_121) );
AOI211_X1 g_15_113 (.ZN (n_15_113), .A (n_11_115), .B (n_6_117), .C1 (n_9_116), .C2 (n_8_120) );
AOI211_X1 g_17_112 (.ZN (n_17_112), .A (n_13_114), .B (n_8_116), .C1 (n_7_115), .C2 (n_10_119) );
AOI211_X1 g_19_111 (.ZN (n_19_111), .A (n_15_113), .B (n_9_114), .C1 (n_6_117), .C2 (n_8_118) );
AOI211_X1 g_21_110 (.ZN (n_21_110), .A (n_17_112), .B (n_11_115), .C1 (n_8_116), .C2 (n_9_116) );
AOI211_X1 g_23_111 (.ZN (n_23_111), .A (n_19_111), .B (n_13_114), .C1 (n_9_114), .C2 (n_7_115) );
AOI211_X1 g_21_112 (.ZN (n_21_112), .A (n_21_110), .B (n_15_113), .C1 (n_11_115), .C2 (n_6_117) );
AOI211_X1 g_19_113 (.ZN (n_19_113), .A (n_23_111), .B (n_17_112), .C1 (n_13_114), .C2 (n_8_116) );
AOI211_X1 g_20_111 (.ZN (n_20_111), .A (n_21_112), .B (n_19_111), .C1 (n_15_113), .C2 (n_9_114) );
AOI211_X1 g_18_112 (.ZN (n_18_112), .A (n_19_113), .B (n_21_110), .C1 (n_17_112), .C2 (n_11_115) );
AOI211_X1 g_16_113 (.ZN (n_16_113), .A (n_20_111), .B (n_23_111), .C1 (n_19_111), .C2 (n_13_114) );
AOI211_X1 g_14_114 (.ZN (n_14_114), .A (n_18_112), .B (n_21_112), .C1 (n_21_110), .C2 (n_15_113) );
AOI211_X1 g_12_115 (.ZN (n_12_115), .A (n_16_113), .B (n_19_113), .C1 (n_23_111), .C2 (n_17_112) );
AOI211_X1 g_10_116 (.ZN (n_10_116), .A (n_14_114), .B (n_20_111), .C1 (n_21_112), .C2 (n_19_111) );
AOI211_X1 g_8_117 (.ZN (n_8_117), .A (n_12_115), .B (n_18_112), .C1 (n_19_113), .C2 (n_21_110) );
AOI211_X1 g_7_119 (.ZN (n_7_119), .A (n_10_116), .B (n_16_113), .C1 (n_20_111), .C2 (n_23_111) );
AOI211_X1 g_9_118 (.ZN (n_9_118), .A (n_8_117), .B (n_14_114), .C1 (n_18_112), .C2 (n_21_112) );
AOI211_X1 g_11_117 (.ZN (n_11_117), .A (n_7_119), .B (n_12_115), .C1 (n_16_113), .C2 (n_19_113) );
AOI211_X1 g_13_116 (.ZN (n_13_116), .A (n_9_118), .B (n_10_116), .C1 (n_14_114), .C2 (n_20_111) );
AOI211_X1 g_15_115 (.ZN (n_15_115), .A (n_11_117), .B (n_8_117), .C1 (n_12_115), .C2 (n_18_112) );
AOI211_X1 g_17_114 (.ZN (n_17_114), .A (n_13_116), .B (n_7_119), .C1 (n_10_116), .C2 (n_16_113) );
AOI211_X1 g_16_116 (.ZN (n_16_116), .A (n_15_115), .B (n_9_118), .C1 (n_8_117), .C2 (n_14_114) );
AOI211_X1 g_15_114 (.ZN (n_15_114), .A (n_17_114), .B (n_11_117), .C1 (n_7_119), .C2 (n_12_115) );
AOI211_X1 g_17_113 (.ZN (n_17_113), .A (n_16_116), .B (n_13_116), .C1 (n_9_118), .C2 (n_10_116) );
AOI211_X1 g_19_112 (.ZN (n_19_112), .A (n_15_114), .B (n_15_115), .C1 (n_11_117), .C2 (n_8_117) );
AOI211_X1 g_18_114 (.ZN (n_18_114), .A (n_17_113), .B (n_17_114), .C1 (n_13_116), .C2 (n_7_119) );
AOI211_X1 g_20_113 (.ZN (n_20_113), .A (n_19_112), .B (n_16_116), .C1 (n_15_115), .C2 (n_9_118) );
AOI211_X1 g_22_112 (.ZN (n_22_112), .A (n_18_114), .B (n_15_114), .C1 (n_17_114), .C2 (n_11_117) );
AOI211_X1 g_24_113 (.ZN (n_24_113), .A (n_20_113), .B (n_17_113), .C1 (n_16_116), .C2 (n_13_116) );
AOI211_X1 g_26_112 (.ZN (n_26_112), .A (n_22_112), .B (n_19_112), .C1 (n_15_114), .C2 (n_15_115) );
AOI211_X1 g_28_111 (.ZN (n_28_111), .A (n_24_113), .B (n_18_114), .C1 (n_17_113), .C2 (n_17_114) );
AOI211_X1 g_26_110 (.ZN (n_26_110), .A (n_26_112), .B (n_20_113), .C1 (n_19_112), .C2 (n_16_116) );
AOI211_X1 g_28_109 (.ZN (n_28_109), .A (n_28_111), .B (n_22_112), .C1 (n_18_114), .C2 (n_15_114) );
AOI211_X1 g_30_108 (.ZN (n_30_108), .A (n_26_110), .B (n_24_113), .C1 (n_20_113), .C2 (n_17_113) );
AOI211_X1 g_29_110 (.ZN (n_29_110), .A (n_28_109), .B (n_26_112), .C1 (n_22_112), .C2 (n_19_112) );
AOI211_X1 g_31_109 (.ZN (n_31_109), .A (n_30_108), .B (n_28_111), .C1 (n_24_113), .C2 (n_18_114) );
AOI211_X1 g_30_111 (.ZN (n_30_111), .A (n_29_110), .B (n_26_110), .C1 (n_26_112), .C2 (n_20_113) );
AOI211_X1 g_28_110 (.ZN (n_28_110), .A (n_31_109), .B (n_28_109), .C1 (n_28_111), .C2 (n_22_112) );
AOI211_X1 g_26_111 (.ZN (n_26_111), .A (n_30_111), .B (n_30_108), .C1 (n_26_110), .C2 (n_24_113) );
AOI211_X1 g_28_112 (.ZN (n_28_112), .A (n_28_110), .B (n_29_110), .C1 (n_28_109), .C2 (n_26_112) );
AOI211_X1 g_26_113 (.ZN (n_26_113), .A (n_26_111), .B (n_31_109), .C1 (n_30_108), .C2 (n_28_111) );
AOI211_X1 g_27_111 (.ZN (n_27_111), .A (n_28_112), .B (n_30_111), .C1 (n_29_110), .C2 (n_26_110) );
AOI211_X1 g_25_112 (.ZN (n_25_112), .A (n_26_113), .B (n_28_110), .C1 (n_31_109), .C2 (n_28_109) );
AOI211_X1 g_23_113 (.ZN (n_23_113), .A (n_27_111), .B (n_26_111), .C1 (n_30_111), .C2 (n_30_108) );
AOI211_X1 g_22_111 (.ZN (n_22_111), .A (n_25_112), .B (n_28_112), .C1 (n_28_110), .C2 (n_29_110) );
AOI211_X1 g_24_112 (.ZN (n_24_112), .A (n_23_113), .B (n_26_113), .C1 (n_26_111), .C2 (n_31_109) );
AOI211_X1 g_22_113 (.ZN (n_22_113), .A (n_22_111), .B (n_27_111), .C1 (n_28_112), .C2 (n_30_111) );
AOI211_X1 g_20_112 (.ZN (n_20_112), .A (n_24_112), .B (n_25_112), .C1 (n_26_113), .C2 (n_28_110) );
AOI211_X1 g_18_113 (.ZN (n_18_113), .A (n_22_113), .B (n_23_113), .C1 (n_27_111), .C2 (n_26_111) );
AOI211_X1 g_16_114 (.ZN (n_16_114), .A (n_20_112), .B (n_22_111), .C1 (n_25_112), .C2 (n_28_112) );
AOI211_X1 g_14_115 (.ZN (n_14_115), .A (n_18_113), .B (n_24_112), .C1 (n_23_113), .C2 (n_26_113) );
AOI211_X1 g_12_116 (.ZN (n_12_116), .A (n_16_114), .B (n_22_113), .C1 (n_22_111), .C2 (n_27_111) );
AOI211_X1 g_10_117 (.ZN (n_10_117), .A (n_14_115), .B (n_20_112), .C1 (n_24_112), .C2 (n_25_112) );
AOI211_X1 g_12_118 (.ZN (n_12_118), .A (n_12_116), .B (n_18_113), .C1 (n_22_113), .C2 (n_23_113) );
AOI211_X1 g_14_117 (.ZN (n_14_117), .A (n_10_117), .B (n_16_114), .C1 (n_20_112), .C2 (n_22_111) );
AOI211_X1 g_13_119 (.ZN (n_13_119), .A (n_12_118), .B (n_14_115), .C1 (n_18_113), .C2 (n_24_112) );
AOI211_X1 g_12_117 (.ZN (n_12_117), .A (n_14_117), .B (n_12_116), .C1 (n_16_114), .C2 (n_22_113) );
AOI211_X1 g_14_116 (.ZN (n_14_116), .A (n_13_119), .B (n_10_117), .C1 (n_14_115), .C2 (n_20_112) );
AOI211_X1 g_16_115 (.ZN (n_16_115), .A (n_12_117), .B (n_12_118), .C1 (n_12_116), .C2 (n_18_113) );
AOI211_X1 g_15_117 (.ZN (n_15_117), .A (n_14_116), .B (n_14_117), .C1 (n_10_117), .C2 (n_16_114) );
AOI211_X1 g_17_116 (.ZN (n_17_116), .A (n_16_115), .B (n_13_119), .C1 (n_12_118), .C2 (n_14_115) );
AOI211_X1 g_19_115 (.ZN (n_19_115), .A (n_15_117), .B (n_12_117), .C1 (n_14_117), .C2 (n_12_116) );
AOI211_X1 g_21_114 (.ZN (n_21_114), .A (n_17_116), .B (n_14_116), .C1 (n_13_119), .C2 (n_10_117) );
AOI211_X1 g_23_115 (.ZN (n_23_115), .A (n_19_115), .B (n_16_115), .C1 (n_12_117), .C2 (n_12_118) );
AOI211_X1 g_25_114 (.ZN (n_25_114), .A (n_21_114), .B (n_15_117), .C1 (n_14_116), .C2 (n_14_117) );
AOI211_X1 g_27_113 (.ZN (n_27_113), .A (n_23_115), .B (n_17_116), .C1 (n_16_115), .C2 (n_13_119) );
AOI211_X1 g_29_112 (.ZN (n_29_112), .A (n_25_114), .B (n_19_115), .C1 (n_15_117), .C2 (n_12_117) );
AOI211_X1 g_30_110 (.ZN (n_30_110), .A (n_27_113), .B (n_21_114), .C1 (n_17_116), .C2 (n_14_116) );
AOI211_X1 g_32_109 (.ZN (n_32_109), .A (n_29_112), .B (n_23_115), .C1 (n_19_115), .C2 (n_16_115) );
AOI211_X1 g_34_108 (.ZN (n_34_108), .A (n_30_110), .B (n_25_114), .C1 (n_21_114), .C2 (n_15_117) );
AOI211_X1 g_36_107 (.ZN (n_36_107), .A (n_32_109), .B (n_27_113), .C1 (n_23_115), .C2 (n_17_116) );
AOI211_X1 g_38_106 (.ZN (n_38_106), .A (n_34_108), .B (n_29_112), .C1 (n_25_114), .C2 (n_19_115) );
AOI211_X1 g_37_108 (.ZN (n_37_108), .A (n_36_107), .B (n_30_110), .C1 (n_27_113), .C2 (n_21_114) );
AOI211_X1 g_39_107 (.ZN (n_39_107), .A (n_38_106), .B (n_32_109), .C1 (n_29_112), .C2 (n_23_115) );
AOI211_X1 g_41_106 (.ZN (n_41_106), .A (n_37_108), .B (n_34_108), .C1 (n_30_110), .C2 (n_25_114) );
AOI211_X1 g_39_105 (.ZN (n_39_105), .A (n_39_107), .B (n_36_107), .C1 (n_32_109), .C2 (n_27_113) );
AOI211_X1 g_41_104 (.ZN (n_41_104), .A (n_41_106), .B (n_38_106), .C1 (n_34_108), .C2 (n_29_112) );
AOI211_X1 g_43_103 (.ZN (n_43_103), .A (n_39_105), .B (n_37_108), .C1 (n_36_107), .C2 (n_30_110) );
AOI211_X1 g_45_102 (.ZN (n_45_102), .A (n_41_104), .B (n_39_107), .C1 (n_38_106), .C2 (n_32_109) );
AOI211_X1 g_47_101 (.ZN (n_47_101), .A (n_43_103), .B (n_41_106), .C1 (n_37_108), .C2 (n_34_108) );
AOI211_X1 g_49_100 (.ZN (n_49_100), .A (n_45_102), .B (n_39_105), .C1 (n_39_107), .C2 (n_36_107) );
AOI211_X1 g_48_102 (.ZN (n_48_102), .A (n_47_101), .B (n_41_104), .C1 (n_41_106), .C2 (n_38_106) );
AOI211_X1 g_50_101 (.ZN (n_50_101), .A (n_49_100), .B (n_43_103), .C1 (n_39_105), .C2 (n_37_108) );
AOI211_X1 g_52_100 (.ZN (n_52_100), .A (n_48_102), .B (n_45_102), .C1 (n_41_104), .C2 (n_39_107) );
AOI211_X1 g_54_99 (.ZN (n_54_99), .A (n_50_101), .B (n_47_101), .C1 (n_43_103), .C2 (n_41_106) );
AOI211_X1 g_56_98 (.ZN (n_56_98), .A (n_52_100), .B (n_49_100), .C1 (n_45_102), .C2 (n_39_105) );
AOI211_X1 g_58_97 (.ZN (n_58_97), .A (n_54_99), .B (n_48_102), .C1 (n_47_101), .C2 (n_41_104) );
AOI211_X1 g_60_96 (.ZN (n_60_96), .A (n_56_98), .B (n_50_101), .C1 (n_49_100), .C2 (n_43_103) );
AOI211_X1 g_62_95 (.ZN (n_62_95), .A (n_58_97), .B (n_52_100), .C1 (n_48_102), .C2 (n_45_102) );
AOI211_X1 g_64_94 (.ZN (n_64_94), .A (n_60_96), .B (n_54_99), .C1 (n_50_101), .C2 (n_47_101) );
AOI211_X1 g_66_93 (.ZN (n_66_93), .A (n_62_95), .B (n_56_98), .C1 (n_52_100), .C2 (n_49_100) );
AOI211_X1 g_68_92 (.ZN (n_68_92), .A (n_64_94), .B (n_58_97), .C1 (n_54_99), .C2 (n_48_102) );
AOI211_X1 g_70_91 (.ZN (n_70_91), .A (n_66_93), .B (n_60_96), .C1 (n_56_98), .C2 (n_50_101) );
AOI211_X1 g_69_93 (.ZN (n_69_93), .A (n_68_92), .B (n_62_95), .C1 (n_58_97), .C2 (n_52_100) );
AOI211_X1 g_67_92 (.ZN (n_67_92), .A (n_70_91), .B (n_64_94), .C1 (n_60_96), .C2 (n_54_99) );
AOI211_X1 g_69_91 (.ZN (n_69_91), .A (n_69_93), .B (n_66_93), .C1 (n_62_95), .C2 (n_56_98) );
AOI211_X1 g_71_90 (.ZN (n_71_90), .A (n_67_92), .B (n_68_92), .C1 (n_64_94), .C2 (n_58_97) );
AOI211_X1 g_73_89 (.ZN (n_73_89), .A (n_69_91), .B (n_70_91), .C1 (n_66_93), .C2 (n_60_96) );
AOI211_X1 g_72_91 (.ZN (n_72_91), .A (n_71_90), .B (n_69_93), .C1 (n_68_92), .C2 (n_62_95) );
AOI211_X1 g_74_90 (.ZN (n_74_90), .A (n_73_89), .B (n_67_92), .C1 (n_70_91), .C2 (n_64_94) );
AOI211_X1 g_73_92 (.ZN (n_73_92), .A (n_72_91), .B (n_69_91), .C1 (n_69_93), .C2 (n_66_93) );
AOI211_X1 g_75_91 (.ZN (n_75_91), .A (n_74_90), .B (n_71_90), .C1 (n_67_92), .C2 (n_68_92) );
AOI211_X1 g_77_90 (.ZN (n_77_90), .A (n_73_92), .B (n_73_89), .C1 (n_69_91), .C2 (n_70_91) );
AOI211_X1 g_78_88 (.ZN (n_78_88), .A (n_75_91), .B (n_72_91), .C1 (n_71_90), .C2 (n_69_93) );
AOI211_X1 g_80_87 (.ZN (n_80_87), .A (n_77_90), .B (n_74_90), .C1 (n_73_89), .C2 (n_67_92) );
AOI211_X1 g_82_86 (.ZN (n_82_86), .A (n_78_88), .B (n_73_92), .C1 (n_72_91), .C2 (n_69_91) );
AOI211_X1 g_84_85 (.ZN (n_84_85), .A (n_80_87), .B (n_75_91), .C1 (n_74_90), .C2 (n_71_90) );
AOI211_X1 g_86_84 (.ZN (n_86_84), .A (n_82_86), .B (n_77_90), .C1 (n_73_92), .C2 (n_73_89) );
AOI211_X1 g_85_86 (.ZN (n_85_86), .A (n_84_85), .B (n_78_88), .C1 (n_75_91), .C2 (n_72_91) );
AOI211_X1 g_87_85 (.ZN (n_87_85), .A (n_86_84), .B (n_80_87), .C1 (n_77_90), .C2 (n_74_90) );
AOI211_X1 g_89_84 (.ZN (n_89_84), .A (n_85_86), .B (n_82_86), .C1 (n_78_88), .C2 (n_73_92) );
AOI211_X1 g_91_83 (.ZN (n_91_83), .A (n_87_85), .B (n_84_85), .C1 (n_80_87), .C2 (n_75_91) );
AOI211_X1 g_93_82 (.ZN (n_93_82), .A (n_89_84), .B (n_86_84), .C1 (n_82_86), .C2 (n_77_90) );
AOI211_X1 g_95_81 (.ZN (n_95_81), .A (n_91_83), .B (n_85_86), .C1 (n_84_85), .C2 (n_78_88) );
AOI211_X1 g_97_80 (.ZN (n_97_80), .A (n_93_82), .B (n_87_85), .C1 (n_86_84), .C2 (n_80_87) );
AOI211_X1 g_99_79 (.ZN (n_99_79), .A (n_95_81), .B (n_89_84), .C1 (n_85_86), .C2 (n_82_86) );
AOI211_X1 g_101_78 (.ZN (n_101_78), .A (n_97_80), .B (n_91_83), .C1 (n_87_85), .C2 (n_84_85) );
AOI211_X1 g_103_77 (.ZN (n_103_77), .A (n_99_79), .B (n_93_82), .C1 (n_89_84), .C2 (n_86_84) );
AOI211_X1 g_105_76 (.ZN (n_105_76), .A (n_101_78), .B (n_95_81), .C1 (n_91_83), .C2 (n_85_86) );
AOI211_X1 g_107_75 (.ZN (n_107_75), .A (n_103_77), .B (n_97_80), .C1 (n_93_82), .C2 (n_87_85) );
AOI211_X1 g_109_74 (.ZN (n_109_74), .A (n_105_76), .B (n_99_79), .C1 (n_95_81), .C2 (n_89_84) );
AOI211_X1 g_111_73 (.ZN (n_111_73), .A (n_107_75), .B (n_101_78), .C1 (n_97_80), .C2 (n_91_83) );
AOI211_X1 g_113_72 (.ZN (n_113_72), .A (n_109_74), .B (n_103_77), .C1 (n_99_79), .C2 (n_93_82) );
AOI211_X1 g_115_71 (.ZN (n_115_71), .A (n_111_73), .B (n_105_76), .C1 (n_101_78), .C2 (n_95_81) );
AOI211_X1 g_117_70 (.ZN (n_117_70), .A (n_113_72), .B (n_107_75), .C1 (n_103_77), .C2 (n_97_80) );
AOI211_X1 g_119_69 (.ZN (n_119_69), .A (n_115_71), .B (n_109_74), .C1 (n_105_76), .C2 (n_99_79) );
AOI211_X1 g_118_71 (.ZN (n_118_71), .A (n_117_70), .B (n_111_73), .C1 (n_107_75), .C2 (n_101_78) );
AOI211_X1 g_120_70 (.ZN (n_120_70), .A (n_119_69), .B (n_113_72), .C1 (n_109_74), .C2 (n_103_77) );
AOI211_X1 g_122_69 (.ZN (n_122_69), .A (n_118_71), .B (n_115_71), .C1 (n_111_73), .C2 (n_105_76) );
AOI211_X1 g_124_68 (.ZN (n_124_68), .A (n_120_70), .B (n_117_70), .C1 (n_113_72), .C2 (n_107_75) );
AOI211_X1 g_126_67 (.ZN (n_126_67), .A (n_122_69), .B (n_119_69), .C1 (n_115_71), .C2 (n_109_74) );
AOI211_X1 g_128_66 (.ZN (n_128_66), .A (n_124_68), .B (n_118_71), .C1 (n_117_70), .C2 (n_111_73) );
AOI211_X1 g_127_68 (.ZN (n_127_68), .A (n_126_67), .B (n_120_70), .C1 (n_119_69), .C2 (n_113_72) );
AOI211_X1 g_125_69 (.ZN (n_125_69), .A (n_128_66), .B (n_122_69), .C1 (n_118_71), .C2 (n_115_71) );
AOI211_X1 g_123_68 (.ZN (n_123_68), .A (n_127_68), .B (n_124_68), .C1 (n_120_70), .C2 (n_117_70) );
AOI211_X1 g_121_69 (.ZN (n_121_69), .A (n_125_69), .B (n_126_67), .C1 (n_122_69), .C2 (n_119_69) );
AOI211_X1 g_119_70 (.ZN (n_119_70), .A (n_123_68), .B (n_128_66), .C1 (n_124_68), .C2 (n_118_71) );
AOI211_X1 g_117_71 (.ZN (n_117_71), .A (n_121_69), .B (n_127_68), .C1 (n_126_67), .C2 (n_120_70) );
AOI211_X1 g_115_72 (.ZN (n_115_72), .A (n_119_70), .B (n_125_69), .C1 (n_128_66), .C2 (n_122_69) );
AOI211_X1 g_113_73 (.ZN (n_113_73), .A (n_117_71), .B (n_123_68), .C1 (n_127_68), .C2 (n_124_68) );
AOI211_X1 g_111_74 (.ZN (n_111_74), .A (n_115_72), .B (n_121_69), .C1 (n_125_69), .C2 (n_126_67) );
AOI211_X1 g_109_75 (.ZN (n_109_75), .A (n_113_73), .B (n_119_70), .C1 (n_123_68), .C2 (n_128_66) );
AOI211_X1 g_107_76 (.ZN (n_107_76), .A (n_111_74), .B (n_117_71), .C1 (n_121_69), .C2 (n_127_68) );
AOI211_X1 g_105_77 (.ZN (n_105_77), .A (n_109_75), .B (n_115_72), .C1 (n_119_70), .C2 (n_125_69) );
AOI211_X1 g_103_78 (.ZN (n_103_78), .A (n_107_76), .B (n_113_73), .C1 (n_117_71), .C2 (n_123_68) );
AOI211_X1 g_101_79 (.ZN (n_101_79), .A (n_105_77), .B (n_111_74), .C1 (n_115_72), .C2 (n_121_69) );
AOI211_X1 g_99_80 (.ZN (n_99_80), .A (n_103_78), .B (n_109_75), .C1 (n_113_73), .C2 (n_119_70) );
AOI211_X1 g_97_79 (.ZN (n_97_79), .A (n_101_79), .B (n_107_76), .C1 (n_111_74), .C2 (n_117_71) );
AOI211_X1 g_95_80 (.ZN (n_95_80), .A (n_99_80), .B (n_105_77), .C1 (n_109_75), .C2 (n_115_72) );
AOI211_X1 g_93_81 (.ZN (n_93_81), .A (n_97_79), .B (n_103_78), .C1 (n_107_76), .C2 (n_113_73) );
AOI211_X1 g_91_82 (.ZN (n_91_82), .A (n_95_80), .B (n_101_79), .C1 (n_105_77), .C2 (n_111_74) );
AOI211_X1 g_90_84 (.ZN (n_90_84), .A (n_93_81), .B (n_99_80), .C1 (n_103_78), .C2 (n_109_75) );
AOI211_X1 g_92_83 (.ZN (n_92_83), .A (n_91_82), .B (n_97_79), .C1 (n_101_79), .C2 (n_107_76) );
AOI211_X1 g_94_82 (.ZN (n_94_82), .A (n_90_84), .B (n_95_80), .C1 (n_99_80), .C2 (n_105_77) );
AOI211_X1 g_96_81 (.ZN (n_96_81), .A (n_92_83), .B (n_93_81), .C1 (n_97_79), .C2 (n_103_78) );
AOI211_X1 g_98_80 (.ZN (n_98_80), .A (n_94_82), .B (n_91_82), .C1 (n_95_80), .C2 (n_101_79) );
AOI211_X1 g_100_79 (.ZN (n_100_79), .A (n_96_81), .B (n_90_84), .C1 (n_93_81), .C2 (n_99_80) );
AOI211_X1 g_102_78 (.ZN (n_102_78), .A (n_98_80), .B (n_92_83), .C1 (n_91_82), .C2 (n_97_79) );
AOI211_X1 g_104_77 (.ZN (n_104_77), .A (n_100_79), .B (n_94_82), .C1 (n_90_84), .C2 (n_95_80) );
AOI211_X1 g_106_76 (.ZN (n_106_76), .A (n_102_78), .B (n_96_81), .C1 (n_92_83), .C2 (n_93_81) );
AOI211_X1 g_105_78 (.ZN (n_105_78), .A (n_104_77), .B (n_98_80), .C1 (n_94_82), .C2 (n_91_82) );
AOI211_X1 g_107_77 (.ZN (n_107_77), .A (n_106_76), .B (n_100_79), .C1 (n_96_81), .C2 (n_90_84) );
AOI211_X1 g_109_76 (.ZN (n_109_76), .A (n_105_78), .B (n_102_78), .C1 (n_98_80), .C2 (n_92_83) );
AOI211_X1 g_111_75 (.ZN (n_111_75), .A (n_107_77), .B (n_104_77), .C1 (n_100_79), .C2 (n_94_82) );
AOI211_X1 g_113_74 (.ZN (n_113_74), .A (n_109_76), .B (n_106_76), .C1 (n_102_78), .C2 (n_96_81) );
AOI211_X1 g_115_73 (.ZN (n_115_73), .A (n_111_75), .B (n_105_78), .C1 (n_104_77), .C2 (n_98_80) );
AOI211_X1 g_117_72 (.ZN (n_117_72), .A (n_113_74), .B (n_107_77), .C1 (n_106_76), .C2 (n_100_79) );
AOI211_X1 g_119_71 (.ZN (n_119_71), .A (n_115_73), .B (n_109_76), .C1 (n_105_78), .C2 (n_102_78) );
AOI211_X1 g_121_70 (.ZN (n_121_70), .A (n_117_72), .B (n_111_75), .C1 (n_107_77), .C2 (n_104_77) );
AOI211_X1 g_123_69 (.ZN (n_123_69), .A (n_119_71), .B (n_113_74), .C1 (n_109_76), .C2 (n_106_76) );
AOI211_X1 g_125_68 (.ZN (n_125_68), .A (n_121_70), .B (n_115_73), .C1 (n_111_75), .C2 (n_105_78) );
AOI211_X1 g_127_67 (.ZN (n_127_67), .A (n_123_69), .B (n_117_72), .C1 (n_113_74), .C2 (n_107_77) );
AOI211_X1 g_129_66 (.ZN (n_129_66), .A (n_125_68), .B (n_119_71), .C1 (n_115_73), .C2 (n_109_76) );
AOI211_X1 g_131_65 (.ZN (n_131_65), .A (n_127_67), .B (n_121_70), .C1 (n_117_72), .C2 (n_111_75) );
AOI211_X1 g_130_67 (.ZN (n_130_67), .A (n_129_66), .B (n_123_69), .C1 (n_119_71), .C2 (n_113_74) );
AOI211_X1 g_128_68 (.ZN (n_128_68), .A (n_131_65), .B (n_125_68), .C1 (n_121_70), .C2 (n_115_73) );
AOI211_X1 g_126_69 (.ZN (n_126_69), .A (n_130_67), .B (n_127_67), .C1 (n_123_69), .C2 (n_117_72) );
AOI211_X1 g_124_70 (.ZN (n_124_70), .A (n_128_68), .B (n_129_66), .C1 (n_125_68), .C2 (n_119_71) );
AOI211_X1 g_122_71 (.ZN (n_122_71), .A (n_126_69), .B (n_131_65), .C1 (n_127_67), .C2 (n_121_70) );
AOI211_X1 g_120_72 (.ZN (n_120_72), .A (n_124_70), .B (n_130_67), .C1 (n_129_66), .C2 (n_123_69) );
AOI211_X1 g_118_73 (.ZN (n_118_73), .A (n_122_71), .B (n_128_68), .C1 (n_131_65), .C2 (n_125_68) );
AOI211_X1 g_116_72 (.ZN (n_116_72), .A (n_120_72), .B (n_126_69), .C1 (n_130_67), .C2 (n_127_67) );
AOI211_X1 g_114_73 (.ZN (n_114_73), .A (n_118_73), .B (n_124_70), .C1 (n_128_68), .C2 (n_129_66) );
AOI211_X1 g_112_74 (.ZN (n_112_74), .A (n_116_72), .B (n_122_71), .C1 (n_126_69), .C2 (n_131_65) );
AOI211_X1 g_110_75 (.ZN (n_110_75), .A (n_114_73), .B (n_120_72), .C1 (n_124_70), .C2 (n_130_67) );
AOI211_X1 g_108_76 (.ZN (n_108_76), .A (n_112_74), .B (n_118_73), .C1 (n_122_71), .C2 (n_128_68) );
AOI211_X1 g_106_77 (.ZN (n_106_77), .A (n_110_75), .B (n_116_72), .C1 (n_120_72), .C2 (n_126_69) );
AOI211_X1 g_104_78 (.ZN (n_104_78), .A (n_108_76), .B (n_114_73), .C1 (n_118_73), .C2 (n_124_70) );
AOI211_X1 g_102_79 (.ZN (n_102_79), .A (n_106_77), .B (n_112_74), .C1 (n_116_72), .C2 (n_122_71) );
AOI211_X1 g_100_80 (.ZN (n_100_80), .A (n_104_78), .B (n_110_75), .C1 (n_114_73), .C2 (n_120_72) );
AOI211_X1 g_98_81 (.ZN (n_98_81), .A (n_102_79), .B (n_108_76), .C1 (n_112_74), .C2 (n_118_73) );
AOI211_X1 g_96_82 (.ZN (n_96_82), .A (n_100_80), .B (n_106_77), .C1 (n_110_75), .C2 (n_116_72) );
AOI211_X1 g_94_83 (.ZN (n_94_83), .A (n_98_81), .B (n_104_78), .C1 (n_108_76), .C2 (n_114_73) );
AOI211_X1 g_92_84 (.ZN (n_92_84), .A (n_96_82), .B (n_102_79), .C1 (n_106_77), .C2 (n_112_74) );
AOI211_X1 g_90_83 (.ZN (n_90_83), .A (n_94_83), .B (n_100_80), .C1 (n_104_78), .C2 (n_110_75) );
AOI211_X1 g_88_84 (.ZN (n_88_84), .A (n_92_84), .B (n_98_81), .C1 (n_102_79), .C2 (n_108_76) );
AOI211_X1 g_86_85 (.ZN (n_86_85), .A (n_90_83), .B (n_96_82), .C1 (n_100_80), .C2 (n_106_77) );
AOI211_X1 g_84_86 (.ZN (n_84_86), .A (n_88_84), .B (n_94_83), .C1 (n_98_81), .C2 (n_104_78) );
AOI211_X1 g_82_87 (.ZN (n_82_87), .A (n_86_85), .B (n_92_84), .C1 (n_96_82), .C2 (n_102_79) );
AOI211_X1 g_80_88 (.ZN (n_80_88), .A (n_84_86), .B (n_90_83), .C1 (n_94_83), .C2 (n_100_80) );
AOI211_X1 g_78_89 (.ZN (n_78_89), .A (n_82_87), .B (n_88_84), .C1 (n_92_84), .C2 (n_98_81) );
AOI211_X1 g_76_90 (.ZN (n_76_90), .A (n_80_88), .B (n_86_85), .C1 (n_90_83), .C2 (n_96_82) );
AOI211_X1 g_74_91 (.ZN (n_74_91), .A (n_78_89), .B (n_84_86), .C1 (n_88_84), .C2 (n_94_83) );
AOI211_X1 g_72_92 (.ZN (n_72_92), .A (n_76_90), .B (n_82_87), .C1 (n_86_85), .C2 (n_92_84) );
AOI211_X1 g_70_93 (.ZN (n_70_93), .A (n_74_91), .B (n_80_88), .C1 (n_84_86), .C2 (n_90_83) );
AOI211_X1 g_68_94 (.ZN (n_68_94), .A (n_72_92), .B (n_78_89), .C1 (n_82_87), .C2 (n_88_84) );
AOI211_X1 g_69_92 (.ZN (n_69_92), .A (n_70_93), .B (n_76_90), .C1 (n_80_88), .C2 (n_86_85) );
AOI211_X1 g_67_93 (.ZN (n_67_93), .A (n_68_94), .B (n_74_91), .C1 (n_78_89), .C2 (n_84_86) );
AOI211_X1 g_65_94 (.ZN (n_65_94), .A (n_69_92), .B (n_72_92), .C1 (n_76_90), .C2 (n_82_87) );
AOI211_X1 g_63_95 (.ZN (n_63_95), .A (n_67_93), .B (n_70_93), .C1 (n_74_91), .C2 (n_80_88) );
AOI211_X1 g_61_96 (.ZN (n_61_96), .A (n_65_94), .B (n_68_94), .C1 (n_72_92), .C2 (n_78_89) );
AOI211_X1 g_59_97 (.ZN (n_59_97), .A (n_63_95), .B (n_69_92), .C1 (n_70_93), .C2 (n_76_90) );
AOI211_X1 g_57_98 (.ZN (n_57_98), .A (n_61_96), .B (n_67_93), .C1 (n_68_94), .C2 (n_74_91) );
AOI211_X1 g_55_99 (.ZN (n_55_99), .A (n_59_97), .B (n_65_94), .C1 (n_69_92), .C2 (n_72_92) );
AOI211_X1 g_53_100 (.ZN (n_53_100), .A (n_57_98), .B (n_63_95), .C1 (n_67_93), .C2 (n_70_93) );
AOI211_X1 g_51_101 (.ZN (n_51_101), .A (n_55_99), .B (n_61_96), .C1 (n_65_94), .C2 (n_68_94) );
AOI211_X1 g_49_102 (.ZN (n_49_102), .A (n_53_100), .B (n_59_97), .C1 (n_63_95), .C2 (n_69_92) );
AOI211_X1 g_47_103 (.ZN (n_47_103), .A (n_51_101), .B (n_57_98), .C1 (n_61_96), .C2 (n_67_93) );
AOI211_X1 g_45_104 (.ZN (n_45_104), .A (n_49_102), .B (n_55_99), .C1 (n_59_97), .C2 (n_65_94) );
AOI211_X1 g_43_105 (.ZN (n_43_105), .A (n_47_103), .B (n_53_100), .C1 (n_57_98), .C2 (n_63_95) );
AOI211_X1 g_42_107 (.ZN (n_42_107), .A (n_45_104), .B (n_51_101), .C1 (n_55_99), .C2 (n_61_96) );
AOI211_X1 g_41_105 (.ZN (n_41_105), .A (n_43_105), .B (n_49_102), .C1 (n_53_100), .C2 (n_59_97) );
AOI211_X1 g_43_104 (.ZN (n_43_104), .A (n_42_107), .B (n_47_103), .C1 (n_51_101), .C2 (n_57_98) );
AOI211_X1 g_42_106 (.ZN (n_42_106), .A (n_41_105), .B (n_45_104), .C1 (n_49_102), .C2 (n_55_99) );
AOI211_X1 g_44_105 (.ZN (n_44_105), .A (n_43_104), .B (n_43_105), .C1 (n_47_103), .C2 (n_53_100) );
AOI211_X1 g_46_104 (.ZN (n_46_104), .A (n_42_106), .B (n_42_107), .C1 (n_45_104), .C2 (n_51_101) );
AOI211_X1 g_47_102 (.ZN (n_47_102), .A (n_44_105), .B (n_41_105), .C1 (n_43_105), .C2 (n_49_102) );
AOI211_X1 g_49_101 (.ZN (n_49_101), .A (n_46_104), .B (n_43_104), .C1 (n_42_107), .C2 (n_47_103) );
AOI211_X1 g_51_100 (.ZN (n_51_100), .A (n_47_102), .B (n_42_106), .C1 (n_41_105), .C2 (n_45_104) );
AOI211_X1 g_53_99 (.ZN (n_53_99), .A (n_49_101), .B (n_44_105), .C1 (n_43_104), .C2 (n_43_105) );
AOI211_X1 g_55_98 (.ZN (n_55_98), .A (n_51_100), .B (n_46_104), .C1 (n_42_106), .C2 (n_42_107) );
AOI211_X1 g_57_97 (.ZN (n_57_97), .A (n_53_99), .B (n_47_102), .C1 (n_44_105), .C2 (n_41_105) );
AOI211_X1 g_59_96 (.ZN (n_59_96), .A (n_55_98), .B (n_49_101), .C1 (n_46_104), .C2 (n_43_104) );
AOI211_X1 g_61_95 (.ZN (n_61_95), .A (n_57_97), .B (n_51_100), .C1 (n_47_102), .C2 (n_42_106) );
AOI211_X1 g_63_94 (.ZN (n_63_94), .A (n_59_96), .B (n_53_99), .C1 (n_49_101), .C2 (n_44_105) );
AOI211_X1 g_65_93 (.ZN (n_65_93), .A (n_61_95), .B (n_55_98), .C1 (n_51_100), .C2 (n_46_104) );
AOI211_X1 g_66_95 (.ZN (n_66_95), .A (n_63_94), .B (n_57_97), .C1 (n_53_99), .C2 (n_47_102) );
AOI211_X1 g_64_96 (.ZN (n_64_96), .A (n_65_93), .B (n_59_96), .C1 (n_55_98), .C2 (n_49_101) );
AOI211_X1 g_62_97 (.ZN (n_62_97), .A (n_66_95), .B (n_61_95), .C1 (n_57_97), .C2 (n_51_100) );
AOI211_X1 g_60_98 (.ZN (n_60_98), .A (n_64_96), .B (n_63_94), .C1 (n_59_96), .C2 (n_53_99) );
AOI211_X1 g_58_99 (.ZN (n_58_99), .A (n_62_97), .B (n_65_93), .C1 (n_61_95), .C2 (n_55_98) );
AOI211_X1 g_56_100 (.ZN (n_56_100), .A (n_60_98), .B (n_66_95), .C1 (n_63_94), .C2 (n_57_97) );
AOI211_X1 g_54_101 (.ZN (n_54_101), .A (n_58_99), .B (n_64_96), .C1 (n_65_93), .C2 (n_59_96) );
AOI211_X1 g_52_102 (.ZN (n_52_102), .A (n_56_100), .B (n_62_97), .C1 (n_66_95), .C2 (n_61_95) );
AOI211_X1 g_50_103 (.ZN (n_50_103), .A (n_54_101), .B (n_60_98), .C1 (n_64_96), .C2 (n_63_94) );
AOI211_X1 g_48_104 (.ZN (n_48_104), .A (n_52_102), .B (n_58_99), .C1 (n_62_97), .C2 (n_65_93) );
AOI211_X1 g_46_103 (.ZN (n_46_103), .A (n_50_103), .B (n_56_100), .C1 (n_60_98), .C2 (n_66_95) );
AOI211_X1 g_44_104 (.ZN (n_44_104), .A (n_48_104), .B (n_54_101), .C1 (n_58_99), .C2 (n_64_96) );
AOI211_X1 g_42_105 (.ZN (n_42_105), .A (n_46_103), .B (n_52_102), .C1 (n_56_100), .C2 (n_62_97) );
AOI211_X1 g_40_106 (.ZN (n_40_106), .A (n_44_104), .B (n_50_103), .C1 (n_54_101), .C2 (n_60_98) );
AOI211_X1 g_38_107 (.ZN (n_38_107), .A (n_42_105), .B (n_48_104), .C1 (n_52_102), .C2 (n_58_99) );
AOI211_X1 g_36_108 (.ZN (n_36_108), .A (n_40_106), .B (n_46_103), .C1 (n_50_103), .C2 (n_56_100) );
AOI211_X1 g_34_109 (.ZN (n_34_109), .A (n_38_107), .B (n_44_104), .C1 (n_48_104), .C2 (n_54_101) );
AOI211_X1 g_32_110 (.ZN (n_32_110), .A (n_36_108), .B (n_42_105), .C1 (n_46_103), .C2 (n_52_102) );
AOI211_X1 g_31_112 (.ZN (n_31_112), .A (n_34_109), .B (n_40_106), .C1 (n_44_104), .C2 (n_50_103) );
AOI211_X1 g_29_111 (.ZN (n_29_111), .A (n_32_110), .B (n_38_107), .C1 (n_42_105), .C2 (n_48_104) );
AOI211_X1 g_31_110 (.ZN (n_31_110), .A (n_31_112), .B (n_36_108), .C1 (n_40_106), .C2 (n_46_103) );
AOI211_X1 g_33_109 (.ZN (n_33_109), .A (n_29_111), .B (n_34_109), .C1 (n_38_107), .C2 (n_44_104) );
AOI211_X1 g_35_108 (.ZN (n_35_108), .A (n_31_110), .B (n_32_110), .C1 (n_36_108), .C2 (n_42_105) );
AOI211_X1 g_37_107 (.ZN (n_37_107), .A (n_33_109), .B (n_31_112), .C1 (n_34_109), .C2 (n_40_106) );
AOI211_X1 g_39_106 (.ZN (n_39_106), .A (n_35_108), .B (n_29_111), .C1 (n_32_110), .C2 (n_38_107) );
AOI211_X1 g_40_108 (.ZN (n_40_108), .A (n_37_107), .B (n_31_110), .C1 (n_31_112), .C2 (n_36_108) );
AOI211_X1 g_38_109 (.ZN (n_38_109), .A (n_39_106), .B (n_33_109), .C1 (n_29_111), .C2 (n_34_109) );
AOI211_X1 g_36_110 (.ZN (n_36_110), .A (n_40_108), .B (n_35_108), .C1 (n_31_110), .C2 (n_32_110) );
AOI211_X1 g_34_111 (.ZN (n_34_111), .A (n_38_109), .B (n_37_107), .C1 (n_33_109), .C2 (n_31_112) );
AOI211_X1 g_35_109 (.ZN (n_35_109), .A (n_36_110), .B (n_39_106), .C1 (n_35_108), .C2 (n_29_111) );
AOI211_X1 g_33_110 (.ZN (n_33_110), .A (n_34_111), .B (n_40_108), .C1 (n_37_107), .C2 (n_31_110) );
AOI211_X1 g_31_111 (.ZN (n_31_111), .A (n_35_109), .B (n_38_109), .C1 (n_39_106), .C2 (n_33_109) );
AOI211_X1 g_30_113 (.ZN (n_30_113), .A (n_33_110), .B (n_36_110), .C1 (n_40_108), .C2 (n_35_108) );
AOI211_X1 g_32_112 (.ZN (n_32_112), .A (n_31_111), .B (n_34_111), .C1 (n_38_109), .C2 (n_37_107) );
AOI211_X1 g_31_114 (.ZN (n_31_114), .A (n_30_113), .B (n_35_109), .C1 (n_36_110), .C2 (n_39_106) );
AOI211_X1 g_30_112 (.ZN (n_30_112), .A (n_32_112), .B (n_33_110), .C1 (n_34_111), .C2 (n_40_108) );
AOI211_X1 g_32_111 (.ZN (n_32_111), .A (n_31_114), .B (n_31_111), .C1 (n_35_109), .C2 (n_38_109) );
AOI211_X1 g_34_110 (.ZN (n_34_110), .A (n_30_112), .B (n_30_113), .C1 (n_33_110), .C2 (n_36_110) );
AOI211_X1 g_36_109 (.ZN (n_36_109), .A (n_32_111), .B (n_32_112), .C1 (n_31_111), .C2 (n_34_111) );
AOI211_X1 g_38_108 (.ZN (n_38_108), .A (n_34_110), .B (n_31_114), .C1 (n_30_113), .C2 (n_35_109) );
AOI211_X1 g_40_107 (.ZN (n_40_107), .A (n_36_109), .B (n_30_112), .C1 (n_32_112), .C2 (n_33_110) );
AOI211_X1 g_39_109 (.ZN (n_39_109), .A (n_38_108), .B (n_32_111), .C1 (n_31_114), .C2 (n_31_111) );
AOI211_X1 g_41_108 (.ZN (n_41_108), .A (n_40_107), .B (n_34_110), .C1 (n_30_112), .C2 (n_30_113) );
AOI211_X1 g_43_107 (.ZN (n_43_107), .A (n_39_109), .B (n_36_109), .C1 (n_32_111), .C2 (n_32_112) );
AOI211_X1 g_45_106 (.ZN (n_45_106), .A (n_41_108), .B (n_38_108), .C1 (n_34_110), .C2 (n_31_114) );
AOI211_X1 g_47_105 (.ZN (n_47_105), .A (n_43_107), .B (n_40_107), .C1 (n_36_109), .C2 (n_30_112) );
AOI211_X1 g_48_103 (.ZN (n_48_103), .A (n_45_106), .B (n_39_109), .C1 (n_38_108), .C2 (n_32_111) );
AOI211_X1 g_50_102 (.ZN (n_50_102), .A (n_47_105), .B (n_41_108), .C1 (n_40_107), .C2 (n_34_110) );
AOI211_X1 g_52_101 (.ZN (n_52_101), .A (n_48_103), .B (n_43_107), .C1 (n_39_109), .C2 (n_36_109) );
AOI211_X1 g_54_100 (.ZN (n_54_100), .A (n_50_102), .B (n_45_106), .C1 (n_41_108), .C2 (n_38_108) );
AOI211_X1 g_56_99 (.ZN (n_56_99), .A (n_52_101), .B (n_47_105), .C1 (n_43_107), .C2 (n_40_107) );
AOI211_X1 g_58_98 (.ZN (n_58_98), .A (n_54_100), .B (n_48_103), .C1 (n_45_106), .C2 (n_39_109) );
AOI211_X1 g_60_97 (.ZN (n_60_97), .A (n_56_99), .B (n_50_102), .C1 (n_47_105), .C2 (n_41_108) );
AOI211_X1 g_62_96 (.ZN (n_62_96), .A (n_58_98), .B (n_52_101), .C1 (n_48_103), .C2 (n_43_107) );
AOI211_X1 g_64_95 (.ZN (n_64_95), .A (n_60_97), .B (n_54_100), .C1 (n_50_102), .C2 (n_45_106) );
AOI211_X1 g_66_94 (.ZN (n_66_94), .A (n_62_96), .B (n_56_99), .C1 (n_52_101), .C2 (n_47_105) );
AOI211_X1 g_68_93 (.ZN (n_68_93), .A (n_64_95), .B (n_58_98), .C1 (n_54_100), .C2 (n_48_103) );
AOI211_X1 g_70_92 (.ZN (n_70_92), .A (n_66_94), .B (n_60_97), .C1 (n_56_99), .C2 (n_50_102) );
AOI211_X1 g_69_94 (.ZN (n_69_94), .A (n_68_93), .B (n_62_96), .C1 (n_58_98), .C2 (n_52_101) );
AOI211_X1 g_71_93 (.ZN (n_71_93), .A (n_70_92), .B (n_64_95), .C1 (n_60_97), .C2 (n_54_100) );
AOI211_X1 g_70_95 (.ZN (n_70_95), .A (n_69_94), .B (n_66_94), .C1 (n_62_96), .C2 (n_56_99) );
AOI211_X1 g_72_94 (.ZN (n_72_94), .A (n_71_93), .B (n_68_93), .C1 (n_64_95), .C2 (n_58_98) );
AOI211_X1 g_71_92 (.ZN (n_71_92), .A (n_70_95), .B (n_70_92), .C1 (n_66_94), .C2 (n_60_97) );
AOI211_X1 g_73_91 (.ZN (n_73_91), .A (n_72_94), .B (n_69_94), .C1 (n_68_93), .C2 (n_62_96) );
AOI211_X1 g_75_90 (.ZN (n_75_90), .A (n_71_92), .B (n_71_93), .C1 (n_70_92), .C2 (n_64_95) );
AOI211_X1 g_77_89 (.ZN (n_77_89), .A (n_73_91), .B (n_70_95), .C1 (n_69_94), .C2 (n_66_94) );
AOI211_X1 g_79_88 (.ZN (n_79_88), .A (n_75_90), .B (n_72_94), .C1 (n_71_93), .C2 (n_68_93) );
AOI211_X1 g_78_90 (.ZN (n_78_90), .A (n_77_89), .B (n_71_92), .C1 (n_70_95), .C2 (n_70_92) );
AOI211_X1 g_80_89 (.ZN (n_80_89), .A (n_79_88), .B (n_73_91), .C1 (n_72_94), .C2 (n_69_94) );
AOI211_X1 g_82_88 (.ZN (n_82_88), .A (n_78_90), .B (n_75_90), .C1 (n_71_92), .C2 (n_71_93) );
AOI211_X1 g_84_87 (.ZN (n_84_87), .A (n_80_89), .B (n_77_89), .C1 (n_73_91), .C2 (n_70_95) );
AOI211_X1 g_86_86 (.ZN (n_86_86), .A (n_82_88), .B (n_79_88), .C1 (n_75_90), .C2 (n_72_94) );
AOI211_X1 g_88_85 (.ZN (n_88_85), .A (n_84_87), .B (n_78_90), .C1 (n_77_89), .C2 (n_71_92) );
AOI211_X1 g_87_87 (.ZN (n_87_87), .A (n_86_86), .B (n_80_89), .C1 (n_79_88), .C2 (n_73_91) );
AOI211_X1 g_89_86 (.ZN (n_89_86), .A (n_88_85), .B (n_82_88), .C1 (n_78_90), .C2 (n_75_90) );
AOI211_X1 g_91_85 (.ZN (n_91_85), .A (n_87_87), .B (n_84_87), .C1 (n_80_89), .C2 (n_77_89) );
AOI211_X1 g_93_84 (.ZN (n_93_84), .A (n_89_86), .B (n_86_86), .C1 (n_82_88), .C2 (n_79_88) );
AOI211_X1 g_95_83 (.ZN (n_95_83), .A (n_91_85), .B (n_88_85), .C1 (n_84_87), .C2 (n_78_90) );
AOI211_X1 g_97_82 (.ZN (n_97_82), .A (n_93_84), .B (n_87_87), .C1 (n_86_86), .C2 (n_80_89) );
AOI211_X1 g_99_81 (.ZN (n_99_81), .A (n_95_83), .B (n_89_86), .C1 (n_88_85), .C2 (n_82_88) );
AOI211_X1 g_101_80 (.ZN (n_101_80), .A (n_97_82), .B (n_91_85), .C1 (n_87_87), .C2 (n_84_87) );
AOI211_X1 g_103_79 (.ZN (n_103_79), .A (n_99_81), .B (n_93_84), .C1 (n_89_86), .C2 (n_86_86) );
AOI211_X1 g_102_81 (.ZN (n_102_81), .A (n_101_80), .B (n_95_83), .C1 (n_91_85), .C2 (n_88_85) );
AOI211_X1 g_104_80 (.ZN (n_104_80), .A (n_103_79), .B (n_97_82), .C1 (n_93_84), .C2 (n_87_87) );
AOI211_X1 g_106_79 (.ZN (n_106_79), .A (n_102_81), .B (n_99_81), .C1 (n_95_83), .C2 (n_89_86) );
AOI211_X1 g_108_78 (.ZN (n_108_78), .A (n_104_80), .B (n_101_80), .C1 (n_97_82), .C2 (n_91_85) );
AOI211_X1 g_110_77 (.ZN (n_110_77), .A (n_106_79), .B (n_103_79), .C1 (n_99_81), .C2 (n_93_84) );
AOI211_X1 g_112_76 (.ZN (n_112_76), .A (n_108_78), .B (n_102_81), .C1 (n_101_80), .C2 (n_95_83) );
AOI211_X1 g_114_75 (.ZN (n_114_75), .A (n_110_77), .B (n_104_80), .C1 (n_103_79), .C2 (n_97_82) );
AOI211_X1 g_116_74 (.ZN (n_116_74), .A (n_112_76), .B (n_106_79), .C1 (n_102_81), .C2 (n_99_81) );
AOI211_X1 g_115_76 (.ZN (n_115_76), .A (n_114_75), .B (n_108_78), .C1 (n_104_80), .C2 (n_101_80) );
AOI211_X1 g_114_74 (.ZN (n_114_74), .A (n_116_74), .B (n_110_77), .C1 (n_106_79), .C2 (n_103_79) );
AOI211_X1 g_116_73 (.ZN (n_116_73), .A (n_115_76), .B (n_112_76), .C1 (n_108_78), .C2 (n_102_81) );
AOI211_X1 g_118_72 (.ZN (n_118_72), .A (n_114_74), .B (n_114_75), .C1 (n_110_77), .C2 (n_104_80) );
AOI211_X1 g_120_71 (.ZN (n_120_71), .A (n_116_73), .B (n_116_74), .C1 (n_112_76), .C2 (n_106_79) );
AOI211_X1 g_122_70 (.ZN (n_122_70), .A (n_118_72), .B (n_115_76), .C1 (n_114_75), .C2 (n_108_78) );
AOI211_X1 g_121_72 (.ZN (n_121_72), .A (n_120_71), .B (n_114_74), .C1 (n_116_74), .C2 (n_110_77) );
AOI211_X1 g_123_71 (.ZN (n_123_71), .A (n_122_70), .B (n_116_73), .C1 (n_115_76), .C2 (n_112_76) );
AOI211_X1 g_125_70 (.ZN (n_125_70), .A (n_121_72), .B (n_118_72), .C1 (n_114_74), .C2 (n_114_75) );
AOI211_X1 g_127_69 (.ZN (n_127_69), .A (n_123_71), .B (n_120_71), .C1 (n_116_73), .C2 (n_116_74) );
AOI211_X1 g_129_68 (.ZN (n_129_68), .A (n_125_70), .B (n_122_70), .C1 (n_118_72), .C2 (n_115_76) );
AOI211_X1 g_131_67 (.ZN (n_131_67), .A (n_127_69), .B (n_121_72), .C1 (n_120_71), .C2 (n_114_74) );
AOI211_X1 g_133_66 (.ZN (n_133_66), .A (n_129_68), .B (n_123_71), .C1 (n_122_70), .C2 (n_116_73) );
AOI211_X1 g_132_68 (.ZN (n_132_68), .A (n_131_67), .B (n_125_70), .C1 (n_121_72), .C2 (n_118_72) );
AOI211_X1 g_130_69 (.ZN (n_130_69), .A (n_133_66), .B (n_127_69), .C1 (n_123_71), .C2 (n_120_71) );
AOI211_X1 g_128_70 (.ZN (n_128_70), .A (n_132_68), .B (n_129_68), .C1 (n_125_70), .C2 (n_122_70) );
AOI211_X1 g_126_71 (.ZN (n_126_71), .A (n_130_69), .B (n_131_67), .C1 (n_127_69), .C2 (n_121_72) );
AOI211_X1 g_124_72 (.ZN (n_124_72), .A (n_128_70), .B (n_133_66), .C1 (n_129_68), .C2 (n_123_71) );
AOI211_X1 g_123_70 (.ZN (n_123_70), .A (n_126_71), .B (n_132_68), .C1 (n_131_67), .C2 (n_125_70) );
AOI211_X1 g_121_71 (.ZN (n_121_71), .A (n_124_72), .B (n_130_69), .C1 (n_133_66), .C2 (n_127_69) );
AOI211_X1 g_119_72 (.ZN (n_119_72), .A (n_123_70), .B (n_128_70), .C1 (n_132_68), .C2 (n_129_68) );
AOI211_X1 g_117_73 (.ZN (n_117_73), .A (n_121_71), .B (n_126_71), .C1 (n_130_69), .C2 (n_131_67) );
AOI211_X1 g_115_74 (.ZN (n_115_74), .A (n_119_72), .B (n_124_72), .C1 (n_128_70), .C2 (n_133_66) );
AOI211_X1 g_113_75 (.ZN (n_113_75), .A (n_117_73), .B (n_123_70), .C1 (n_126_71), .C2 (n_132_68) );
AOI211_X1 g_111_76 (.ZN (n_111_76), .A (n_115_74), .B (n_121_71), .C1 (n_124_72), .C2 (n_130_69) );
AOI211_X1 g_109_77 (.ZN (n_109_77), .A (n_113_75), .B (n_119_72), .C1 (n_123_70), .C2 (n_128_70) );
AOI211_X1 g_107_78 (.ZN (n_107_78), .A (n_111_76), .B (n_117_73), .C1 (n_121_71), .C2 (n_126_71) );
AOI211_X1 g_105_79 (.ZN (n_105_79), .A (n_109_77), .B (n_115_74), .C1 (n_119_72), .C2 (n_124_72) );
AOI211_X1 g_103_80 (.ZN (n_103_80), .A (n_107_78), .B (n_113_75), .C1 (n_117_73), .C2 (n_123_70) );
AOI211_X1 g_101_81 (.ZN (n_101_81), .A (n_105_79), .B (n_111_76), .C1 (n_115_74), .C2 (n_121_71) );
AOI211_X1 g_99_82 (.ZN (n_99_82), .A (n_103_80), .B (n_109_77), .C1 (n_113_75), .C2 (n_119_72) );
AOI211_X1 g_97_81 (.ZN (n_97_81), .A (n_101_81), .B (n_107_78), .C1 (n_111_76), .C2 (n_117_73) );
AOI211_X1 g_95_82 (.ZN (n_95_82), .A (n_99_82), .B (n_105_79), .C1 (n_109_77), .C2 (n_115_74) );
AOI211_X1 g_93_83 (.ZN (n_93_83), .A (n_97_81), .B (n_103_80), .C1 (n_107_78), .C2 (n_113_75) );
AOI211_X1 g_91_84 (.ZN (n_91_84), .A (n_95_82), .B (n_101_81), .C1 (n_105_79), .C2 (n_111_76) );
AOI211_X1 g_89_85 (.ZN (n_89_85), .A (n_93_83), .B (n_99_82), .C1 (n_103_80), .C2 (n_109_77) );
AOI211_X1 g_87_86 (.ZN (n_87_86), .A (n_91_84), .B (n_97_81), .C1 (n_101_81), .C2 (n_107_78) );
AOI211_X1 g_85_87 (.ZN (n_85_87), .A (n_89_85), .B (n_95_82), .C1 (n_99_82), .C2 (n_105_79) );
AOI211_X1 g_83_88 (.ZN (n_83_88), .A (n_87_86), .B (n_93_83), .C1 (n_97_81), .C2 (n_103_80) );
AOI211_X1 g_81_89 (.ZN (n_81_89), .A (n_85_87), .B (n_91_84), .C1 (n_95_82), .C2 (n_101_81) );
AOI211_X1 g_79_90 (.ZN (n_79_90), .A (n_83_88), .B (n_89_85), .C1 (n_93_83), .C2 (n_99_82) );
AOI211_X1 g_77_91 (.ZN (n_77_91), .A (n_81_89), .B (n_87_86), .C1 (n_91_84), .C2 (n_97_81) );
AOI211_X1 g_75_92 (.ZN (n_75_92), .A (n_79_90), .B (n_85_87), .C1 (n_89_85), .C2 (n_95_82) );
AOI211_X1 g_73_93 (.ZN (n_73_93), .A (n_77_91), .B (n_83_88), .C1 (n_87_86), .C2 (n_93_83) );
AOI211_X1 g_71_94 (.ZN (n_71_94), .A (n_75_92), .B (n_81_89), .C1 (n_85_87), .C2 (n_91_84) );
AOI211_X1 g_69_95 (.ZN (n_69_95), .A (n_73_93), .B (n_79_90), .C1 (n_83_88), .C2 (n_89_85) );
AOI211_X1 g_67_94 (.ZN (n_67_94), .A (n_71_94), .B (n_77_91), .C1 (n_81_89), .C2 (n_87_86) );
AOI211_X1 g_65_95 (.ZN (n_65_95), .A (n_69_95), .B (n_75_92), .C1 (n_79_90), .C2 (n_85_87) );
AOI211_X1 g_63_96 (.ZN (n_63_96), .A (n_67_94), .B (n_73_93), .C1 (n_77_91), .C2 (n_83_88) );
AOI211_X1 g_61_97 (.ZN (n_61_97), .A (n_65_95), .B (n_71_94), .C1 (n_75_92), .C2 (n_81_89) );
AOI211_X1 g_59_98 (.ZN (n_59_98), .A (n_63_96), .B (n_69_95), .C1 (n_73_93), .C2 (n_79_90) );
AOI211_X1 g_57_99 (.ZN (n_57_99), .A (n_61_97), .B (n_67_94), .C1 (n_71_94), .C2 (n_77_91) );
AOI211_X1 g_55_100 (.ZN (n_55_100), .A (n_59_98), .B (n_65_95), .C1 (n_69_95), .C2 (n_75_92) );
AOI211_X1 g_53_101 (.ZN (n_53_101), .A (n_57_99), .B (n_63_96), .C1 (n_67_94), .C2 (n_73_93) );
AOI211_X1 g_51_102 (.ZN (n_51_102), .A (n_55_100), .B (n_61_97), .C1 (n_65_95), .C2 (n_71_94) );
AOI211_X1 g_49_103 (.ZN (n_49_103), .A (n_53_101), .B (n_59_98), .C1 (n_63_96), .C2 (n_69_95) );
AOI211_X1 g_47_104 (.ZN (n_47_104), .A (n_51_102), .B (n_57_99), .C1 (n_61_97), .C2 (n_67_94) );
AOI211_X1 g_45_105 (.ZN (n_45_105), .A (n_49_103), .B (n_55_100), .C1 (n_59_98), .C2 (n_65_95) );
AOI211_X1 g_43_106 (.ZN (n_43_106), .A (n_47_104), .B (n_53_101), .C1 (n_57_99), .C2 (n_63_96) );
AOI211_X1 g_41_107 (.ZN (n_41_107), .A (n_45_105), .B (n_51_102), .C1 (n_55_100), .C2 (n_61_97) );
AOI211_X1 g_39_108 (.ZN (n_39_108), .A (n_43_106), .B (n_49_103), .C1 (n_53_101), .C2 (n_59_98) );
AOI211_X1 g_37_109 (.ZN (n_37_109), .A (n_41_107), .B (n_47_104), .C1 (n_51_102), .C2 (n_57_99) );
AOI211_X1 g_35_110 (.ZN (n_35_110), .A (n_39_108), .B (n_45_105), .C1 (n_49_103), .C2 (n_55_100) );
AOI211_X1 g_33_111 (.ZN (n_33_111), .A (n_37_109), .B (n_43_106), .C1 (n_47_104), .C2 (n_53_101) );
AOI211_X1 g_32_113 (.ZN (n_32_113), .A (n_35_110), .B (n_41_107), .C1 (n_45_105), .C2 (n_51_102) );
AOI211_X1 g_34_112 (.ZN (n_34_112), .A (n_33_111), .B (n_39_108), .C1 (n_43_106), .C2 (n_49_103) );
AOI211_X1 g_36_111 (.ZN (n_36_111), .A (n_32_113), .B (n_37_109), .C1 (n_41_107), .C2 (n_47_104) );
AOI211_X1 g_38_110 (.ZN (n_38_110), .A (n_34_112), .B (n_35_110), .C1 (n_39_108), .C2 (n_45_105) );
AOI211_X1 g_40_109 (.ZN (n_40_109), .A (n_36_111), .B (n_33_111), .C1 (n_37_109), .C2 (n_43_106) );
AOI211_X1 g_42_108 (.ZN (n_42_108), .A (n_38_110), .B (n_32_113), .C1 (n_35_110), .C2 (n_41_107) );
AOI211_X1 g_44_107 (.ZN (n_44_107), .A (n_40_109), .B (n_34_112), .C1 (n_33_111), .C2 (n_39_108) );
AOI211_X1 g_46_106 (.ZN (n_46_106), .A (n_42_108), .B (n_36_111), .C1 (n_32_113), .C2 (n_37_109) );
AOI211_X1 g_48_105 (.ZN (n_48_105), .A (n_44_107), .B (n_38_110), .C1 (n_34_112), .C2 (n_35_110) );
AOI211_X1 g_50_104 (.ZN (n_50_104), .A (n_46_106), .B (n_40_109), .C1 (n_36_111), .C2 (n_33_111) );
AOI211_X1 g_52_103 (.ZN (n_52_103), .A (n_48_105), .B (n_42_108), .C1 (n_38_110), .C2 (n_32_113) );
AOI211_X1 g_54_102 (.ZN (n_54_102), .A (n_50_104), .B (n_44_107), .C1 (n_40_109), .C2 (n_34_112) );
AOI211_X1 g_56_101 (.ZN (n_56_101), .A (n_52_103), .B (n_46_106), .C1 (n_42_108), .C2 (n_36_111) );
AOI211_X1 g_58_100 (.ZN (n_58_100), .A (n_54_102), .B (n_48_105), .C1 (n_44_107), .C2 (n_38_110) );
AOI211_X1 g_60_99 (.ZN (n_60_99), .A (n_56_101), .B (n_50_104), .C1 (n_46_106), .C2 (n_40_109) );
AOI211_X1 g_62_98 (.ZN (n_62_98), .A (n_58_100), .B (n_52_103), .C1 (n_48_105), .C2 (n_42_108) );
AOI211_X1 g_64_97 (.ZN (n_64_97), .A (n_60_99), .B (n_54_102), .C1 (n_50_104), .C2 (n_44_107) );
AOI211_X1 g_66_96 (.ZN (n_66_96), .A (n_62_98), .B (n_56_101), .C1 (n_52_103), .C2 (n_46_106) );
AOI211_X1 g_68_95 (.ZN (n_68_95), .A (n_64_97), .B (n_58_100), .C1 (n_54_102), .C2 (n_48_105) );
AOI211_X1 g_70_94 (.ZN (n_70_94), .A (n_66_96), .B (n_60_99), .C1 (n_56_101), .C2 (n_50_104) );
AOI211_X1 g_72_93 (.ZN (n_72_93), .A (n_68_95), .B (n_62_98), .C1 (n_58_100), .C2 (n_52_103) );
AOI211_X1 g_74_92 (.ZN (n_74_92), .A (n_70_94), .B (n_64_97), .C1 (n_60_99), .C2 (n_54_102) );
AOI211_X1 g_76_91 (.ZN (n_76_91), .A (n_72_93), .B (n_66_96), .C1 (n_62_98), .C2 (n_56_101) );
AOI211_X1 g_75_93 (.ZN (n_75_93), .A (n_74_92), .B (n_68_95), .C1 (n_64_97), .C2 (n_58_100) );
AOI211_X1 g_77_92 (.ZN (n_77_92), .A (n_76_91), .B (n_70_94), .C1 (n_66_96), .C2 (n_60_99) );
AOI211_X1 g_79_91 (.ZN (n_79_91), .A (n_75_93), .B (n_72_93), .C1 (n_68_95), .C2 (n_62_98) );
AOI211_X1 g_81_90 (.ZN (n_81_90), .A (n_77_92), .B (n_74_92), .C1 (n_70_94), .C2 (n_64_97) );
AOI211_X1 g_79_89 (.ZN (n_79_89), .A (n_79_91), .B (n_76_91), .C1 (n_72_93), .C2 (n_66_96) );
AOI211_X1 g_81_88 (.ZN (n_81_88), .A (n_81_90), .B (n_75_93), .C1 (n_74_92), .C2 (n_68_95) );
AOI211_X1 g_83_87 (.ZN (n_83_87), .A (n_79_89), .B (n_77_92), .C1 (n_76_91), .C2 (n_70_94) );
AOI211_X1 g_85_88 (.ZN (n_85_88), .A (n_81_88), .B (n_79_91), .C1 (n_75_93), .C2 (n_72_93) );
AOI211_X1 g_83_89 (.ZN (n_83_89), .A (n_83_87), .B (n_81_90), .C1 (n_77_92), .C2 (n_74_92) );
AOI211_X1 g_82_91 (.ZN (n_82_91), .A (n_85_88), .B (n_79_89), .C1 (n_79_91), .C2 (n_76_91) );
AOI211_X1 g_80_90 (.ZN (n_80_90), .A (n_83_89), .B (n_81_88), .C1 (n_81_90), .C2 (n_75_93) );
AOI211_X1 g_82_89 (.ZN (n_82_89), .A (n_82_91), .B (n_83_87), .C1 (n_79_89), .C2 (n_77_92) );
AOI211_X1 g_84_88 (.ZN (n_84_88), .A (n_80_90), .B (n_85_88), .C1 (n_81_88), .C2 (n_79_91) );
AOI211_X1 g_86_87 (.ZN (n_86_87), .A (n_82_89), .B (n_83_89), .C1 (n_83_87), .C2 (n_81_90) );
AOI211_X1 g_88_86 (.ZN (n_88_86), .A (n_84_88), .B (n_82_91), .C1 (n_85_88), .C2 (n_79_89) );
AOI211_X1 g_90_85 (.ZN (n_90_85), .A (n_86_87), .B (n_80_90), .C1 (n_83_89), .C2 (n_81_88) );
AOI211_X1 g_89_87 (.ZN (n_89_87), .A (n_88_86), .B (n_82_89), .C1 (n_82_91), .C2 (n_83_87) );
AOI211_X1 g_91_86 (.ZN (n_91_86), .A (n_90_85), .B (n_84_88), .C1 (n_80_90), .C2 (n_85_88) );
AOI211_X1 g_93_85 (.ZN (n_93_85), .A (n_89_87), .B (n_86_87), .C1 (n_82_89), .C2 (n_83_89) );
AOI211_X1 g_95_84 (.ZN (n_95_84), .A (n_91_86), .B (n_88_86), .C1 (n_84_88), .C2 (n_82_91) );
AOI211_X1 g_97_83 (.ZN (n_97_83), .A (n_93_85), .B (n_90_85), .C1 (n_86_87), .C2 (n_80_90) );
AOI211_X1 g_96_85 (.ZN (n_96_85), .A (n_95_84), .B (n_89_87), .C1 (n_88_86), .C2 (n_82_89) );
AOI211_X1 g_94_84 (.ZN (n_94_84), .A (n_97_83), .B (n_91_86), .C1 (n_90_85), .C2 (n_84_88) );
AOI211_X1 g_96_83 (.ZN (n_96_83), .A (n_96_85), .B (n_93_85), .C1 (n_89_87), .C2 (n_86_87) );
AOI211_X1 g_98_82 (.ZN (n_98_82), .A (n_94_84), .B (n_95_84), .C1 (n_91_86), .C2 (n_88_86) );
AOI211_X1 g_100_81 (.ZN (n_100_81), .A (n_96_83), .B (n_97_83), .C1 (n_93_85), .C2 (n_90_85) );
AOI211_X1 g_102_80 (.ZN (n_102_80), .A (n_98_82), .B (n_96_85), .C1 (n_95_84), .C2 (n_89_87) );
AOI211_X1 g_104_79 (.ZN (n_104_79), .A (n_100_81), .B (n_94_84), .C1 (n_97_83), .C2 (n_91_86) );
AOI211_X1 g_106_78 (.ZN (n_106_78), .A (n_102_80), .B (n_96_83), .C1 (n_96_85), .C2 (n_93_85) );
AOI211_X1 g_108_77 (.ZN (n_108_77), .A (n_104_79), .B (n_98_82), .C1 (n_94_84), .C2 (n_95_84) );
AOI211_X1 g_110_76 (.ZN (n_110_76), .A (n_106_78), .B (n_100_81), .C1 (n_96_83), .C2 (n_97_83) );
AOI211_X1 g_112_75 (.ZN (n_112_75), .A (n_108_77), .B (n_102_80), .C1 (n_98_82), .C2 (n_96_85) );
AOI211_X1 g_113_77 (.ZN (n_113_77), .A (n_110_76), .B (n_104_79), .C1 (n_100_81), .C2 (n_94_84) );
AOI211_X1 g_111_78 (.ZN (n_111_78), .A (n_112_75), .B (n_106_78), .C1 (n_102_80), .C2 (n_96_83) );
AOI211_X1 g_109_79 (.ZN (n_109_79), .A (n_113_77), .B (n_108_77), .C1 (n_104_79), .C2 (n_98_82) );
AOI211_X1 g_107_80 (.ZN (n_107_80), .A (n_111_78), .B (n_110_76), .C1 (n_106_78), .C2 (n_100_81) );
AOI211_X1 g_105_81 (.ZN (n_105_81), .A (n_109_79), .B (n_112_75), .C1 (n_108_77), .C2 (n_102_80) );
AOI211_X1 g_103_82 (.ZN (n_103_82), .A (n_107_80), .B (n_113_77), .C1 (n_110_76), .C2 (n_104_79) );
AOI211_X1 g_101_83 (.ZN (n_101_83), .A (n_105_81), .B (n_111_78), .C1 (n_112_75), .C2 (n_106_78) );
AOI211_X1 g_99_84 (.ZN (n_99_84), .A (n_103_82), .B (n_109_79), .C1 (n_113_77), .C2 (n_108_77) );
AOI211_X1 g_100_82 (.ZN (n_100_82), .A (n_101_83), .B (n_107_80), .C1 (n_111_78), .C2 (n_110_76) );
AOI211_X1 g_98_83 (.ZN (n_98_83), .A (n_99_84), .B (n_105_81), .C1 (n_109_79), .C2 (n_112_75) );
AOI211_X1 g_96_84 (.ZN (n_96_84), .A (n_100_82), .B (n_103_82), .C1 (n_107_80), .C2 (n_113_77) );
AOI211_X1 g_94_85 (.ZN (n_94_85), .A (n_98_83), .B (n_101_83), .C1 (n_105_81), .C2 (n_111_78) );
AOI211_X1 g_92_86 (.ZN (n_92_86), .A (n_96_84), .B (n_99_84), .C1 (n_103_82), .C2 (n_109_79) );
AOI211_X1 g_90_87 (.ZN (n_90_87), .A (n_94_85), .B (n_100_82), .C1 (n_101_83), .C2 (n_107_80) );
AOI211_X1 g_88_88 (.ZN (n_88_88), .A (n_92_86), .B (n_98_83), .C1 (n_99_84), .C2 (n_105_81) );
AOI211_X1 g_86_89 (.ZN (n_86_89), .A (n_90_87), .B (n_96_84), .C1 (n_100_82), .C2 (n_103_82) );
AOI211_X1 g_84_90 (.ZN (n_84_90), .A (n_88_88), .B (n_94_85), .C1 (n_98_83), .C2 (n_101_83) );
AOI211_X1 g_83_92 (.ZN (n_83_92), .A (n_86_89), .B (n_92_86), .C1 (n_96_84), .C2 (n_99_84) );
AOI211_X1 g_82_90 (.ZN (n_82_90), .A (n_84_90), .B (n_90_87), .C1 (n_94_85), .C2 (n_100_82) );
AOI211_X1 g_84_89 (.ZN (n_84_89), .A (n_83_92), .B (n_88_88), .C1 (n_92_86), .C2 (n_98_83) );
AOI211_X1 g_86_88 (.ZN (n_86_88), .A (n_82_90), .B (n_86_89), .C1 (n_90_87), .C2 (n_96_84) );
AOI211_X1 g_88_87 (.ZN (n_88_87), .A (n_84_89), .B (n_84_90), .C1 (n_88_88), .C2 (n_94_85) );
AOI211_X1 g_90_86 (.ZN (n_90_86), .A (n_86_88), .B (n_83_92), .C1 (n_86_89), .C2 (n_92_86) );
AOI211_X1 g_92_85 (.ZN (n_92_85), .A (n_88_87), .B (n_82_90), .C1 (n_84_90), .C2 (n_90_87) );
AOI211_X1 g_94_86 (.ZN (n_94_86), .A (n_90_86), .B (n_84_89), .C1 (n_83_92), .C2 (n_88_88) );
AOI211_X1 g_92_87 (.ZN (n_92_87), .A (n_92_85), .B (n_86_88), .C1 (n_82_90), .C2 (n_86_89) );
AOI211_X1 g_90_88 (.ZN (n_90_88), .A (n_94_86), .B (n_88_87), .C1 (n_84_89), .C2 (n_84_90) );
AOI211_X1 g_88_89 (.ZN (n_88_89), .A (n_92_87), .B (n_90_86), .C1 (n_86_88), .C2 (n_83_92) );
AOI211_X1 g_86_90 (.ZN (n_86_90), .A (n_90_88), .B (n_92_85), .C1 (n_88_87), .C2 (n_82_90) );
AOI211_X1 g_87_88 (.ZN (n_87_88), .A (n_88_89), .B (n_94_86), .C1 (n_90_86), .C2 (n_84_89) );
AOI211_X1 g_85_89 (.ZN (n_85_89), .A (n_86_90), .B (n_92_87), .C1 (n_92_85), .C2 (n_86_88) );
AOI211_X1 g_83_90 (.ZN (n_83_90), .A (n_87_88), .B (n_90_88), .C1 (n_94_86), .C2 (n_88_87) );
AOI211_X1 g_81_91 (.ZN (n_81_91), .A (n_85_89), .B (n_88_89), .C1 (n_92_87), .C2 (n_90_86) );
AOI211_X1 g_79_92 (.ZN (n_79_92), .A (n_83_90), .B (n_86_90), .C1 (n_90_88), .C2 (n_92_85) );
AOI211_X1 g_77_93 (.ZN (n_77_93), .A (n_81_91), .B (n_87_88), .C1 (n_88_89), .C2 (n_94_86) );
AOI211_X1 g_78_91 (.ZN (n_78_91), .A (n_79_92), .B (n_85_89), .C1 (n_86_90), .C2 (n_92_87) );
AOI211_X1 g_76_92 (.ZN (n_76_92), .A (n_77_93), .B (n_83_90), .C1 (n_87_88), .C2 (n_90_88) );
AOI211_X1 g_74_93 (.ZN (n_74_93), .A (n_78_91), .B (n_81_91), .C1 (n_85_89), .C2 (n_88_89) );
AOI211_X1 g_73_95 (.ZN (n_73_95), .A (n_76_92), .B (n_79_92), .C1 (n_83_90), .C2 (n_86_90) );
AOI211_X1 g_75_94 (.ZN (n_75_94), .A (n_74_93), .B (n_77_93), .C1 (n_81_91), .C2 (n_87_88) );
AOI211_X1 g_74_96 (.ZN (n_74_96), .A (n_73_95), .B (n_78_91), .C1 (n_79_92), .C2 (n_85_89) );
AOI211_X1 g_73_94 (.ZN (n_73_94), .A (n_75_94), .B (n_76_92), .C1 (n_77_93), .C2 (n_83_90) );
AOI211_X1 g_71_95 (.ZN (n_71_95), .A (n_74_96), .B (n_74_93), .C1 (n_78_91), .C2 (n_81_91) );
AOI211_X1 g_69_96 (.ZN (n_69_96), .A (n_73_94), .B (n_73_95), .C1 (n_76_92), .C2 (n_79_92) );
AOI211_X1 g_67_95 (.ZN (n_67_95), .A (n_71_95), .B (n_75_94), .C1 (n_74_93), .C2 (n_77_93) );
AOI211_X1 g_65_96 (.ZN (n_65_96), .A (n_69_96), .B (n_74_96), .C1 (n_73_95), .C2 (n_78_91) );
AOI211_X1 g_63_97 (.ZN (n_63_97), .A (n_67_95), .B (n_73_94), .C1 (n_75_94), .C2 (n_76_92) );
AOI211_X1 g_61_98 (.ZN (n_61_98), .A (n_65_96), .B (n_71_95), .C1 (n_74_96), .C2 (n_74_93) );
AOI211_X1 g_59_99 (.ZN (n_59_99), .A (n_63_97), .B (n_69_96), .C1 (n_73_94), .C2 (n_73_95) );
AOI211_X1 g_57_100 (.ZN (n_57_100), .A (n_61_98), .B (n_67_95), .C1 (n_71_95), .C2 (n_75_94) );
AOI211_X1 g_55_101 (.ZN (n_55_101), .A (n_59_99), .B (n_65_96), .C1 (n_69_96), .C2 (n_74_96) );
AOI211_X1 g_53_102 (.ZN (n_53_102), .A (n_57_100), .B (n_63_97), .C1 (n_67_95), .C2 (n_73_94) );
AOI211_X1 g_51_103 (.ZN (n_51_103), .A (n_55_101), .B (n_61_98), .C1 (n_65_96), .C2 (n_71_95) );
AOI211_X1 g_49_104 (.ZN (n_49_104), .A (n_53_102), .B (n_59_99), .C1 (n_63_97), .C2 (n_69_96) );
AOI211_X1 g_51_105 (.ZN (n_51_105), .A (n_51_103), .B (n_57_100), .C1 (n_61_98), .C2 (n_67_95) );
AOI211_X1 g_53_104 (.ZN (n_53_104), .A (n_49_104), .B (n_55_101), .C1 (n_59_99), .C2 (n_65_96) );
AOI211_X1 g_55_103 (.ZN (n_55_103), .A (n_51_105), .B (n_53_102), .C1 (n_57_100), .C2 (n_63_97) );
AOI211_X1 g_57_102 (.ZN (n_57_102), .A (n_53_104), .B (n_51_103), .C1 (n_55_101), .C2 (n_61_98) );
AOI211_X1 g_59_101 (.ZN (n_59_101), .A (n_55_103), .B (n_49_104), .C1 (n_53_102), .C2 (n_59_99) );
AOI211_X1 g_61_100 (.ZN (n_61_100), .A (n_57_102), .B (n_51_105), .C1 (n_51_103), .C2 (n_57_100) );
AOI211_X1 g_63_99 (.ZN (n_63_99), .A (n_59_101), .B (n_53_104), .C1 (n_49_104), .C2 (n_55_101) );
AOI211_X1 g_65_98 (.ZN (n_65_98), .A (n_61_100), .B (n_55_103), .C1 (n_51_105), .C2 (n_53_102) );
AOI211_X1 g_67_97 (.ZN (n_67_97), .A (n_63_99), .B (n_57_102), .C1 (n_53_104), .C2 (n_51_103) );
AOI211_X1 g_66_99 (.ZN (n_66_99), .A (n_65_98), .B (n_59_101), .C1 (n_55_103), .C2 (n_49_104) );
AOI211_X1 g_65_97 (.ZN (n_65_97), .A (n_67_97), .B (n_61_100), .C1 (n_57_102), .C2 (n_51_105) );
AOI211_X1 g_67_96 (.ZN (n_67_96), .A (n_66_99), .B (n_63_99), .C1 (n_59_101), .C2 (n_53_104) );
AOI211_X1 g_66_98 (.ZN (n_66_98), .A (n_65_97), .B (n_65_98), .C1 (n_61_100), .C2 (n_55_103) );
AOI211_X1 g_68_97 (.ZN (n_68_97), .A (n_67_96), .B (n_67_97), .C1 (n_63_99), .C2 (n_57_102) );
AOI211_X1 g_70_96 (.ZN (n_70_96), .A (n_66_98), .B (n_66_99), .C1 (n_65_98), .C2 (n_59_101) );
AOI211_X1 g_72_95 (.ZN (n_72_95), .A (n_68_97), .B (n_65_97), .C1 (n_67_97), .C2 (n_61_100) );
AOI211_X1 g_74_94 (.ZN (n_74_94), .A (n_70_96), .B (n_67_96), .C1 (n_66_99), .C2 (n_63_99) );
AOI211_X1 g_76_93 (.ZN (n_76_93), .A (n_72_95), .B (n_66_98), .C1 (n_65_97), .C2 (n_65_98) );
AOI211_X1 g_78_92 (.ZN (n_78_92), .A (n_74_94), .B (n_68_97), .C1 (n_67_96), .C2 (n_67_97) );
AOI211_X1 g_80_91 (.ZN (n_80_91), .A (n_76_93), .B (n_70_96), .C1 (n_66_98), .C2 (n_66_99) );
AOI211_X1 g_81_93 (.ZN (n_81_93), .A (n_78_92), .B (n_72_95), .C1 (n_68_97), .C2 (n_65_97) );
AOI211_X1 g_79_94 (.ZN (n_79_94), .A (n_80_91), .B (n_74_94), .C1 (n_70_96), .C2 (n_67_96) );
AOI211_X1 g_80_92 (.ZN (n_80_92), .A (n_81_93), .B (n_76_93), .C1 (n_72_95), .C2 (n_66_98) );
AOI211_X1 g_78_93 (.ZN (n_78_93), .A (n_79_94), .B (n_78_92), .C1 (n_74_94), .C2 (n_68_97) );
AOI211_X1 g_76_94 (.ZN (n_76_94), .A (n_80_92), .B (n_80_91), .C1 (n_76_93), .C2 (n_70_96) );
AOI211_X1 g_74_95 (.ZN (n_74_95), .A (n_78_93), .B (n_81_93), .C1 (n_78_92), .C2 (n_72_95) );
AOI211_X1 g_72_96 (.ZN (n_72_96), .A (n_76_94), .B (n_79_94), .C1 (n_80_91), .C2 (n_74_94) );
AOI211_X1 g_70_97 (.ZN (n_70_97), .A (n_74_95), .B (n_80_92), .C1 (n_81_93), .C2 (n_76_93) );
AOI211_X1 g_68_96 (.ZN (n_68_96), .A (n_72_96), .B (n_78_93), .C1 (n_79_94), .C2 (n_78_92) );
AOI211_X1 g_66_97 (.ZN (n_66_97), .A (n_70_97), .B (n_76_94), .C1 (n_80_92), .C2 (n_80_91) );
AOI211_X1 g_64_98 (.ZN (n_64_98), .A (n_68_96), .B (n_74_95), .C1 (n_78_93), .C2 (n_81_93) );
AOI211_X1 g_62_99 (.ZN (n_62_99), .A (n_66_97), .B (n_72_96), .C1 (n_76_94), .C2 (n_79_94) );
AOI211_X1 g_60_100 (.ZN (n_60_100), .A (n_64_98), .B (n_70_97), .C1 (n_74_95), .C2 (n_80_92) );
AOI211_X1 g_58_101 (.ZN (n_58_101), .A (n_62_99), .B (n_68_96), .C1 (n_72_96), .C2 (n_78_93) );
AOI211_X1 g_56_102 (.ZN (n_56_102), .A (n_60_100), .B (n_66_97), .C1 (n_70_97), .C2 (n_76_94) );
AOI211_X1 g_54_103 (.ZN (n_54_103), .A (n_58_101), .B (n_64_98), .C1 (n_68_96), .C2 (n_74_95) );
AOI211_X1 g_52_104 (.ZN (n_52_104), .A (n_56_102), .B (n_62_99), .C1 (n_66_97), .C2 (n_72_96) );
AOI211_X1 g_50_105 (.ZN (n_50_105), .A (n_54_103), .B (n_60_100), .C1 (n_64_98), .C2 (n_70_97) );
AOI211_X1 g_48_106 (.ZN (n_48_106), .A (n_52_104), .B (n_58_101), .C1 (n_62_99), .C2 (n_68_96) );
AOI211_X1 g_46_105 (.ZN (n_46_105), .A (n_50_105), .B (n_56_102), .C1 (n_60_100), .C2 (n_66_97) );
AOI211_X1 g_44_106 (.ZN (n_44_106), .A (n_48_106), .B (n_54_103), .C1 (n_58_101), .C2 (n_64_98) );
AOI211_X1 g_46_107 (.ZN (n_46_107), .A (n_46_105), .B (n_52_104), .C1 (n_56_102), .C2 (n_62_99) );
AOI211_X1 g_44_108 (.ZN (n_44_108), .A (n_44_106), .B (n_50_105), .C1 (n_54_103), .C2 (n_60_100) );
AOI211_X1 g_42_109 (.ZN (n_42_109), .A (n_46_107), .B (n_48_106), .C1 (n_52_104), .C2 (n_58_101) );
AOI211_X1 g_40_110 (.ZN (n_40_110), .A (n_44_108), .B (n_46_105), .C1 (n_50_105), .C2 (n_56_102) );
AOI211_X1 g_38_111 (.ZN (n_38_111), .A (n_42_109), .B (n_44_106), .C1 (n_48_106), .C2 (n_54_103) );
AOI211_X1 g_36_112 (.ZN (n_36_112), .A (n_40_110), .B (n_46_107), .C1 (n_46_105), .C2 (n_52_104) );
AOI211_X1 g_37_110 (.ZN (n_37_110), .A (n_38_111), .B (n_44_108), .C1 (n_44_106), .C2 (n_50_105) );
AOI211_X1 g_35_111 (.ZN (n_35_111), .A (n_36_112), .B (n_42_109), .C1 (n_46_107), .C2 (n_48_106) );
AOI211_X1 g_33_112 (.ZN (n_33_112), .A (n_37_110), .B (n_40_110), .C1 (n_44_108), .C2 (n_46_105) );
AOI211_X1 g_31_113 (.ZN (n_31_113), .A (n_35_111), .B (n_38_111), .C1 (n_42_109), .C2 (n_44_106) );
AOI211_X1 g_29_114 (.ZN (n_29_114), .A (n_33_112), .B (n_36_112), .C1 (n_40_110), .C2 (n_46_107) );
AOI211_X1 g_27_115 (.ZN (n_27_115), .A (n_31_113), .B (n_37_110), .C1 (n_38_111), .C2 (n_44_108) );
AOI211_X1 g_28_113 (.ZN (n_28_113), .A (n_29_114), .B (n_35_111), .C1 (n_36_112), .C2 (n_42_109) );
AOI211_X1 g_30_114 (.ZN (n_30_114), .A (n_27_115), .B (n_33_112), .C1 (n_37_110), .C2 (n_40_110) );
AOI211_X1 g_28_115 (.ZN (n_28_115), .A (n_28_113), .B (n_31_113), .C1 (n_35_111), .C2 (n_38_111) );
AOI211_X1 g_29_113 (.ZN (n_29_113), .A (n_30_114), .B (n_29_114), .C1 (n_33_112), .C2 (n_36_112) );
AOI211_X1 g_27_112 (.ZN (n_27_112), .A (n_28_115), .B (n_27_115), .C1 (n_31_113), .C2 (n_37_110) );
AOI211_X1 g_26_114 (.ZN (n_26_114), .A (n_29_113), .B (n_28_113), .C1 (n_29_114), .C2 (n_35_111) );
AOI211_X1 g_25_116 (.ZN (n_25_116), .A (n_27_112), .B (n_30_114), .C1 (n_27_115), .C2 (n_33_112) );
AOI211_X1 g_24_114 (.ZN (n_24_114), .A (n_26_114), .B (n_28_115), .C1 (n_28_113), .C2 (n_31_113) );
AOI211_X1 g_22_115 (.ZN (n_22_115), .A (n_25_116), .B (n_29_113), .C1 (n_30_114), .C2 (n_29_114) );
AOI211_X1 g_21_113 (.ZN (n_21_113), .A (n_24_114), .B (n_27_112), .C1 (n_28_115), .C2 (n_27_115) );
AOI211_X1 g_19_114 (.ZN (n_19_114), .A (n_22_115), .B (n_26_114), .C1 (n_29_113), .C2 (n_28_113) );
AOI211_X1 g_17_115 (.ZN (n_17_115), .A (n_21_113), .B (n_25_116), .C1 (n_27_112), .C2 (n_30_114) );
AOI211_X1 g_15_116 (.ZN (n_15_116), .A (n_19_114), .B (n_24_114), .C1 (n_26_114), .C2 (n_28_115) );
AOI211_X1 g_13_117 (.ZN (n_13_117), .A (n_17_115), .B (n_22_115), .C1 (n_25_116), .C2 (n_29_113) );
AOI211_X1 g_11_118 (.ZN (n_11_118), .A (n_15_116), .B (n_21_113), .C1 (n_24_114), .C2 (n_27_112) );
AOI211_X1 g_9_119 (.ZN (n_9_119), .A (n_13_117), .B (n_19_114), .C1 (n_22_115), .C2 (n_26_114) );
AOI211_X1 g_7_120 (.ZN (n_7_120), .A (n_11_118), .B (n_17_115), .C1 (n_21_113), .C2 (n_25_116) );
AOI211_X1 g_6_122 (.ZN (n_6_122), .A (n_9_119), .B (n_15_116), .C1 (n_19_114), .C2 (n_24_114) );
AOI211_X1 g_8_121 (.ZN (n_8_121), .A (n_7_120), .B (n_13_117), .C1 (n_17_115), .C2 (n_22_115) );
AOI211_X1 g_10_120 (.ZN (n_10_120), .A (n_6_122), .B (n_11_118), .C1 (n_15_116), .C2 (n_21_113) );
AOI211_X1 g_12_119 (.ZN (n_12_119), .A (n_8_121), .B (n_9_119), .C1 (n_13_117), .C2 (n_19_114) );
AOI211_X1 g_14_118 (.ZN (n_14_118), .A (n_10_120), .B (n_7_120), .C1 (n_11_118), .C2 (n_17_115) );
AOI211_X1 g_16_117 (.ZN (n_16_117), .A (n_12_119), .B (n_6_122), .C1 (n_9_119), .C2 (n_15_116) );
AOI211_X1 g_18_116 (.ZN (n_18_116), .A (n_14_118), .B (n_8_121), .C1 (n_7_120), .C2 (n_13_117) );
AOI211_X1 g_20_115 (.ZN (n_20_115), .A (n_16_117), .B (n_10_120), .C1 (n_6_122), .C2 (n_11_118) );
AOI211_X1 g_22_114 (.ZN (n_22_114), .A (n_18_116), .B (n_12_119), .C1 (n_8_121), .C2 (n_9_119) );
AOI211_X1 g_21_116 (.ZN (n_21_116), .A (n_20_115), .B (n_14_118), .C1 (n_10_120), .C2 (n_7_120) );
AOI211_X1 g_20_114 (.ZN (n_20_114), .A (n_22_114), .B (n_16_117), .C1 (n_12_119), .C2 (n_6_122) );
AOI211_X1 g_18_115 (.ZN (n_18_115), .A (n_21_116), .B (n_18_116), .C1 (n_14_118), .C2 (n_8_121) );
AOI211_X1 g_19_117 (.ZN (n_19_117), .A (n_20_114), .B (n_20_115), .C1 (n_16_117), .C2 (n_10_120) );
AOI211_X1 g_17_118 (.ZN (n_17_118), .A (n_18_115), .B (n_22_114), .C1 (n_18_116), .C2 (n_12_119) );
AOI211_X1 g_15_119 (.ZN (n_15_119), .A (n_19_117), .B (n_21_116), .C1 (n_20_115), .C2 (n_14_118) );
AOI211_X1 g_13_118 (.ZN (n_13_118), .A (n_17_118), .B (n_20_114), .C1 (n_22_114), .C2 (n_16_117) );
AOI211_X1 g_11_119 (.ZN (n_11_119), .A (n_15_119), .B (n_18_115), .C1 (n_21_116), .C2 (n_18_116) );
AOI211_X1 g_9_120 (.ZN (n_9_120), .A (n_13_118), .B (n_19_117), .C1 (n_20_114), .C2 (n_20_115) );
AOI211_X1 g_8_122 (.ZN (n_8_122), .A (n_11_119), .B (n_17_118), .C1 (n_18_115), .C2 (n_22_114) );
AOI211_X1 g_6_123 (.ZN (n_6_123), .A (n_9_120), .B (n_15_119), .C1 (n_19_117), .C2 (n_21_116) );
AOI211_X1 g_5_125 (.ZN (n_5_125), .A (n_8_122), .B (n_13_118), .C1 (n_17_118), .C2 (n_20_114) );
AOI211_X1 g_7_124 (.ZN (n_7_124), .A (n_6_123), .B (n_11_119), .C1 (n_15_119), .C2 (n_18_115) );
AOI211_X1 g_9_123 (.ZN (n_9_123), .A (n_5_125), .B (n_9_120), .C1 (n_13_118), .C2 (n_19_117) );
AOI211_X1 g_10_121 (.ZN (n_10_121), .A (n_7_124), .B (n_8_122), .C1 (n_11_119), .C2 (n_17_118) );
AOI211_X1 g_12_120 (.ZN (n_12_120), .A (n_9_123), .B (n_6_123), .C1 (n_9_120), .C2 (n_15_119) );
AOI211_X1 g_14_119 (.ZN (n_14_119), .A (n_10_121), .B (n_5_125), .C1 (n_8_122), .C2 (n_13_118) );
AOI211_X1 g_16_118 (.ZN (n_16_118), .A (n_12_120), .B (n_7_124), .C1 (n_6_123), .C2 (n_11_119) );
AOI211_X1 g_18_117 (.ZN (n_18_117), .A (n_14_119), .B (n_9_123), .C1 (n_5_125), .C2 (n_9_120) );
AOI211_X1 g_20_116 (.ZN (n_20_116), .A (n_16_118), .B (n_10_121), .C1 (n_7_124), .C2 (n_8_122) );
AOI211_X1 g_19_118 (.ZN (n_19_118), .A (n_18_117), .B (n_12_120), .C1 (n_9_123), .C2 (n_6_123) );
AOI211_X1 g_17_117 (.ZN (n_17_117), .A (n_20_116), .B (n_14_119), .C1 (n_10_121), .C2 (n_5_125) );
AOI211_X1 g_15_118 (.ZN (n_15_118), .A (n_19_118), .B (n_16_118), .C1 (n_12_120), .C2 (n_7_124) );
AOI211_X1 g_17_119 (.ZN (n_17_119), .A (n_17_117), .B (n_18_117), .C1 (n_14_119), .C2 (n_9_123) );
AOI211_X1 g_15_120 (.ZN (n_15_120), .A (n_15_118), .B (n_20_116), .C1 (n_16_118), .C2 (n_10_121) );
AOI211_X1 g_13_121 (.ZN (n_13_121), .A (n_17_119), .B (n_19_118), .C1 (n_18_117), .C2 (n_12_120) );
AOI211_X1 g_11_120 (.ZN (n_11_120), .A (n_15_120), .B (n_17_117), .C1 (n_20_116), .C2 (n_14_119) );
AOI211_X1 g_9_121 (.ZN (n_9_121), .A (n_13_121), .B (n_15_118), .C1 (n_19_118), .C2 (n_16_118) );
AOI211_X1 g_11_122 (.ZN (n_11_122), .A (n_11_120), .B (n_17_119), .C1 (n_17_117), .C2 (n_18_117) );
AOI211_X1 g_10_124 (.ZN (n_10_124), .A (n_9_121), .B (n_15_120), .C1 (n_15_118), .C2 (n_20_116) );
AOI211_X1 g_8_123 (.ZN (n_8_123), .A (n_11_122), .B (n_13_121), .C1 (n_17_119), .C2 (n_19_118) );
AOI211_X1 g_10_122 (.ZN (n_10_122), .A (n_10_124), .B (n_11_120), .C1 (n_15_120), .C2 (n_17_117) );
AOI211_X1 g_12_121 (.ZN (n_12_121), .A (n_8_123), .B (n_9_121), .C1 (n_13_121), .C2 (n_15_118) );
AOI211_X1 g_14_120 (.ZN (n_14_120), .A (n_10_122), .B (n_11_122), .C1 (n_11_120), .C2 (n_17_119) );
AOI211_X1 g_16_119 (.ZN (n_16_119), .A (n_12_121), .B (n_10_124), .C1 (n_9_121), .C2 (n_15_120) );
AOI211_X1 g_18_118 (.ZN (n_18_118), .A (n_14_120), .B (n_8_123), .C1 (n_11_122), .C2 (n_13_121) );
AOI211_X1 g_19_116 (.ZN (n_19_116), .A (n_16_119), .B (n_10_122), .C1 (n_10_124), .C2 (n_11_120) );
AOI211_X1 g_21_115 (.ZN (n_21_115), .A (n_18_118), .B (n_12_121), .C1 (n_8_123), .C2 (n_9_121) );
AOI211_X1 g_23_114 (.ZN (n_23_114), .A (n_19_116), .B (n_14_120), .C1 (n_10_122), .C2 (n_11_122) );
AOI211_X1 g_25_113 (.ZN (n_25_113), .A (n_21_115), .B (n_16_119), .C1 (n_12_121), .C2 (n_10_124) );
AOI211_X1 g_24_115 (.ZN (n_24_115), .A (n_23_114), .B (n_18_118), .C1 (n_14_120), .C2 (n_8_123) );
AOI211_X1 g_22_116 (.ZN (n_22_116), .A (n_25_113), .B (n_19_116), .C1 (n_16_119), .C2 (n_10_122) );
AOI211_X1 g_20_117 (.ZN (n_20_117), .A (n_24_115), .B (n_21_115), .C1 (n_18_118), .C2 (n_12_121) );
AOI211_X1 g_19_119 (.ZN (n_19_119), .A (n_22_116), .B (n_23_114), .C1 (n_19_116), .C2 (n_14_120) );
AOI211_X1 g_21_118 (.ZN (n_21_118), .A (n_20_117), .B (n_25_113), .C1 (n_21_115), .C2 (n_16_119) );
AOI211_X1 g_23_117 (.ZN (n_23_117), .A (n_19_119), .B (n_24_115), .C1 (n_23_114), .C2 (n_18_118) );
AOI211_X1 g_22_119 (.ZN (n_22_119), .A (n_21_118), .B (n_22_116), .C1 (n_25_113), .C2 (n_19_116) );
AOI211_X1 g_21_117 (.ZN (n_21_117), .A (n_23_117), .B (n_20_117), .C1 (n_24_115), .C2 (n_21_115) );
AOI211_X1 g_23_116 (.ZN (n_23_116), .A (n_22_119), .B (n_19_119), .C1 (n_22_116), .C2 (n_23_114) );
AOI211_X1 g_25_115 (.ZN (n_25_115), .A (n_21_117), .B (n_21_118), .C1 (n_20_117), .C2 (n_25_113) );
AOI211_X1 g_27_114 (.ZN (n_27_114), .A (n_23_116), .B (n_23_117), .C1 (n_19_119), .C2 (n_24_115) );
AOI211_X1 g_26_116 (.ZN (n_26_116), .A (n_25_115), .B (n_22_119), .C1 (n_21_118), .C2 (n_22_116) );
AOI211_X1 g_24_117 (.ZN (n_24_117), .A (n_27_114), .B (n_21_117), .C1 (n_23_117), .C2 (n_20_117) );
AOI211_X1 g_22_118 (.ZN (n_22_118), .A (n_26_116), .B (n_23_116), .C1 (n_22_119), .C2 (n_19_119) );
AOI211_X1 g_20_119 (.ZN (n_20_119), .A (n_24_117), .B (n_25_115), .C1 (n_21_117), .C2 (n_21_118) );
AOI211_X1 g_18_120 (.ZN (n_18_120), .A (n_22_118), .B (n_27_114), .C1 (n_23_116), .C2 (n_23_117) );
AOI211_X1 g_16_121 (.ZN (n_16_121), .A (n_20_119), .B (n_26_116), .C1 (n_25_115), .C2 (n_22_119) );
AOI211_X1 g_14_122 (.ZN (n_14_122), .A (n_18_120), .B (n_24_117), .C1 (n_27_114), .C2 (n_21_117) );
AOI211_X1 g_13_120 (.ZN (n_13_120), .A (n_16_121), .B (n_22_118), .C1 (n_26_116), .C2 (n_23_116) );
AOI211_X1 g_11_121 (.ZN (n_11_121), .A (n_14_122), .B (n_20_119), .C1 (n_24_117), .C2 (n_25_115) );
AOI211_X1 g_9_122 (.ZN (n_9_122), .A (n_13_120), .B (n_18_120), .C1 (n_22_118), .C2 (n_27_114) );
AOI211_X1 g_7_123 (.ZN (n_7_123), .A (n_11_121), .B (n_16_121), .C1 (n_20_119), .C2 (n_26_116) );
AOI211_X1 g_5_124 (.ZN (n_5_124), .A (n_9_122), .B (n_14_122), .C1 (n_18_120), .C2 (n_24_117) );
AOI211_X1 g_4_126 (.ZN (n_4_126), .A (n_7_123), .B (n_13_120), .C1 (n_16_121), .C2 (n_22_118) );
AOI211_X1 g_6_125 (.ZN (n_6_125), .A (n_5_124), .B (n_11_121), .C1 (n_14_122), .C2 (n_20_119) );
AOI211_X1 g_8_124 (.ZN (n_8_124), .A (n_4_126), .B (n_9_122), .C1 (n_13_120), .C2 (n_18_120) );
AOI211_X1 g_10_123 (.ZN (n_10_123), .A (n_6_125), .B (n_7_123), .C1 (n_11_121), .C2 (n_16_121) );
AOI211_X1 g_12_122 (.ZN (n_12_122), .A (n_8_124), .B (n_5_124), .C1 (n_9_122), .C2 (n_14_122) );
AOI211_X1 g_14_121 (.ZN (n_14_121), .A (n_10_123), .B (n_4_126), .C1 (n_7_123), .C2 (n_13_120) );
AOI211_X1 g_16_120 (.ZN (n_16_120), .A (n_12_122), .B (n_6_125), .C1 (n_5_124), .C2 (n_11_121) );
AOI211_X1 g_18_119 (.ZN (n_18_119), .A (n_14_121), .B (n_8_124), .C1 (n_4_126), .C2 (n_9_122) );
AOI211_X1 g_20_118 (.ZN (n_20_118), .A (n_16_120), .B (n_10_123), .C1 (n_6_125), .C2 (n_7_123) );
AOI211_X1 g_22_117 (.ZN (n_22_117), .A (n_18_119), .B (n_12_122), .C1 (n_8_124), .C2 (n_5_124) );
AOI211_X1 g_24_116 (.ZN (n_24_116), .A (n_20_118), .B (n_14_121), .C1 (n_10_123), .C2 (n_4_126) );
AOI211_X1 g_26_115 (.ZN (n_26_115), .A (n_22_117), .B (n_16_120), .C1 (n_12_122), .C2 (n_6_125) );
AOI211_X1 g_28_114 (.ZN (n_28_114), .A (n_24_116), .B (n_18_119), .C1 (n_14_121), .C2 (n_8_124) );
AOI211_X1 g_27_116 (.ZN (n_27_116), .A (n_26_115), .B (n_20_118), .C1 (n_16_120), .C2 (n_10_123) );
AOI211_X1 g_29_115 (.ZN (n_29_115), .A (n_28_114), .B (n_22_117), .C1 (n_18_119), .C2 (n_12_122) );
AOI211_X1 g_28_117 (.ZN (n_28_117), .A (n_27_116), .B (n_24_116), .C1 (n_20_118), .C2 (n_14_121) );
AOI211_X1 g_30_116 (.ZN (n_30_116), .A (n_29_115), .B (n_26_115), .C1 (n_22_117), .C2 (n_16_120) );
AOI211_X1 g_32_115 (.ZN (n_32_115), .A (n_28_117), .B (n_28_114), .C1 (n_24_116), .C2 (n_18_119) );
AOI211_X1 g_33_113 (.ZN (n_33_113), .A (n_30_116), .B (n_27_116), .C1 (n_26_115), .C2 (n_20_118) );
AOI211_X1 g_35_112 (.ZN (n_35_112), .A (n_32_115), .B (n_29_115), .C1 (n_28_114), .C2 (n_22_117) );
AOI211_X1 g_37_111 (.ZN (n_37_111), .A (n_33_113), .B (n_28_117), .C1 (n_27_116), .C2 (n_24_116) );
AOI211_X1 g_39_110 (.ZN (n_39_110), .A (n_35_112), .B (n_30_116), .C1 (n_29_115), .C2 (n_26_115) );
AOI211_X1 g_41_109 (.ZN (n_41_109), .A (n_37_111), .B (n_32_115), .C1 (n_28_117), .C2 (n_28_114) );
AOI211_X1 g_43_108 (.ZN (n_43_108), .A (n_39_110), .B (n_33_113), .C1 (n_30_116), .C2 (n_27_116) );
AOI211_X1 g_45_107 (.ZN (n_45_107), .A (n_41_109), .B (n_35_112), .C1 (n_32_115), .C2 (n_29_115) );
AOI211_X1 g_47_106 (.ZN (n_47_106), .A (n_43_108), .B (n_37_111), .C1 (n_33_113), .C2 (n_28_117) );
AOI211_X1 g_49_105 (.ZN (n_49_105), .A (n_45_107), .B (n_39_110), .C1 (n_35_112), .C2 (n_30_116) );
AOI211_X1 g_51_104 (.ZN (n_51_104), .A (n_47_106), .B (n_41_109), .C1 (n_37_111), .C2 (n_32_115) );
AOI211_X1 g_53_103 (.ZN (n_53_103), .A (n_49_105), .B (n_43_108), .C1 (n_39_110), .C2 (n_33_113) );
AOI211_X1 g_55_102 (.ZN (n_55_102), .A (n_51_104), .B (n_45_107), .C1 (n_41_109), .C2 (n_35_112) );
AOI211_X1 g_57_101 (.ZN (n_57_101), .A (n_53_103), .B (n_47_106), .C1 (n_43_108), .C2 (n_37_111) );
AOI211_X1 g_59_100 (.ZN (n_59_100), .A (n_55_102), .B (n_49_105), .C1 (n_45_107), .C2 (n_39_110) );
AOI211_X1 g_61_99 (.ZN (n_61_99), .A (n_57_101), .B (n_51_104), .C1 (n_47_106), .C2 (n_41_109) );
AOI211_X1 g_63_98 (.ZN (n_63_98), .A (n_59_100), .B (n_53_103), .C1 (n_49_105), .C2 (n_43_108) );
AOI211_X1 g_64_100 (.ZN (n_64_100), .A (n_61_99), .B (n_55_102), .C1 (n_51_104), .C2 (n_45_107) );
AOI211_X1 g_62_101 (.ZN (n_62_101), .A (n_63_98), .B (n_57_101), .C1 (n_53_103), .C2 (n_47_106) );
AOI211_X1 g_60_102 (.ZN (n_60_102), .A (n_64_100), .B (n_59_100), .C1 (n_55_102), .C2 (n_49_105) );
AOI211_X1 g_58_103 (.ZN (n_58_103), .A (n_62_101), .B (n_61_99), .C1 (n_57_101), .C2 (n_51_104) );
AOI211_X1 g_56_104 (.ZN (n_56_104), .A (n_60_102), .B (n_63_98), .C1 (n_59_100), .C2 (n_53_103) );
AOI211_X1 g_54_105 (.ZN (n_54_105), .A (n_58_103), .B (n_64_100), .C1 (n_61_99), .C2 (n_55_102) );
AOI211_X1 g_52_106 (.ZN (n_52_106), .A (n_56_104), .B (n_62_101), .C1 (n_63_98), .C2 (n_57_101) );
AOI211_X1 g_50_107 (.ZN (n_50_107), .A (n_54_105), .B (n_60_102), .C1 (n_64_100), .C2 (n_59_100) );
AOI211_X1 g_48_108 (.ZN (n_48_108), .A (n_52_106), .B (n_58_103), .C1 (n_62_101), .C2 (n_61_99) );
AOI211_X1 g_49_106 (.ZN (n_49_106), .A (n_50_107), .B (n_56_104), .C1 (n_60_102), .C2 (n_63_98) );
AOI211_X1 g_47_107 (.ZN (n_47_107), .A (n_48_108), .B (n_54_105), .C1 (n_58_103), .C2 (n_64_100) );
AOI211_X1 g_45_108 (.ZN (n_45_108), .A (n_49_106), .B (n_52_106), .C1 (n_56_104), .C2 (n_62_101) );
AOI211_X1 g_43_109 (.ZN (n_43_109), .A (n_47_107), .B (n_50_107), .C1 (n_54_105), .C2 (n_60_102) );
AOI211_X1 g_41_110 (.ZN (n_41_110), .A (n_45_108), .B (n_48_108), .C1 (n_52_106), .C2 (n_58_103) );
AOI211_X1 g_39_111 (.ZN (n_39_111), .A (n_43_109), .B (n_49_106), .C1 (n_50_107), .C2 (n_56_104) );
AOI211_X1 g_37_112 (.ZN (n_37_112), .A (n_41_110), .B (n_47_107), .C1 (n_48_108), .C2 (n_54_105) );
AOI211_X1 g_35_113 (.ZN (n_35_113), .A (n_39_111), .B (n_45_108), .C1 (n_49_106), .C2 (n_52_106) );
AOI211_X1 g_33_114 (.ZN (n_33_114), .A (n_37_112), .B (n_43_109), .C1 (n_47_107), .C2 (n_50_107) );
AOI211_X1 g_31_115 (.ZN (n_31_115), .A (n_35_113), .B (n_41_110), .C1 (n_45_108), .C2 (n_48_108) );
AOI211_X1 g_29_116 (.ZN (n_29_116), .A (n_33_114), .B (n_39_111), .C1 (n_43_109), .C2 (n_49_106) );
AOI211_X1 g_27_117 (.ZN (n_27_117), .A (n_31_115), .B (n_37_112), .C1 (n_41_110), .C2 (n_47_107) );
AOI211_X1 g_25_118 (.ZN (n_25_118), .A (n_29_116), .B (n_35_113), .C1 (n_39_111), .C2 (n_45_108) );
AOI211_X1 g_23_119 (.ZN (n_23_119), .A (n_27_117), .B (n_33_114), .C1 (n_37_112), .C2 (n_43_109) );
AOI211_X1 g_21_120 (.ZN (n_21_120), .A (n_25_118), .B (n_31_115), .C1 (n_35_113), .C2 (n_41_110) );
AOI211_X1 g_19_121 (.ZN (n_19_121), .A (n_23_119), .B (n_29_116), .C1 (n_33_114), .C2 (n_39_111) );
AOI211_X1 g_17_120 (.ZN (n_17_120), .A (n_21_120), .B (n_27_117), .C1 (n_31_115), .C2 (n_37_112) );
AOI211_X1 g_15_121 (.ZN (n_15_121), .A (n_19_121), .B (n_25_118), .C1 (n_29_116), .C2 (n_35_113) );
AOI211_X1 g_13_122 (.ZN (n_13_122), .A (n_17_120), .B (n_23_119), .C1 (n_27_117), .C2 (n_33_114) );
AOI211_X1 g_11_123 (.ZN (n_11_123), .A (n_15_121), .B (n_21_120), .C1 (n_25_118), .C2 (n_31_115) );
AOI211_X1 g_9_124 (.ZN (n_9_124), .A (n_13_122), .B (n_19_121), .C1 (n_23_119), .C2 (n_29_116) );
AOI211_X1 g_7_125 (.ZN (n_7_125), .A (n_11_123), .B (n_17_120), .C1 (n_21_120), .C2 (n_27_117) );
AOI211_X1 g_6_127 (.ZN (n_6_127), .A (n_9_124), .B (n_15_121), .C1 (n_19_121), .C2 (n_25_118) );
AOI211_X1 g_8_126 (.ZN (n_8_126), .A (n_7_125), .B (n_13_122), .C1 (n_17_120), .C2 (n_23_119) );
AOI211_X1 g_10_125 (.ZN (n_10_125), .A (n_6_127), .B (n_11_123), .C1 (n_15_121), .C2 (n_21_120) );
AOI211_X1 g_12_124 (.ZN (n_12_124), .A (n_8_126), .B (n_9_124), .C1 (n_13_122), .C2 (n_19_121) );
AOI211_X1 g_14_123 (.ZN (n_14_123), .A (n_10_125), .B (n_7_125), .C1 (n_11_123), .C2 (n_17_120) );
AOI211_X1 g_16_122 (.ZN (n_16_122), .A (n_12_124), .B (n_6_127), .C1 (n_9_124), .C2 (n_15_121) );
AOI211_X1 g_18_121 (.ZN (n_18_121), .A (n_14_123), .B (n_8_126), .C1 (n_7_125), .C2 (n_13_122) );
AOI211_X1 g_20_120 (.ZN (n_20_120), .A (n_16_122), .B (n_10_125), .C1 (n_6_127), .C2 (n_11_123) );
AOI211_X1 g_19_122 (.ZN (n_19_122), .A (n_18_121), .B (n_12_124), .C1 (n_8_126), .C2 (n_9_124) );
AOI211_X1 g_17_121 (.ZN (n_17_121), .A (n_20_120), .B (n_14_123), .C1 (n_10_125), .C2 (n_7_125) );
AOI211_X1 g_19_120 (.ZN (n_19_120), .A (n_19_122), .B (n_16_122), .C1 (n_12_124), .C2 (n_6_127) );
AOI211_X1 g_21_119 (.ZN (n_21_119), .A (n_17_121), .B (n_18_121), .C1 (n_14_123), .C2 (n_8_126) );
AOI211_X1 g_23_118 (.ZN (n_23_118), .A (n_19_120), .B (n_20_120), .C1 (n_16_122), .C2 (n_10_125) );
AOI211_X1 g_25_117 (.ZN (n_25_117), .A (n_21_119), .B (n_19_122), .C1 (n_18_121), .C2 (n_12_124) );
AOI211_X1 g_24_119 (.ZN (n_24_119), .A (n_23_118), .B (n_17_121), .C1 (n_20_120), .C2 (n_14_123) );
AOI211_X1 g_26_118 (.ZN (n_26_118), .A (n_25_117), .B (n_19_120), .C1 (n_19_122), .C2 (n_16_122) );
AOI211_X1 g_25_120 (.ZN (n_25_120), .A (n_24_119), .B (n_21_119), .C1 (n_17_121), .C2 (n_18_121) );
AOI211_X1 g_24_118 (.ZN (n_24_118), .A (n_26_118), .B (n_23_118), .C1 (n_19_120), .C2 (n_20_120) );
AOI211_X1 g_26_117 (.ZN (n_26_117), .A (n_25_120), .B (n_25_117), .C1 (n_21_119), .C2 (n_19_122) );
AOI211_X1 g_28_116 (.ZN (n_28_116), .A (n_24_118), .B (n_24_119), .C1 (n_23_118), .C2 (n_17_121) );
AOI211_X1 g_30_115 (.ZN (n_30_115), .A (n_26_117), .B (n_26_118), .C1 (n_25_117), .C2 (n_19_120) );
AOI211_X1 g_32_114 (.ZN (n_32_114), .A (n_28_116), .B (n_25_120), .C1 (n_24_119), .C2 (n_21_119) );
AOI211_X1 g_34_113 (.ZN (n_34_113), .A (n_30_115), .B (n_24_118), .C1 (n_26_118), .C2 (n_23_118) );
AOI211_X1 g_33_115 (.ZN (n_33_115), .A (n_32_114), .B (n_26_117), .C1 (n_25_120), .C2 (n_25_117) );
AOI211_X1 g_35_114 (.ZN (n_35_114), .A (n_34_113), .B (n_28_116), .C1 (n_24_118), .C2 (n_24_119) );
AOI211_X1 g_37_113 (.ZN (n_37_113), .A (n_33_115), .B (n_30_115), .C1 (n_26_117), .C2 (n_26_118) );
AOI211_X1 g_39_112 (.ZN (n_39_112), .A (n_35_114), .B (n_32_114), .C1 (n_28_116), .C2 (n_25_120) );
AOI211_X1 g_41_111 (.ZN (n_41_111), .A (n_37_113), .B (n_34_113), .C1 (n_30_115), .C2 (n_24_118) );
AOI211_X1 g_43_110 (.ZN (n_43_110), .A (n_39_112), .B (n_33_115), .C1 (n_32_114), .C2 (n_26_117) );
AOI211_X1 g_45_109 (.ZN (n_45_109), .A (n_41_111), .B (n_35_114), .C1 (n_34_113), .C2 (n_28_116) );
AOI211_X1 g_47_108 (.ZN (n_47_108), .A (n_43_110), .B (n_37_113), .C1 (n_33_115), .C2 (n_30_115) );
AOI211_X1 g_49_107 (.ZN (n_49_107), .A (n_45_109), .B (n_39_112), .C1 (n_35_114), .C2 (n_32_114) );
AOI211_X1 g_51_106 (.ZN (n_51_106), .A (n_47_108), .B (n_41_111), .C1 (n_37_113), .C2 (n_34_113) );
AOI211_X1 g_53_105 (.ZN (n_53_105), .A (n_49_107), .B (n_43_110), .C1 (n_39_112), .C2 (n_33_115) );
AOI211_X1 g_55_104 (.ZN (n_55_104), .A (n_51_106), .B (n_45_109), .C1 (n_41_111), .C2 (n_35_114) );
AOI211_X1 g_57_103 (.ZN (n_57_103), .A (n_53_105), .B (n_47_108), .C1 (n_43_110), .C2 (n_37_113) );
AOI211_X1 g_59_102 (.ZN (n_59_102), .A (n_55_104), .B (n_49_107), .C1 (n_45_109), .C2 (n_39_112) );
AOI211_X1 g_61_101 (.ZN (n_61_101), .A (n_57_103), .B (n_51_106), .C1 (n_47_108), .C2 (n_41_111) );
AOI211_X1 g_63_100 (.ZN (n_63_100), .A (n_59_102), .B (n_53_105), .C1 (n_49_107), .C2 (n_43_110) );
AOI211_X1 g_65_99 (.ZN (n_65_99), .A (n_61_101), .B (n_55_104), .C1 (n_51_106), .C2 (n_45_109) );
AOI211_X1 g_67_98 (.ZN (n_67_98), .A (n_63_100), .B (n_57_103), .C1 (n_53_105), .C2 (n_47_108) );
AOI211_X1 g_69_97 (.ZN (n_69_97), .A (n_65_99), .B (n_59_102), .C1 (n_55_104), .C2 (n_49_107) );
AOI211_X1 g_71_96 (.ZN (n_71_96), .A (n_67_98), .B (n_61_101), .C1 (n_57_103), .C2 (n_51_106) );
AOI211_X1 g_70_98 (.ZN (n_70_98), .A (n_69_97), .B (n_63_100), .C1 (n_59_102), .C2 (n_53_105) );
AOI211_X1 g_72_97 (.ZN (n_72_97), .A (n_71_96), .B (n_65_99), .C1 (n_61_101), .C2 (n_55_104) );
AOI211_X1 g_71_99 (.ZN (n_71_99), .A (n_70_98), .B (n_67_98), .C1 (n_63_100), .C2 (n_57_103) );
AOI211_X1 g_69_98 (.ZN (n_69_98), .A (n_72_97), .B (n_69_97), .C1 (n_65_99), .C2 (n_59_102) );
AOI211_X1 g_71_97 (.ZN (n_71_97), .A (n_71_99), .B (n_71_96), .C1 (n_67_98), .C2 (n_61_101) );
AOI211_X1 g_73_96 (.ZN (n_73_96), .A (n_69_98), .B (n_70_98), .C1 (n_69_97), .C2 (n_63_100) );
AOI211_X1 g_75_95 (.ZN (n_75_95), .A (n_71_97), .B (n_72_97), .C1 (n_71_96), .C2 (n_65_99) );
AOI211_X1 g_77_94 (.ZN (n_77_94), .A (n_73_96), .B (n_71_99), .C1 (n_70_98), .C2 (n_67_98) );
AOI211_X1 g_79_93 (.ZN (n_79_93), .A (n_75_95), .B (n_69_98), .C1 (n_72_97), .C2 (n_69_97) );
AOI211_X1 g_81_92 (.ZN (n_81_92), .A (n_77_94), .B (n_71_97), .C1 (n_71_99), .C2 (n_71_96) );
AOI211_X1 g_83_91 (.ZN (n_83_91), .A (n_79_93), .B (n_73_96), .C1 (n_69_98), .C2 (n_70_98) );
AOI211_X1 g_85_90 (.ZN (n_85_90), .A (n_81_92), .B (n_75_95), .C1 (n_71_97), .C2 (n_72_97) );
AOI211_X1 g_87_89 (.ZN (n_87_89), .A (n_83_91), .B (n_77_94), .C1 (n_73_96), .C2 (n_71_99) );
AOI211_X1 g_89_88 (.ZN (n_89_88), .A (n_85_90), .B (n_79_93), .C1 (n_75_95), .C2 (n_69_98) );
AOI211_X1 g_91_87 (.ZN (n_91_87), .A (n_87_89), .B (n_81_92), .C1 (n_77_94), .C2 (n_71_97) );
AOI211_X1 g_93_86 (.ZN (n_93_86), .A (n_89_88), .B (n_83_91), .C1 (n_79_93), .C2 (n_73_96) );
AOI211_X1 g_95_85 (.ZN (n_95_85), .A (n_91_87), .B (n_85_90), .C1 (n_81_92), .C2 (n_75_95) );
AOI211_X1 g_97_84 (.ZN (n_97_84), .A (n_93_86), .B (n_87_89), .C1 (n_83_91), .C2 (n_77_94) );
AOI211_X1 g_99_83 (.ZN (n_99_83), .A (n_95_85), .B (n_89_88), .C1 (n_85_90), .C2 (n_79_93) );
AOI211_X1 g_101_82 (.ZN (n_101_82), .A (n_97_84), .B (n_91_87), .C1 (n_87_89), .C2 (n_81_92) );
AOI211_X1 g_103_81 (.ZN (n_103_81), .A (n_99_83), .B (n_93_86), .C1 (n_89_88), .C2 (n_83_91) );
AOI211_X1 g_105_80 (.ZN (n_105_80), .A (n_101_82), .B (n_95_85), .C1 (n_91_87), .C2 (n_85_90) );
AOI211_X1 g_107_79 (.ZN (n_107_79), .A (n_103_81), .B (n_97_84), .C1 (n_93_86), .C2 (n_87_89) );
AOI211_X1 g_109_78 (.ZN (n_109_78), .A (n_105_80), .B (n_99_83), .C1 (n_95_85), .C2 (n_89_88) );
AOI211_X1 g_111_77 (.ZN (n_111_77), .A (n_107_79), .B (n_101_82), .C1 (n_97_84), .C2 (n_91_87) );
AOI211_X1 g_113_76 (.ZN (n_113_76), .A (n_109_78), .B (n_103_81), .C1 (n_99_83), .C2 (n_93_86) );
AOI211_X1 g_115_75 (.ZN (n_115_75), .A (n_111_77), .B (n_105_80), .C1 (n_101_82), .C2 (n_95_85) );
AOI211_X1 g_117_74 (.ZN (n_117_74), .A (n_113_76), .B (n_107_79), .C1 (n_103_81), .C2 (n_97_84) );
AOI211_X1 g_119_73 (.ZN (n_119_73), .A (n_115_75), .B (n_109_78), .C1 (n_105_80), .C2 (n_99_83) );
AOI211_X1 g_118_75 (.ZN (n_118_75), .A (n_117_74), .B (n_111_77), .C1 (n_107_79), .C2 (n_101_82) );
AOI211_X1 g_120_74 (.ZN (n_120_74), .A (n_119_73), .B (n_113_76), .C1 (n_109_78), .C2 (n_103_81) );
AOI211_X1 g_122_73 (.ZN (n_122_73), .A (n_118_75), .B (n_115_75), .C1 (n_111_77), .C2 (n_105_80) );
AOI211_X1 g_121_75 (.ZN (n_121_75), .A (n_120_74), .B (n_117_74), .C1 (n_113_76), .C2 (n_107_79) );
AOI211_X1 g_120_73 (.ZN (n_120_73), .A (n_122_73), .B (n_119_73), .C1 (n_115_75), .C2 (n_109_78) );
AOI211_X1 g_122_72 (.ZN (n_122_72), .A (n_121_75), .B (n_118_75), .C1 (n_117_74), .C2 (n_111_77) );
AOI211_X1 g_124_71 (.ZN (n_124_71), .A (n_120_73), .B (n_120_74), .C1 (n_119_73), .C2 (n_113_76) );
AOI211_X1 g_126_70 (.ZN (n_126_70), .A (n_122_72), .B (n_122_73), .C1 (n_118_75), .C2 (n_115_75) );
AOI211_X1 g_128_69 (.ZN (n_128_69), .A (n_124_71), .B (n_121_75), .C1 (n_120_74), .C2 (n_117_74) );
AOI211_X1 g_130_68 (.ZN (n_130_68), .A (n_126_70), .B (n_120_73), .C1 (n_122_73), .C2 (n_119_73) );
AOI211_X1 g_132_67 (.ZN (n_132_67), .A (n_128_69), .B (n_122_72), .C1 (n_121_75), .C2 (n_118_75) );
AOI211_X1 g_131_69 (.ZN (n_131_69), .A (n_130_68), .B (n_124_71), .C1 (n_120_73), .C2 (n_120_74) );
AOI211_X1 g_133_68 (.ZN (n_133_68), .A (n_132_67), .B (n_126_70), .C1 (n_122_72), .C2 (n_122_73) );
AOI211_X1 g_135_67 (.ZN (n_135_67), .A (n_131_69), .B (n_128_69), .C1 (n_124_71), .C2 (n_121_75) );
AOI211_X1 g_137_66 (.ZN (n_137_66), .A (n_133_68), .B (n_130_68), .C1 (n_126_70), .C2 (n_120_73) );
AOI211_X1 g_139_65 (.ZN (n_139_65), .A (n_135_67), .B (n_132_67), .C1 (n_128_69), .C2 (n_122_72) );
AOI211_X1 g_141_64 (.ZN (n_141_64), .A (n_137_66), .B (n_131_69), .C1 (n_130_68), .C2 (n_124_71) );
AOI211_X1 g_143_63 (.ZN (n_143_63), .A (n_139_65), .B (n_133_68), .C1 (n_132_67), .C2 (n_126_70) );
AOI211_X1 g_141_62 (.ZN (n_141_62), .A (n_141_64), .B (n_135_67), .C1 (n_131_69), .C2 (n_128_69) );
AOI211_X1 g_143_61 (.ZN (n_143_61), .A (n_143_63), .B (n_137_66), .C1 (n_133_68), .C2 (n_130_68) );
AOI211_X1 g_145_60 (.ZN (n_145_60), .A (n_141_62), .B (n_139_65), .C1 (n_135_67), .C2 (n_132_67) );
AOI211_X1 g_147_61 (.ZN (n_147_61), .A (n_143_61), .B (n_141_64), .C1 (n_137_66), .C2 (n_131_69) );
AOI211_X1 g_145_62 (.ZN (n_145_62), .A (n_145_60), .B (n_143_63), .C1 (n_139_65), .C2 (n_133_68) );
AOI211_X1 g_144_64 (.ZN (n_144_64), .A (n_147_61), .B (n_141_62), .C1 (n_141_64), .C2 (n_135_67) );
AOI211_X1 g_146_63 (.ZN (n_146_63), .A (n_145_62), .B (n_143_61), .C1 (n_143_63), .C2 (n_137_66) );
AOI211_X1 g_144_62 (.ZN (n_144_62), .A (n_144_64), .B (n_145_60), .C1 (n_141_62), .C2 (n_139_65) );
AOI211_X1 g_142_63 (.ZN (n_142_63), .A (n_146_63), .B (n_147_61), .C1 (n_143_61), .C2 (n_141_64) );
AOI211_X1 g_140_64 (.ZN (n_140_64), .A (n_144_62), .B (n_145_62), .C1 (n_145_60), .C2 (n_143_63) );
AOI211_X1 g_138_65 (.ZN (n_138_65), .A (n_142_63), .B (n_144_64), .C1 (n_147_61), .C2 (n_141_62) );
AOI211_X1 g_136_66 (.ZN (n_136_66), .A (n_140_64), .B (n_146_63), .C1 (n_145_62), .C2 (n_143_61) );
AOI211_X1 g_135_68 (.ZN (n_135_68), .A (n_138_65), .B (n_144_62), .C1 (n_144_64), .C2 (n_145_60) );
AOI211_X1 g_133_67 (.ZN (n_133_67), .A (n_136_66), .B (n_142_63), .C1 (n_146_63), .C2 (n_147_61) );
AOI211_X1 g_135_66 (.ZN (n_135_66), .A (n_135_68), .B (n_140_64), .C1 (n_144_62), .C2 (n_145_62) );
AOI211_X1 g_137_65 (.ZN (n_137_65), .A (n_133_67), .B (n_138_65), .C1 (n_142_63), .C2 (n_144_64) );
AOI211_X1 g_136_67 (.ZN (n_136_67), .A (n_135_66), .B (n_136_66), .C1 (n_140_64), .C2 (n_146_63) );
AOI211_X1 g_138_66 (.ZN (n_138_66), .A (n_137_65), .B (n_135_68), .C1 (n_138_65), .C2 (n_144_62) );
AOI211_X1 g_140_65 (.ZN (n_140_65), .A (n_136_67), .B (n_133_67), .C1 (n_136_66), .C2 (n_142_63) );
AOI211_X1 g_142_64 (.ZN (n_142_64), .A (n_138_66), .B (n_135_66), .C1 (n_135_68), .C2 (n_140_64) );
AOI211_X1 g_144_63 (.ZN (n_144_63), .A (n_140_65), .B (n_137_65), .C1 (n_133_67), .C2 (n_138_65) );
AOI211_X1 g_146_62 (.ZN (n_146_62), .A (n_142_64), .B (n_136_67), .C1 (n_135_66), .C2 (n_136_66) );
AOI211_X1 g_147_64 (.ZN (n_147_64), .A (n_144_63), .B (n_138_66), .C1 (n_137_65), .C2 (n_135_68) );
AOI211_X1 g_149_65 (.ZN (n_149_65), .A (n_146_62), .B (n_140_65), .C1 (n_136_67), .C2 (n_133_67) );
AOI211_X1 g_148_63 (.ZN (n_148_63), .A (n_147_64), .B (n_142_64), .C1 (n_138_66), .C2 (n_135_66) );
AOI211_X1 g_146_64 (.ZN (n_146_64), .A (n_149_65), .B (n_144_63), .C1 (n_140_65), .C2 (n_137_65) );
AOI211_X1 g_147_66 (.ZN (n_147_66), .A (n_148_63), .B (n_146_62), .C1 (n_142_64), .C2 (n_136_67) );
AOI211_X1 g_145_65 (.ZN (n_145_65), .A (n_146_64), .B (n_147_64), .C1 (n_144_63), .C2 (n_138_66) );
AOI211_X1 g_143_64 (.ZN (n_143_64), .A (n_147_66), .B (n_149_65), .C1 (n_146_62), .C2 (n_140_65) );
AOI211_X1 g_141_65 (.ZN (n_141_65), .A (n_145_65), .B (n_148_63), .C1 (n_147_64), .C2 (n_142_64) );
AOI211_X1 g_139_66 (.ZN (n_139_66), .A (n_143_64), .B (n_146_64), .C1 (n_149_65), .C2 (n_144_63) );
AOI211_X1 g_137_67 (.ZN (n_137_67), .A (n_141_65), .B (n_147_66), .C1 (n_148_63), .C2 (n_146_62) );
AOI211_X1 g_136_69 (.ZN (n_136_69), .A (n_139_66), .B (n_145_65), .C1 (n_146_64), .C2 (n_147_64) );
AOI211_X1 g_134_68 (.ZN (n_134_68), .A (n_137_67), .B (n_143_64), .C1 (n_147_66), .C2 (n_149_65) );
AOI211_X1 g_132_69 (.ZN (n_132_69), .A (n_136_69), .B (n_141_65), .C1 (n_145_65), .C2 (n_148_63) );
AOI211_X1 g_134_70 (.ZN (n_134_70), .A (n_134_68), .B (n_139_66), .C1 (n_143_64), .C2 (n_146_64) );
AOI211_X1 g_132_71 (.ZN (n_132_71), .A (n_132_69), .B (n_137_67), .C1 (n_141_65), .C2 (n_147_66) );
AOI211_X1 g_133_69 (.ZN (n_133_69), .A (n_134_70), .B (n_136_69), .C1 (n_139_66), .C2 (n_145_65) );
AOI211_X1 g_131_68 (.ZN (n_131_68), .A (n_132_71), .B (n_134_68), .C1 (n_137_67), .C2 (n_143_64) );
AOI211_X1 g_130_70 (.ZN (n_130_70), .A (n_133_69), .B (n_132_69), .C1 (n_136_69), .C2 (n_141_65) );
AOI211_X1 g_128_71 (.ZN (n_128_71), .A (n_131_68), .B (n_134_70), .C1 (n_134_68), .C2 (n_139_66) );
AOI211_X1 g_129_69 (.ZN (n_129_69), .A (n_130_70), .B (n_132_71), .C1 (n_132_69), .C2 (n_137_67) );
AOI211_X1 g_127_70 (.ZN (n_127_70), .A (n_128_71), .B (n_133_69), .C1 (n_134_70), .C2 (n_136_69) );
AOI211_X1 g_125_71 (.ZN (n_125_71), .A (n_129_69), .B (n_131_68), .C1 (n_132_71), .C2 (n_134_68) );
AOI211_X1 g_123_72 (.ZN (n_123_72), .A (n_127_70), .B (n_130_70), .C1 (n_133_69), .C2 (n_132_69) );
AOI211_X1 g_121_73 (.ZN (n_121_73), .A (n_125_71), .B (n_128_71), .C1 (n_131_68), .C2 (n_134_70) );
AOI211_X1 g_119_74 (.ZN (n_119_74), .A (n_123_72), .B (n_129_69), .C1 (n_130_70), .C2 (n_132_71) );
AOI211_X1 g_117_75 (.ZN (n_117_75), .A (n_121_73), .B (n_127_70), .C1 (n_128_71), .C2 (n_133_69) );
AOI211_X1 g_119_76 (.ZN (n_119_76), .A (n_119_74), .B (n_125_71), .C1 (n_129_69), .C2 (n_131_68) );
AOI211_X1 g_118_74 (.ZN (n_118_74), .A (n_117_75), .B (n_123_72), .C1 (n_127_70), .C2 (n_130_70) );
AOI211_X1 g_116_75 (.ZN (n_116_75), .A (n_119_76), .B (n_121_73), .C1 (n_125_71), .C2 (n_128_71) );
AOI211_X1 g_114_76 (.ZN (n_114_76), .A (n_118_74), .B (n_119_74), .C1 (n_123_72), .C2 (n_129_69) );
AOI211_X1 g_112_77 (.ZN (n_112_77), .A (n_116_75), .B (n_117_75), .C1 (n_121_73), .C2 (n_127_70) );
AOI211_X1 g_110_78 (.ZN (n_110_78), .A (n_114_76), .B (n_119_76), .C1 (n_119_74), .C2 (n_125_71) );
AOI211_X1 g_108_79 (.ZN (n_108_79), .A (n_112_77), .B (n_118_74), .C1 (n_117_75), .C2 (n_123_72) );
AOI211_X1 g_106_80 (.ZN (n_106_80), .A (n_110_78), .B (n_116_75), .C1 (n_119_76), .C2 (n_121_73) );
AOI211_X1 g_104_81 (.ZN (n_104_81), .A (n_108_79), .B (n_114_76), .C1 (n_118_74), .C2 (n_119_74) );
AOI211_X1 g_102_82 (.ZN (n_102_82), .A (n_106_80), .B (n_112_77), .C1 (n_116_75), .C2 (n_117_75) );
AOI211_X1 g_100_83 (.ZN (n_100_83), .A (n_104_81), .B (n_110_78), .C1 (n_114_76), .C2 (n_119_76) );
AOI211_X1 g_98_84 (.ZN (n_98_84), .A (n_102_82), .B (n_108_79), .C1 (n_112_77), .C2 (n_118_74) );
AOI211_X1 g_97_86 (.ZN (n_97_86), .A (n_100_83), .B (n_106_80), .C1 (n_110_78), .C2 (n_116_75) );
AOI211_X1 g_99_85 (.ZN (n_99_85), .A (n_98_84), .B (n_104_81), .C1 (n_108_79), .C2 (n_114_76) );
AOI211_X1 g_101_84 (.ZN (n_101_84), .A (n_97_86), .B (n_102_82), .C1 (n_106_80), .C2 (n_112_77) );
AOI211_X1 g_103_83 (.ZN (n_103_83), .A (n_99_85), .B (n_100_83), .C1 (n_104_81), .C2 (n_110_78) );
AOI211_X1 g_105_82 (.ZN (n_105_82), .A (n_101_84), .B (n_98_84), .C1 (n_102_82), .C2 (n_108_79) );
AOI211_X1 g_107_81 (.ZN (n_107_81), .A (n_103_83), .B (n_97_86), .C1 (n_100_83), .C2 (n_106_80) );
AOI211_X1 g_109_80 (.ZN (n_109_80), .A (n_105_82), .B (n_99_85), .C1 (n_98_84), .C2 (n_104_81) );
AOI211_X1 g_111_79 (.ZN (n_111_79), .A (n_107_81), .B (n_101_84), .C1 (n_97_86), .C2 (n_102_82) );
AOI211_X1 g_113_78 (.ZN (n_113_78), .A (n_109_80), .B (n_103_83), .C1 (n_99_85), .C2 (n_100_83) );
AOI211_X1 g_115_77 (.ZN (n_115_77), .A (n_111_79), .B (n_105_82), .C1 (n_101_84), .C2 (n_98_84) );
AOI211_X1 g_117_76 (.ZN (n_117_76), .A (n_113_78), .B (n_107_81), .C1 (n_103_83), .C2 (n_97_86) );
AOI211_X1 g_119_75 (.ZN (n_119_75), .A (n_115_77), .B (n_109_80), .C1 (n_105_82), .C2 (n_99_85) );
AOI211_X1 g_121_74 (.ZN (n_121_74), .A (n_117_76), .B (n_111_79), .C1 (n_107_81), .C2 (n_101_84) );
AOI211_X1 g_123_73 (.ZN (n_123_73), .A (n_119_75), .B (n_113_78), .C1 (n_109_80), .C2 (n_103_83) );
AOI211_X1 g_125_72 (.ZN (n_125_72), .A (n_121_74), .B (n_115_77), .C1 (n_111_79), .C2 (n_105_82) );
AOI211_X1 g_127_71 (.ZN (n_127_71), .A (n_123_73), .B (n_117_76), .C1 (n_113_78), .C2 (n_107_81) );
AOI211_X1 g_129_70 (.ZN (n_129_70), .A (n_125_72), .B (n_119_75), .C1 (n_115_77), .C2 (n_109_80) );
AOI211_X1 g_128_72 (.ZN (n_128_72), .A (n_127_71), .B (n_121_74), .C1 (n_117_76), .C2 (n_111_79) );
AOI211_X1 g_130_71 (.ZN (n_130_71), .A (n_129_70), .B (n_123_73), .C1 (n_119_75), .C2 (n_113_78) );
AOI211_X1 g_132_70 (.ZN (n_132_70), .A (n_128_72), .B (n_125_72), .C1 (n_121_74), .C2 (n_115_77) );
AOI211_X1 g_134_69 (.ZN (n_134_69), .A (n_130_71), .B (n_127_71), .C1 (n_123_73), .C2 (n_117_76) );
AOI211_X1 g_136_68 (.ZN (n_136_68), .A (n_132_70), .B (n_129_70), .C1 (n_125_72), .C2 (n_119_75) );
AOI211_X1 g_138_67 (.ZN (n_138_67), .A (n_134_69), .B (n_128_72), .C1 (n_127_71), .C2 (n_121_74) );
AOI211_X1 g_140_66 (.ZN (n_140_66), .A (n_136_68), .B (n_130_71), .C1 (n_129_70), .C2 (n_123_73) );
AOI211_X1 g_142_65 (.ZN (n_142_65), .A (n_138_67), .B (n_132_70), .C1 (n_128_72), .C2 (n_125_72) );
AOI211_X1 g_141_67 (.ZN (n_141_67), .A (n_140_66), .B (n_134_69), .C1 (n_130_71), .C2 (n_127_71) );
AOI211_X1 g_143_66 (.ZN (n_143_66), .A (n_142_65), .B (n_136_68), .C1 (n_132_70), .C2 (n_129_70) );
AOI211_X1 g_145_67 (.ZN (n_145_67), .A (n_141_67), .B (n_138_67), .C1 (n_134_69), .C2 (n_128_72) );
AOI211_X1 g_144_65 (.ZN (n_144_65), .A (n_143_66), .B (n_140_66), .C1 (n_136_68), .C2 (n_130_71) );
AOI211_X1 g_142_66 (.ZN (n_142_66), .A (n_145_67), .B (n_142_65), .C1 (n_138_67), .C2 (n_132_70) );
AOI211_X1 g_140_67 (.ZN (n_140_67), .A (n_144_65), .B (n_141_67), .C1 (n_140_66), .C2 (n_134_69) );
AOI211_X1 g_138_68 (.ZN (n_138_68), .A (n_142_66), .B (n_143_66), .C1 (n_142_65), .C2 (n_136_68) );
AOI211_X1 g_137_70 (.ZN (n_137_70), .A (n_140_67), .B (n_145_67), .C1 (n_141_67), .C2 (n_138_67) );
AOI211_X1 g_135_69 (.ZN (n_135_69), .A (n_138_68), .B (n_144_65), .C1 (n_143_66), .C2 (n_140_66) );
AOI211_X1 g_137_68 (.ZN (n_137_68), .A (n_137_70), .B (n_142_66), .C1 (n_145_67), .C2 (n_142_65) );
AOI211_X1 g_139_67 (.ZN (n_139_67), .A (n_135_69), .B (n_140_67), .C1 (n_144_65), .C2 (n_141_67) );
AOI211_X1 g_141_66 (.ZN (n_141_66), .A (n_137_68), .B (n_138_68), .C1 (n_142_66), .C2 (n_143_66) );
AOI211_X1 g_143_65 (.ZN (n_143_65), .A (n_139_67), .B (n_137_70), .C1 (n_140_67), .C2 (n_145_67) );
AOI211_X1 g_145_64 (.ZN (n_145_64), .A (n_141_66), .B (n_135_69), .C1 (n_138_68), .C2 (n_144_65) );
AOI211_X1 g_147_65 (.ZN (n_147_65), .A (n_143_65), .B (n_137_68), .C1 (n_137_70), .C2 (n_142_66) );
AOI211_X1 g_145_66 (.ZN (n_145_66), .A (n_145_64), .B (n_139_67), .C1 (n_135_69), .C2 (n_140_67) );
AOI211_X1 g_143_67 (.ZN (n_143_67), .A (n_147_65), .B (n_141_66), .C1 (n_137_68), .C2 (n_138_68) );
AOI211_X1 g_141_68 (.ZN (n_141_68), .A (n_145_66), .B (n_143_65), .C1 (n_139_67), .C2 (n_137_70) );
AOI211_X1 g_139_69 (.ZN (n_139_69), .A (n_143_67), .B (n_145_64), .C1 (n_141_66), .C2 (n_135_69) );
AOI211_X1 g_138_71 (.ZN (n_138_71), .A (n_141_68), .B (n_147_65), .C1 (n_143_65), .C2 (n_137_68) );
AOI211_X1 g_137_69 (.ZN (n_137_69), .A (n_139_69), .B (n_145_66), .C1 (n_145_64), .C2 (n_139_67) );
AOI211_X1 g_139_68 (.ZN (n_139_68), .A (n_138_71), .B (n_143_67), .C1 (n_147_65), .C2 (n_141_66) );
AOI211_X1 g_138_70 (.ZN (n_138_70), .A (n_137_69), .B (n_141_68), .C1 (n_145_66), .C2 (n_143_65) );
AOI211_X1 g_140_69 (.ZN (n_140_69), .A (n_139_68), .B (n_139_69), .C1 (n_143_67), .C2 (n_145_64) );
AOI211_X1 g_142_68 (.ZN (n_142_68), .A (n_138_70), .B (n_138_71), .C1 (n_141_68), .C2 (n_147_65) );
AOI211_X1 g_144_67 (.ZN (n_144_67), .A (n_140_69), .B (n_137_69), .C1 (n_139_69), .C2 (n_145_66) );
AOI211_X1 g_146_66 (.ZN (n_146_66), .A (n_142_68), .B (n_139_68), .C1 (n_138_71), .C2 (n_143_67) );
AOI211_X1 g_147_68 (.ZN (n_147_68), .A (n_144_67), .B (n_138_70), .C1 (n_137_69), .C2 (n_141_68) );
AOI211_X1 g_149_69 (.ZN (n_149_69), .A (n_146_66), .B (n_140_69), .C1 (n_139_68), .C2 (n_139_69) );
AOI211_X1 g_148_67 (.ZN (n_148_67), .A (n_147_68), .B (n_142_68), .C1 (n_138_70), .C2 (n_138_71) );
AOI211_X1 g_146_68 (.ZN (n_146_68), .A (n_149_69), .B (n_144_67), .C1 (n_140_69), .C2 (n_137_69) );
AOI211_X1 g_147_70 (.ZN (n_147_70), .A (n_148_67), .B (n_146_66), .C1 (n_142_68), .C2 (n_139_68) );
AOI211_X1 g_145_69 (.ZN (n_145_69), .A (n_146_68), .B (n_147_68), .C1 (n_144_67), .C2 (n_138_70) );
AOI211_X1 g_146_67 (.ZN (n_146_67), .A (n_147_70), .B (n_149_69), .C1 (n_146_66), .C2 (n_140_69) );
AOI211_X1 g_144_66 (.ZN (n_144_66), .A (n_145_69), .B (n_148_67), .C1 (n_147_68), .C2 (n_142_68) );
AOI211_X1 g_143_68 (.ZN (n_143_68), .A (n_146_67), .B (n_146_68), .C1 (n_149_69), .C2 (n_144_67) );
AOI211_X1 g_141_69 (.ZN (n_141_69), .A (n_144_66), .B (n_147_70), .C1 (n_148_67), .C2 (n_146_66) );
AOI211_X1 g_142_67 (.ZN (n_142_67), .A (n_143_68), .B (n_145_69), .C1 (n_146_68), .C2 (n_147_68) );
AOI211_X1 g_144_68 (.ZN (n_144_68), .A (n_141_69), .B (n_146_67), .C1 (n_147_70), .C2 (n_149_69) );
AOI211_X1 g_143_70 (.ZN (n_143_70), .A (n_142_67), .B (n_144_66), .C1 (n_145_69), .C2 (n_148_67) );
AOI211_X1 g_145_71 (.ZN (n_145_71), .A (n_144_68), .B (n_143_68), .C1 (n_146_67), .C2 (n_146_68) );
AOI211_X1 g_144_69 (.ZN (n_144_69), .A (n_143_70), .B (n_141_69), .C1 (n_144_66), .C2 (n_147_70) );
AOI211_X1 g_142_70 (.ZN (n_142_70), .A (n_145_71), .B (n_142_67), .C1 (n_143_68), .C2 (n_145_69) );
AOI211_X1 g_140_71 (.ZN (n_140_71), .A (n_144_69), .B (n_144_68), .C1 (n_141_69), .C2 (n_146_67) );
AOI211_X1 g_138_72 (.ZN (n_138_72), .A (n_142_70), .B (n_143_70), .C1 (n_142_67), .C2 (n_144_66) );
AOI211_X1 g_136_71 (.ZN (n_136_71), .A (n_140_71), .B (n_145_71), .C1 (n_144_68), .C2 (n_143_68) );
AOI211_X1 g_134_72 (.ZN (n_134_72), .A (n_138_72), .B (n_144_69), .C1 (n_143_70), .C2 (n_141_69) );
AOI211_X1 g_135_70 (.ZN (n_135_70), .A (n_136_71), .B (n_142_70), .C1 (n_145_71), .C2 (n_142_67) );
AOI211_X1 g_133_71 (.ZN (n_133_71), .A (n_134_72), .B (n_140_71), .C1 (n_144_69), .C2 (n_144_68) );
AOI211_X1 g_131_70 (.ZN (n_131_70), .A (n_135_70), .B (n_138_72), .C1 (n_142_70), .C2 (n_143_70) );
AOI211_X1 g_129_71 (.ZN (n_129_71), .A (n_133_71), .B (n_136_71), .C1 (n_140_71), .C2 (n_145_71) );
AOI211_X1 g_127_72 (.ZN (n_127_72), .A (n_131_70), .B (n_134_72), .C1 (n_138_72), .C2 (n_144_69) );
AOI211_X1 g_125_73 (.ZN (n_125_73), .A (n_129_71), .B (n_135_70), .C1 (n_136_71), .C2 (n_142_70) );
AOI211_X1 g_123_74 (.ZN (n_123_74), .A (n_127_72), .B (n_133_71), .C1 (n_134_72), .C2 (n_140_71) );
AOI211_X1 g_122_76 (.ZN (n_122_76), .A (n_125_73), .B (n_131_70), .C1 (n_135_70), .C2 (n_138_72) );
AOI211_X1 g_120_75 (.ZN (n_120_75), .A (n_123_74), .B (n_129_71), .C1 (n_133_71), .C2 (n_136_71) );
AOI211_X1 g_122_74 (.ZN (n_122_74), .A (n_122_76), .B (n_127_72), .C1 (n_131_70), .C2 (n_134_72) );
AOI211_X1 g_124_73 (.ZN (n_124_73), .A (n_120_75), .B (n_125_73), .C1 (n_129_71), .C2 (n_135_70) );
AOI211_X1 g_126_72 (.ZN (n_126_72), .A (n_122_74), .B (n_123_74), .C1 (n_127_72), .C2 (n_133_71) );
AOI211_X1 g_125_74 (.ZN (n_125_74), .A (n_124_73), .B (n_122_76), .C1 (n_125_73), .C2 (n_131_70) );
AOI211_X1 g_127_73 (.ZN (n_127_73), .A (n_126_72), .B (n_120_75), .C1 (n_123_74), .C2 (n_129_71) );
AOI211_X1 g_129_72 (.ZN (n_129_72), .A (n_125_74), .B (n_122_74), .C1 (n_122_76), .C2 (n_127_72) );
AOI211_X1 g_131_71 (.ZN (n_131_71), .A (n_127_73), .B (n_124_73), .C1 (n_120_75), .C2 (n_125_73) );
AOI211_X1 g_133_70 (.ZN (n_133_70), .A (n_129_72), .B (n_126_72), .C1 (n_122_74), .C2 (n_123_74) );
AOI211_X1 g_135_71 (.ZN (n_135_71), .A (n_131_71), .B (n_125_74), .C1 (n_124_73), .C2 (n_122_76) );
AOI211_X1 g_133_72 (.ZN (n_133_72), .A (n_133_70), .B (n_127_73), .C1 (n_126_72), .C2 (n_120_75) );
AOI211_X1 g_131_73 (.ZN (n_131_73), .A (n_135_71), .B (n_129_72), .C1 (n_125_74), .C2 (n_122_74) );
AOI211_X1 g_129_74 (.ZN (n_129_74), .A (n_133_72), .B (n_131_71), .C1 (n_127_73), .C2 (n_124_73) );
AOI211_X1 g_130_72 (.ZN (n_130_72), .A (n_131_73), .B (n_133_70), .C1 (n_129_72), .C2 (n_126_72) );
AOI211_X1 g_128_73 (.ZN (n_128_73), .A (n_129_74), .B (n_135_71), .C1 (n_131_71), .C2 (n_125_74) );
AOI211_X1 g_126_74 (.ZN (n_126_74), .A (n_130_72), .B (n_133_72), .C1 (n_133_70), .C2 (n_127_73) );
AOI211_X1 g_124_75 (.ZN (n_124_75), .A (n_128_73), .B (n_131_73), .C1 (n_135_71), .C2 (n_129_72) );
AOI211_X1 g_126_76 (.ZN (n_126_76), .A (n_126_74), .B (n_129_74), .C1 (n_133_72), .C2 (n_131_71) );
AOI211_X1 g_127_74 (.ZN (n_127_74), .A (n_124_75), .B (n_130_72), .C1 (n_131_73), .C2 (n_133_70) );
AOI211_X1 g_129_73 (.ZN (n_129_73), .A (n_126_76), .B (n_128_73), .C1 (n_129_74), .C2 (n_135_71) );
AOI211_X1 g_131_72 (.ZN (n_131_72), .A (n_127_74), .B (n_126_74), .C1 (n_130_72), .C2 (n_133_72) );
AOI211_X1 g_130_74 (.ZN (n_130_74), .A (n_129_73), .B (n_124_75), .C1 (n_128_73), .C2 (n_131_73) );
AOI211_X1 g_132_73 (.ZN (n_132_73), .A (n_131_72), .B (n_126_76), .C1 (n_126_74), .C2 (n_129_74) );
AOI211_X1 g_131_75 (.ZN (n_131_75), .A (n_130_74), .B (n_127_74), .C1 (n_124_75), .C2 (n_130_72) );
AOI211_X1 g_130_73 (.ZN (n_130_73), .A (n_132_73), .B (n_129_73), .C1 (n_126_76), .C2 (n_128_73) );
AOI211_X1 g_132_72 (.ZN (n_132_72), .A (n_131_75), .B (n_131_72), .C1 (n_127_74), .C2 (n_126_74) );
AOI211_X1 g_134_71 (.ZN (n_134_71), .A (n_130_73), .B (n_130_74), .C1 (n_129_73), .C2 (n_124_75) );
AOI211_X1 g_136_70 (.ZN (n_136_70), .A (n_132_72), .B (n_132_73), .C1 (n_131_72), .C2 (n_126_76) );
AOI211_X1 g_138_69 (.ZN (n_138_69), .A (n_134_71), .B (n_131_75), .C1 (n_130_74), .C2 (n_127_74) );
AOI211_X1 g_140_68 (.ZN (n_140_68), .A (n_136_70), .B (n_130_73), .C1 (n_132_73), .C2 (n_129_73) );
AOI211_X1 g_139_70 (.ZN (n_139_70), .A (n_138_69), .B (n_132_72), .C1 (n_131_75), .C2 (n_131_72) );
AOI211_X1 g_137_71 (.ZN (n_137_71), .A (n_140_68), .B (n_134_71), .C1 (n_130_73), .C2 (n_130_74) );
AOI211_X1 g_135_72 (.ZN (n_135_72), .A (n_139_70), .B (n_136_70), .C1 (n_132_72), .C2 (n_132_73) );
AOI211_X1 g_133_73 (.ZN (n_133_73), .A (n_137_71), .B (n_138_69), .C1 (n_134_71), .C2 (n_131_75) );
AOI211_X1 g_131_74 (.ZN (n_131_74), .A (n_135_72), .B (n_140_68), .C1 (n_136_70), .C2 (n_130_73) );
AOI211_X1 g_129_75 (.ZN (n_129_75), .A (n_133_73), .B (n_139_70), .C1 (n_138_69), .C2 (n_132_72) );
AOI211_X1 g_127_76 (.ZN (n_127_76), .A (n_131_74), .B (n_137_71), .C1 (n_140_68), .C2 (n_134_71) );
AOI211_X1 g_128_74 (.ZN (n_128_74), .A (n_129_75), .B (n_135_72), .C1 (n_139_70), .C2 (n_136_70) );
AOI211_X1 g_126_73 (.ZN (n_126_73), .A (n_127_76), .B (n_133_73), .C1 (n_137_71), .C2 (n_138_69) );
AOI211_X1 g_125_75 (.ZN (n_125_75), .A (n_128_74), .B (n_131_74), .C1 (n_135_72), .C2 (n_140_68) );
AOI211_X1 g_123_76 (.ZN (n_123_76), .A (n_126_73), .B (n_129_75), .C1 (n_133_73), .C2 (n_139_70) );
AOI211_X1 g_124_74 (.ZN (n_124_74), .A (n_125_75), .B (n_127_76), .C1 (n_131_74), .C2 (n_137_71) );
AOI211_X1 g_122_75 (.ZN (n_122_75), .A (n_123_76), .B (n_128_74), .C1 (n_129_75), .C2 (n_135_72) );
AOI211_X1 g_120_76 (.ZN (n_120_76), .A (n_124_74), .B (n_126_73), .C1 (n_127_76), .C2 (n_133_73) );
AOI211_X1 g_118_77 (.ZN (n_118_77), .A (n_122_75), .B (n_125_75), .C1 (n_128_74), .C2 (n_131_74) );
AOI211_X1 g_116_76 (.ZN (n_116_76), .A (n_120_76), .B (n_123_76), .C1 (n_126_73), .C2 (n_129_75) );
AOI211_X1 g_114_77 (.ZN (n_114_77), .A (n_118_77), .B (n_124_74), .C1 (n_125_75), .C2 (n_127_76) );
AOI211_X1 g_112_78 (.ZN (n_112_78), .A (n_116_76), .B (n_122_75), .C1 (n_123_76), .C2 (n_128_74) );
AOI211_X1 g_110_79 (.ZN (n_110_79), .A (n_114_77), .B (n_120_76), .C1 (n_124_74), .C2 (n_126_73) );
AOI211_X1 g_108_80 (.ZN (n_108_80), .A (n_112_78), .B (n_118_77), .C1 (n_122_75), .C2 (n_125_75) );
AOI211_X1 g_106_81 (.ZN (n_106_81), .A (n_110_79), .B (n_116_76), .C1 (n_120_76), .C2 (n_123_76) );
AOI211_X1 g_104_82 (.ZN (n_104_82), .A (n_108_80), .B (n_114_77), .C1 (n_118_77), .C2 (n_124_74) );
AOI211_X1 g_102_83 (.ZN (n_102_83), .A (n_106_81), .B (n_112_78), .C1 (n_116_76), .C2 (n_122_75) );
AOI211_X1 g_100_84 (.ZN (n_100_84), .A (n_104_82), .B (n_110_79), .C1 (n_114_77), .C2 (n_120_76) );
AOI211_X1 g_98_85 (.ZN (n_98_85), .A (n_102_83), .B (n_108_80), .C1 (n_112_78), .C2 (n_118_77) );
AOI211_X1 g_96_86 (.ZN (n_96_86), .A (n_100_84), .B (n_106_81), .C1 (n_110_79), .C2 (n_116_76) );
AOI211_X1 g_94_87 (.ZN (n_94_87), .A (n_98_85), .B (n_104_82), .C1 (n_108_80), .C2 (n_114_77) );
AOI211_X1 g_92_88 (.ZN (n_92_88), .A (n_96_86), .B (n_102_83), .C1 (n_106_81), .C2 (n_112_78) );
AOI211_X1 g_90_89 (.ZN (n_90_89), .A (n_94_87), .B (n_100_84), .C1 (n_104_82), .C2 (n_110_79) );
AOI211_X1 g_88_90 (.ZN (n_88_90), .A (n_92_88), .B (n_98_85), .C1 (n_102_83), .C2 (n_108_80) );
AOI211_X1 g_86_91 (.ZN (n_86_91), .A (n_90_89), .B (n_96_86), .C1 (n_100_84), .C2 (n_106_81) );
AOI211_X1 g_84_92 (.ZN (n_84_92), .A (n_88_90), .B (n_94_87), .C1 (n_98_85), .C2 (n_104_82) );
AOI211_X1 g_82_93 (.ZN (n_82_93), .A (n_86_91), .B (n_92_88), .C1 (n_96_86), .C2 (n_102_83) );
AOI211_X1 g_80_94 (.ZN (n_80_94), .A (n_84_92), .B (n_90_89), .C1 (n_94_87), .C2 (n_100_84) );
AOI211_X1 g_78_95 (.ZN (n_78_95), .A (n_82_93), .B (n_88_90), .C1 (n_92_88), .C2 (n_98_85) );
AOI211_X1 g_76_96 (.ZN (n_76_96), .A (n_80_94), .B (n_86_91), .C1 (n_90_89), .C2 (n_96_86) );
AOI211_X1 g_74_97 (.ZN (n_74_97), .A (n_78_95), .B (n_84_92), .C1 (n_88_90), .C2 (n_94_87) );
AOI211_X1 g_72_98 (.ZN (n_72_98), .A (n_76_96), .B (n_82_93), .C1 (n_86_91), .C2 (n_92_88) );
AOI211_X1 g_70_99 (.ZN (n_70_99), .A (n_74_97), .B (n_80_94), .C1 (n_84_92), .C2 (n_90_89) );
AOI211_X1 g_68_98 (.ZN (n_68_98), .A (n_72_98), .B (n_78_95), .C1 (n_82_93), .C2 (n_88_90) );
AOI211_X1 g_67_100 (.ZN (n_67_100), .A (n_70_99), .B (n_76_96), .C1 (n_80_94), .C2 (n_86_91) );
AOI211_X1 g_69_99 (.ZN (n_69_99), .A (n_68_98), .B (n_74_97), .C1 (n_78_95), .C2 (n_84_92) );
AOI211_X1 g_71_98 (.ZN (n_71_98), .A (n_67_100), .B (n_72_98), .C1 (n_76_96), .C2 (n_82_93) );
AOI211_X1 g_73_97 (.ZN (n_73_97), .A (n_69_99), .B (n_70_99), .C1 (n_74_97), .C2 (n_80_94) );
AOI211_X1 g_75_96 (.ZN (n_75_96), .A (n_71_98), .B (n_68_98), .C1 (n_72_98), .C2 (n_78_95) );
AOI211_X1 g_77_95 (.ZN (n_77_95), .A (n_73_97), .B (n_67_100), .C1 (n_70_99), .C2 (n_76_96) );
AOI211_X1 g_76_97 (.ZN (n_76_97), .A (n_75_96), .B (n_69_99), .C1 (n_68_98), .C2 (n_74_97) );
AOI211_X1 g_74_98 (.ZN (n_74_98), .A (n_77_95), .B (n_71_98), .C1 (n_67_100), .C2 (n_72_98) );
AOI211_X1 g_72_99 (.ZN (n_72_99), .A (n_76_97), .B (n_73_97), .C1 (n_69_99), .C2 (n_70_99) );
AOI211_X1 g_70_100 (.ZN (n_70_100), .A (n_74_98), .B (n_75_96), .C1 (n_71_98), .C2 (n_68_98) );
AOI211_X1 g_68_99 (.ZN (n_68_99), .A (n_72_99), .B (n_77_95), .C1 (n_73_97), .C2 (n_67_100) );
AOI211_X1 g_66_100 (.ZN (n_66_100), .A (n_70_100), .B (n_76_97), .C1 (n_75_96), .C2 (n_69_99) );
AOI211_X1 g_64_99 (.ZN (n_64_99), .A (n_68_99), .B (n_74_98), .C1 (n_77_95), .C2 (n_71_98) );
AOI211_X1 g_62_100 (.ZN (n_62_100), .A (n_66_100), .B (n_72_99), .C1 (n_76_97), .C2 (n_73_97) );
AOI211_X1 g_60_101 (.ZN (n_60_101), .A (n_64_99), .B (n_70_100), .C1 (n_74_98), .C2 (n_75_96) );
AOI211_X1 g_58_102 (.ZN (n_58_102), .A (n_62_100), .B (n_68_99), .C1 (n_72_99), .C2 (n_77_95) );
AOI211_X1 g_56_103 (.ZN (n_56_103), .A (n_60_101), .B (n_66_100), .C1 (n_70_100), .C2 (n_76_97) );
AOI211_X1 g_54_104 (.ZN (n_54_104), .A (n_58_102), .B (n_64_99), .C1 (n_68_99), .C2 (n_74_98) );
AOI211_X1 g_52_105 (.ZN (n_52_105), .A (n_56_103), .B (n_62_100), .C1 (n_66_100), .C2 (n_72_99) );
AOI211_X1 g_50_106 (.ZN (n_50_106), .A (n_54_104), .B (n_60_101), .C1 (n_64_99), .C2 (n_70_100) );
AOI211_X1 g_48_107 (.ZN (n_48_107), .A (n_52_105), .B (n_58_102), .C1 (n_62_100), .C2 (n_68_99) );
AOI211_X1 g_46_108 (.ZN (n_46_108), .A (n_50_106), .B (n_56_103), .C1 (n_60_101), .C2 (n_66_100) );
AOI211_X1 g_44_109 (.ZN (n_44_109), .A (n_48_107), .B (n_54_104), .C1 (n_58_102), .C2 (n_64_99) );
AOI211_X1 g_42_110 (.ZN (n_42_110), .A (n_46_108), .B (n_52_105), .C1 (n_56_103), .C2 (n_62_100) );
AOI211_X1 g_40_111 (.ZN (n_40_111), .A (n_44_109), .B (n_50_106), .C1 (n_54_104), .C2 (n_60_101) );
AOI211_X1 g_38_112 (.ZN (n_38_112), .A (n_42_110), .B (n_48_107), .C1 (n_52_105), .C2 (n_58_102) );
AOI211_X1 g_36_113 (.ZN (n_36_113), .A (n_40_111), .B (n_46_108), .C1 (n_50_106), .C2 (n_56_103) );
AOI211_X1 g_34_114 (.ZN (n_34_114), .A (n_38_112), .B (n_44_109), .C1 (n_48_107), .C2 (n_54_104) );
AOI211_X1 g_33_116 (.ZN (n_33_116), .A (n_36_113), .B (n_42_110), .C1 (n_46_108), .C2 (n_52_105) );
AOI211_X1 g_35_115 (.ZN (n_35_115), .A (n_34_114), .B (n_40_111), .C1 (n_44_109), .C2 (n_50_106) );
AOI211_X1 g_37_114 (.ZN (n_37_114), .A (n_33_116), .B (n_38_112), .C1 (n_42_110), .C2 (n_48_107) );
AOI211_X1 g_39_113 (.ZN (n_39_113), .A (n_35_115), .B (n_36_113), .C1 (n_40_111), .C2 (n_46_108) );
AOI211_X1 g_41_112 (.ZN (n_41_112), .A (n_37_114), .B (n_34_114), .C1 (n_38_112), .C2 (n_44_109) );
AOI211_X1 g_43_111 (.ZN (n_43_111), .A (n_39_113), .B (n_33_116), .C1 (n_36_113), .C2 (n_42_110) );
AOI211_X1 g_45_110 (.ZN (n_45_110), .A (n_41_112), .B (n_35_115), .C1 (n_34_114), .C2 (n_40_111) );
AOI211_X1 g_47_109 (.ZN (n_47_109), .A (n_43_111), .B (n_37_114), .C1 (n_33_116), .C2 (n_38_112) );
AOI211_X1 g_49_108 (.ZN (n_49_108), .A (n_45_110), .B (n_39_113), .C1 (n_35_115), .C2 (n_36_113) );
AOI211_X1 g_51_107 (.ZN (n_51_107), .A (n_47_109), .B (n_41_112), .C1 (n_37_114), .C2 (n_34_114) );
AOI211_X1 g_53_106 (.ZN (n_53_106), .A (n_49_108), .B (n_43_111), .C1 (n_39_113), .C2 (n_33_116) );
AOI211_X1 g_55_105 (.ZN (n_55_105), .A (n_51_107), .B (n_45_110), .C1 (n_41_112), .C2 (n_35_115) );
AOI211_X1 g_57_104 (.ZN (n_57_104), .A (n_53_106), .B (n_47_109), .C1 (n_43_111), .C2 (n_37_114) );
AOI211_X1 g_59_103 (.ZN (n_59_103), .A (n_55_105), .B (n_49_108), .C1 (n_45_110), .C2 (n_39_113) );
AOI211_X1 g_61_102 (.ZN (n_61_102), .A (n_57_104), .B (n_51_107), .C1 (n_47_109), .C2 (n_41_112) );
AOI211_X1 g_63_101 (.ZN (n_63_101), .A (n_59_103), .B (n_53_106), .C1 (n_49_108), .C2 (n_43_111) );
AOI211_X1 g_65_100 (.ZN (n_65_100), .A (n_61_102), .B (n_55_105), .C1 (n_51_107), .C2 (n_45_110) );
AOI211_X1 g_67_99 (.ZN (n_67_99), .A (n_63_101), .B (n_57_104), .C1 (n_53_106), .C2 (n_47_109) );
AOI211_X1 g_68_101 (.ZN (n_68_101), .A (n_65_100), .B (n_59_103), .C1 (n_55_105), .C2 (n_49_108) );
AOI211_X1 g_66_102 (.ZN (n_66_102), .A (n_67_99), .B (n_61_102), .C1 (n_57_104), .C2 (n_51_107) );
AOI211_X1 g_64_101 (.ZN (n_64_101), .A (n_68_101), .B (n_63_101), .C1 (n_59_103), .C2 (n_53_106) );
AOI211_X1 g_62_102 (.ZN (n_62_102), .A (n_66_102), .B (n_65_100), .C1 (n_61_102), .C2 (n_55_105) );
AOI211_X1 g_60_103 (.ZN (n_60_103), .A (n_64_101), .B (n_67_99), .C1 (n_63_101), .C2 (n_57_104) );
AOI211_X1 g_58_104 (.ZN (n_58_104), .A (n_62_102), .B (n_68_101), .C1 (n_65_100), .C2 (n_59_103) );
AOI211_X1 g_56_105 (.ZN (n_56_105), .A (n_60_103), .B (n_66_102), .C1 (n_67_99), .C2 (n_61_102) );
AOI211_X1 g_54_106 (.ZN (n_54_106), .A (n_58_104), .B (n_64_101), .C1 (n_68_101), .C2 (n_63_101) );
AOI211_X1 g_52_107 (.ZN (n_52_107), .A (n_56_105), .B (n_62_102), .C1 (n_66_102), .C2 (n_65_100) );
AOI211_X1 g_50_108 (.ZN (n_50_108), .A (n_54_106), .B (n_60_103), .C1 (n_64_101), .C2 (n_67_99) );
AOI211_X1 g_48_109 (.ZN (n_48_109), .A (n_52_107), .B (n_58_104), .C1 (n_62_102), .C2 (n_68_101) );
AOI211_X1 g_46_110 (.ZN (n_46_110), .A (n_50_108), .B (n_56_105), .C1 (n_60_103), .C2 (n_66_102) );
AOI211_X1 g_44_111 (.ZN (n_44_111), .A (n_48_109), .B (n_54_106), .C1 (n_58_104), .C2 (n_64_101) );
AOI211_X1 g_42_112 (.ZN (n_42_112), .A (n_46_110), .B (n_52_107), .C1 (n_56_105), .C2 (n_62_102) );
AOI211_X1 g_40_113 (.ZN (n_40_113), .A (n_44_111), .B (n_50_108), .C1 (n_54_106), .C2 (n_60_103) );
AOI211_X1 g_38_114 (.ZN (n_38_114), .A (n_42_112), .B (n_48_109), .C1 (n_52_107), .C2 (n_58_104) );
AOI211_X1 g_36_115 (.ZN (n_36_115), .A (n_40_113), .B (n_46_110), .C1 (n_50_108), .C2 (n_56_105) );
AOI211_X1 g_34_116 (.ZN (n_34_116), .A (n_38_114), .B (n_44_111), .C1 (n_48_109), .C2 (n_54_106) );
AOI211_X1 g_32_117 (.ZN (n_32_117), .A (n_36_115), .B (n_42_112), .C1 (n_46_110), .C2 (n_52_107) );
AOI211_X1 g_30_118 (.ZN (n_30_118), .A (n_34_116), .B (n_40_113), .C1 (n_44_111), .C2 (n_50_108) );
AOI211_X1 g_31_116 (.ZN (n_31_116), .A (n_32_117), .B (n_38_114), .C1 (n_42_112), .C2 (n_48_109) );
AOI211_X1 g_29_117 (.ZN (n_29_117), .A (n_30_118), .B (n_36_115), .C1 (n_40_113), .C2 (n_46_110) );
AOI211_X1 g_27_118 (.ZN (n_27_118), .A (n_31_116), .B (n_34_116), .C1 (n_38_114), .C2 (n_44_111) );
AOI211_X1 g_25_119 (.ZN (n_25_119), .A (n_29_117), .B (n_32_117), .C1 (n_36_115), .C2 (n_42_112) );
AOI211_X1 g_23_120 (.ZN (n_23_120), .A (n_27_118), .B (n_30_118), .C1 (n_34_116), .C2 (n_40_113) );
AOI211_X1 g_21_121 (.ZN (n_21_121), .A (n_25_119), .B (n_31_116), .C1 (n_32_117), .C2 (n_38_114) );
AOI211_X1 g_20_123 (.ZN (n_20_123), .A (n_23_120), .B (n_29_117), .C1 (n_30_118), .C2 (n_36_115) );
AOI211_X1 g_18_122 (.ZN (n_18_122), .A (n_21_121), .B (n_27_118), .C1 (n_31_116), .C2 (n_34_116) );
AOI211_X1 g_20_121 (.ZN (n_20_121), .A (n_20_123), .B (n_25_119), .C1 (n_29_117), .C2 (n_32_117) );
AOI211_X1 g_22_120 (.ZN (n_22_120), .A (n_18_122), .B (n_23_120), .C1 (n_27_118), .C2 (n_30_118) );
AOI211_X1 g_21_122 (.ZN (n_21_122), .A (n_20_121), .B (n_21_121), .C1 (n_25_119), .C2 (n_31_116) );
AOI211_X1 g_23_121 (.ZN (n_23_121), .A (n_22_120), .B (n_20_123), .C1 (n_23_120), .C2 (n_29_117) );
AOI211_X1 g_22_123 (.ZN (n_22_123), .A (n_21_122), .B (n_18_122), .C1 (n_21_121), .C2 (n_27_118) );
AOI211_X1 g_20_122 (.ZN (n_20_122), .A (n_23_121), .B (n_20_121), .C1 (n_20_123), .C2 (n_25_119) );
AOI211_X1 g_22_121 (.ZN (n_22_121), .A (n_22_123), .B (n_22_120), .C1 (n_18_122), .C2 (n_23_120) );
AOI211_X1 g_24_120 (.ZN (n_24_120), .A (n_20_122), .B (n_21_122), .C1 (n_20_121), .C2 (n_21_121) );
AOI211_X1 g_26_119 (.ZN (n_26_119), .A (n_22_121), .B (n_23_121), .C1 (n_22_120), .C2 (n_20_123) );
AOI211_X1 g_28_118 (.ZN (n_28_118), .A (n_24_120), .B (n_22_123), .C1 (n_21_122), .C2 (n_18_122) );
AOI211_X1 g_30_117 (.ZN (n_30_117), .A (n_26_119), .B (n_20_122), .C1 (n_23_121), .C2 (n_20_121) );
AOI211_X1 g_32_116 (.ZN (n_32_116), .A (n_28_118), .B (n_22_121), .C1 (n_22_123), .C2 (n_22_120) );
AOI211_X1 g_34_115 (.ZN (n_34_115), .A (n_30_117), .B (n_24_120), .C1 (n_20_122), .C2 (n_21_122) );
AOI211_X1 g_36_114 (.ZN (n_36_114), .A (n_32_116), .B (n_26_119), .C1 (n_22_121), .C2 (n_23_121) );
AOI211_X1 g_38_113 (.ZN (n_38_113), .A (n_34_115), .B (n_28_118), .C1 (n_24_120), .C2 (n_22_123) );
AOI211_X1 g_40_112 (.ZN (n_40_112), .A (n_36_114), .B (n_30_117), .C1 (n_26_119), .C2 (n_20_122) );
AOI211_X1 g_42_111 (.ZN (n_42_111), .A (n_38_113), .B (n_32_116), .C1 (n_28_118), .C2 (n_22_121) );
AOI211_X1 g_44_110 (.ZN (n_44_110), .A (n_40_112), .B (n_34_115), .C1 (n_30_117), .C2 (n_24_120) );
AOI211_X1 g_46_109 (.ZN (n_46_109), .A (n_42_111), .B (n_36_114), .C1 (n_32_116), .C2 (n_26_119) );
AOI211_X1 g_45_111 (.ZN (n_45_111), .A (n_44_110), .B (n_38_113), .C1 (n_34_115), .C2 (n_28_118) );
AOI211_X1 g_47_110 (.ZN (n_47_110), .A (n_46_109), .B (n_40_112), .C1 (n_36_114), .C2 (n_30_117) );
AOI211_X1 g_49_109 (.ZN (n_49_109), .A (n_45_111), .B (n_42_111), .C1 (n_38_113), .C2 (n_32_116) );
AOI211_X1 g_51_108 (.ZN (n_51_108), .A (n_47_110), .B (n_44_110), .C1 (n_40_112), .C2 (n_34_115) );
AOI211_X1 g_53_107 (.ZN (n_53_107), .A (n_49_109), .B (n_46_109), .C1 (n_42_111), .C2 (n_36_114) );
AOI211_X1 g_55_106 (.ZN (n_55_106), .A (n_51_108), .B (n_45_111), .C1 (n_44_110), .C2 (n_38_113) );
AOI211_X1 g_57_105 (.ZN (n_57_105), .A (n_53_107), .B (n_47_110), .C1 (n_46_109), .C2 (n_40_112) );
AOI211_X1 g_59_104 (.ZN (n_59_104), .A (n_55_106), .B (n_49_109), .C1 (n_45_111), .C2 (n_42_111) );
AOI211_X1 g_61_103 (.ZN (n_61_103), .A (n_57_105), .B (n_51_108), .C1 (n_47_110), .C2 (n_44_110) );
AOI211_X1 g_63_102 (.ZN (n_63_102), .A (n_59_104), .B (n_53_107), .C1 (n_49_109), .C2 (n_46_109) );
AOI211_X1 g_65_101 (.ZN (n_65_101), .A (n_61_103), .B (n_55_106), .C1 (n_51_108), .C2 (n_45_111) );
AOI211_X1 g_64_103 (.ZN (n_64_103), .A (n_63_102), .B (n_57_105), .C1 (n_53_107), .C2 (n_47_110) );
AOI211_X1 g_62_104 (.ZN (n_62_104), .A (n_65_101), .B (n_59_104), .C1 (n_55_106), .C2 (n_49_109) );
AOI211_X1 g_60_105 (.ZN (n_60_105), .A (n_64_103), .B (n_61_103), .C1 (n_57_105), .C2 (n_51_108) );
AOI211_X1 g_58_106 (.ZN (n_58_106), .A (n_62_104), .B (n_63_102), .C1 (n_59_104), .C2 (n_53_107) );
AOI211_X1 g_56_107 (.ZN (n_56_107), .A (n_60_105), .B (n_65_101), .C1 (n_61_103), .C2 (n_55_106) );
AOI211_X1 g_54_108 (.ZN (n_54_108), .A (n_58_106), .B (n_64_103), .C1 (n_63_102), .C2 (n_57_105) );
AOI211_X1 g_52_109 (.ZN (n_52_109), .A (n_56_107), .B (n_62_104), .C1 (n_65_101), .C2 (n_59_104) );
AOI211_X1 g_50_110 (.ZN (n_50_110), .A (n_54_108), .B (n_60_105), .C1 (n_64_103), .C2 (n_61_103) );
AOI211_X1 g_48_111 (.ZN (n_48_111), .A (n_52_109), .B (n_58_106), .C1 (n_62_104), .C2 (n_63_102) );
AOI211_X1 g_46_112 (.ZN (n_46_112), .A (n_50_110), .B (n_56_107), .C1 (n_60_105), .C2 (n_65_101) );
AOI211_X1 g_44_113 (.ZN (n_44_113), .A (n_48_111), .B (n_54_108), .C1 (n_58_106), .C2 (n_64_103) );
AOI211_X1 g_42_114 (.ZN (n_42_114), .A (n_46_112), .B (n_52_109), .C1 (n_56_107), .C2 (n_62_104) );
AOI211_X1 g_43_112 (.ZN (n_43_112), .A (n_44_113), .B (n_50_110), .C1 (n_54_108), .C2 (n_60_105) );
AOI211_X1 g_41_113 (.ZN (n_41_113), .A (n_42_114), .B (n_48_111), .C1 (n_52_109), .C2 (n_58_106) );
AOI211_X1 g_39_114 (.ZN (n_39_114), .A (n_43_112), .B (n_46_112), .C1 (n_50_110), .C2 (n_56_107) );
AOI211_X1 g_37_115 (.ZN (n_37_115), .A (n_41_113), .B (n_44_113), .C1 (n_48_111), .C2 (n_54_108) );
AOI211_X1 g_35_116 (.ZN (n_35_116), .A (n_39_114), .B (n_42_114), .C1 (n_46_112), .C2 (n_52_109) );
AOI211_X1 g_33_117 (.ZN (n_33_117), .A (n_37_115), .B (n_43_112), .C1 (n_44_113), .C2 (n_50_110) );
AOI211_X1 g_31_118 (.ZN (n_31_118), .A (n_35_116), .B (n_41_113), .C1 (n_42_114), .C2 (n_48_111) );
AOI211_X1 g_29_119 (.ZN (n_29_119), .A (n_33_117), .B (n_39_114), .C1 (n_43_112), .C2 (n_46_112) );
AOI211_X1 g_27_120 (.ZN (n_27_120), .A (n_31_118), .B (n_37_115), .C1 (n_41_113), .C2 (n_44_113) );
AOI211_X1 g_25_121 (.ZN (n_25_121), .A (n_29_119), .B (n_35_116), .C1 (n_39_114), .C2 (n_42_114) );
AOI211_X1 g_23_122 (.ZN (n_23_122), .A (n_27_120), .B (n_33_117), .C1 (n_37_115), .C2 (n_43_112) );
AOI211_X1 g_21_123 (.ZN (n_21_123), .A (n_25_121), .B (n_31_118), .C1 (n_35_116), .C2 (n_41_113) );
AOI211_X1 g_19_124 (.ZN (n_19_124), .A (n_23_122), .B (n_29_119), .C1 (n_33_117), .C2 (n_39_114) );
AOI211_X1 g_17_123 (.ZN (n_17_123), .A (n_21_123), .B (n_27_120), .C1 (n_31_118), .C2 (n_37_115) );
AOI211_X1 g_15_122 (.ZN (n_15_122), .A (n_19_124), .B (n_25_121), .C1 (n_29_119), .C2 (n_35_116) );
AOI211_X1 g_13_123 (.ZN (n_13_123), .A (n_17_123), .B (n_23_122), .C1 (n_27_120), .C2 (n_33_117) );
AOI211_X1 g_11_124 (.ZN (n_11_124), .A (n_15_122), .B (n_21_123), .C1 (n_25_121), .C2 (n_31_118) );
AOI211_X1 g_9_125 (.ZN (n_9_125), .A (n_13_123), .B (n_19_124), .C1 (n_23_122), .C2 (n_29_119) );
AOI211_X1 g_7_126 (.ZN (n_7_126), .A (n_11_124), .B (n_17_123), .C1 (n_21_123), .C2 (n_27_120) );
AOI211_X1 g_5_127 (.ZN (n_5_127), .A (n_9_125), .B (n_15_122), .C1 (n_19_124), .C2 (n_25_121) );
AOI211_X1 g_3_128 (.ZN (n_3_128), .A (n_7_126), .B (n_13_123), .C1 (n_17_123), .C2 (n_23_122) );
AOI211_X1 g_2_130 (.ZN (n_2_130), .A (n_5_127), .B (n_11_124), .C1 (n_15_122), .C2 (n_21_123) );
AOI211_X1 g_1_132 (.ZN (n_1_132), .A (n_3_128), .B (n_9_125), .C1 (n_13_123), .C2 (n_19_124) );
AOI211_X1 g_3_131 (.ZN (n_3_131), .A (n_2_130), .B (n_7_126), .C1 (n_11_124), .C2 (n_17_123) );
AOI211_X1 g_4_129 (.ZN (n_4_129), .A (n_1_132), .B (n_5_127), .C1 (n_9_125), .C2 (n_15_122) );
AOI211_X1 g_6_128 (.ZN (n_6_128), .A (n_3_131), .B (n_3_128), .C1 (n_7_126), .C2 (n_13_123) );
AOI211_X1 g_4_127 (.ZN (n_4_127), .A (n_4_129), .B (n_2_130), .C1 (n_5_127), .C2 (n_11_124) );
AOI211_X1 g_3_129 (.ZN (n_3_129), .A (n_6_128), .B (n_1_132), .C1 (n_3_128), .C2 (n_9_125) );
AOI211_X1 g_5_130 (.ZN (n_5_130), .A (n_4_127), .B (n_3_131), .C1 (n_2_130), .C2 (n_7_126) );
AOI211_X1 g_7_129 (.ZN (n_7_129), .A (n_3_129), .B (n_4_129), .C1 (n_1_132), .C2 (n_5_127) );
AOI211_X1 g_8_127 (.ZN (n_8_127), .A (n_5_130), .B (n_6_128), .C1 (n_3_131), .C2 (n_3_128) );
AOI211_X1 g_6_126 (.ZN (n_6_126), .A (n_7_129), .B (n_4_127), .C1 (n_4_129), .C2 (n_2_130) );
AOI211_X1 g_8_125 (.ZN (n_8_125), .A (n_8_127), .B (n_3_129), .C1 (n_6_128), .C2 (n_1_132) );
AOI211_X1 g_10_126 (.ZN (n_10_126), .A (n_6_126), .B (n_5_130), .C1 (n_4_127), .C2 (n_3_131) );
AOI211_X1 g_12_125 (.ZN (n_12_125), .A (n_8_125), .B (n_7_129), .C1 (n_3_129), .C2 (n_4_129) );
AOI211_X1 g_14_124 (.ZN (n_14_124), .A (n_10_126), .B (n_8_127), .C1 (n_5_130), .C2 (n_6_128) );
AOI211_X1 g_12_123 (.ZN (n_12_123), .A (n_12_125), .B (n_6_126), .C1 (n_7_129), .C2 (n_4_127) );
AOI211_X1 g_11_125 (.ZN (n_11_125), .A (n_14_124), .B (n_8_125), .C1 (n_8_127), .C2 (n_3_129) );
AOI211_X1 g_13_124 (.ZN (n_13_124), .A (n_12_123), .B (n_10_126), .C1 (n_6_126), .C2 (n_5_130) );
AOI211_X1 g_15_123 (.ZN (n_15_123), .A (n_11_125), .B (n_12_125), .C1 (n_8_125), .C2 (n_7_129) );
AOI211_X1 g_17_122 (.ZN (n_17_122), .A (n_13_124), .B (n_14_124), .C1 (n_10_126), .C2 (n_8_127) );
AOI211_X1 g_19_123 (.ZN (n_19_123), .A (n_15_123), .B (n_12_123), .C1 (n_12_125), .C2 (n_6_126) );
AOI211_X1 g_17_124 (.ZN (n_17_124), .A (n_17_122), .B (n_11_125), .C1 (n_14_124), .C2 (n_8_125) );
AOI211_X1 g_15_125 (.ZN (n_15_125), .A (n_19_123), .B (n_13_124), .C1 (n_12_123), .C2 (n_10_126) );
AOI211_X1 g_16_123 (.ZN (n_16_123), .A (n_17_124), .B (n_15_123), .C1 (n_11_125), .C2 (n_12_125) );
AOI211_X1 g_18_124 (.ZN (n_18_124), .A (n_15_125), .B (n_17_122), .C1 (n_13_124), .C2 (n_14_124) );
AOI211_X1 g_16_125 (.ZN (n_16_125), .A (n_16_123), .B (n_19_123), .C1 (n_15_123), .C2 (n_12_123) );
AOI211_X1 g_14_126 (.ZN (n_14_126), .A (n_18_124), .B (n_17_124), .C1 (n_17_122), .C2 (n_11_125) );
AOI211_X1 g_15_124 (.ZN (n_15_124), .A (n_16_125), .B (n_15_125), .C1 (n_19_123), .C2 (n_13_124) );
AOI211_X1 g_13_125 (.ZN (n_13_125), .A (n_14_126), .B (n_16_123), .C1 (n_17_124), .C2 (n_15_123) );
AOI211_X1 g_11_126 (.ZN (n_11_126), .A (n_15_124), .B (n_18_124), .C1 (n_15_125), .C2 (n_17_122) );
AOI211_X1 g_9_127 (.ZN (n_9_127), .A (n_13_125), .B (n_16_125), .C1 (n_16_123), .C2 (n_19_123) );
AOI211_X1 g_7_128 (.ZN (n_7_128), .A (n_11_126), .B (n_14_126), .C1 (n_18_124), .C2 (n_17_124) );
AOI211_X1 g_5_129 (.ZN (n_5_129), .A (n_9_127), .B (n_15_124), .C1 (n_16_125), .C2 (n_15_125) );
AOI211_X1 g_4_131 (.ZN (n_4_131), .A (n_7_128), .B (n_13_125), .C1 (n_14_126), .C2 (n_16_123) );
AOI211_X1 g_3_133 (.ZN (n_3_133), .A (n_5_129), .B (n_11_126), .C1 (n_15_124), .C2 (n_18_124) );
AOI211_X1 g_5_134 (.ZN (n_5_134), .A (n_4_131), .B (n_9_127), .C1 (n_13_125), .C2 (n_16_125) );
AOI211_X1 g_3_135 (.ZN (n_3_135), .A (n_3_133), .B (n_7_128), .C1 (n_11_126), .C2 (n_14_126) );
AOI211_X1 g_1_136 (.ZN (n_1_136), .A (n_5_134), .B (n_5_129), .C1 (n_9_127), .C2 (n_15_124) );
AOI211_X1 g_2_134 (.ZN (n_2_134), .A (n_3_135), .B (n_4_131), .C1 (n_7_128), .C2 (n_13_125) );
AOI211_X1 g_4_133 (.ZN (n_4_133), .A (n_1_136), .B (n_3_133), .C1 (n_5_129), .C2 (n_11_126) );
AOI211_X1 g_6_132 (.ZN (n_6_132), .A (n_2_134), .B (n_5_134), .C1 (n_4_131), .C2 (n_9_127) );
AOI211_X1 g_7_130 (.ZN (n_7_130), .A (n_4_133), .B (n_3_135), .C1 (n_3_133), .C2 (n_7_128) );
AOI211_X1 g_5_131 (.ZN (n_5_131), .A (n_6_132), .B (n_1_136), .C1 (n_5_134), .C2 (n_5_129) );
AOI211_X1 g_3_132 (.ZN (n_3_132), .A (n_7_130), .B (n_2_134), .C1 (n_3_135), .C2 (n_4_131) );
AOI211_X1 g_4_130 (.ZN (n_4_130), .A (n_5_131), .B (n_4_133), .C1 (n_1_136), .C2 (n_3_133) );
AOI211_X1 g_5_128 (.ZN (n_5_128), .A (n_3_132), .B (n_6_132), .C1 (n_2_134), .C2 (n_5_134) );
AOI211_X1 g_7_127 (.ZN (n_7_127), .A (n_4_130), .B (n_7_130), .C1 (n_4_133), .C2 (n_3_135) );
AOI211_X1 g_9_126 (.ZN (n_9_126), .A (n_5_128), .B (n_5_131), .C1 (n_6_132), .C2 (n_1_136) );
AOI211_X1 g_8_128 (.ZN (n_8_128), .A (n_7_127), .B (n_3_132), .C1 (n_7_130), .C2 (n_2_134) );
AOI211_X1 g_6_129 (.ZN (n_6_129), .A (n_9_126), .B (n_4_130), .C1 (n_5_131), .C2 (n_4_133) );
AOI211_X1 g_7_131 (.ZN (n_7_131), .A (n_8_128), .B (n_5_128), .C1 (n_3_132), .C2 (n_6_132) );
AOI211_X1 g_8_129 (.ZN (n_8_129), .A (n_6_129), .B (n_7_127), .C1 (n_4_130), .C2 (n_7_130) );
AOI211_X1 g_6_130 (.ZN (n_6_130), .A (n_7_131), .B (n_9_126), .C1 (n_5_128), .C2 (n_5_131) );
AOI211_X1 g_5_132 (.ZN (n_5_132), .A (n_8_129), .B (n_8_128), .C1 (n_7_127), .C2 (n_3_132) );
AOI211_X1 g_4_134 (.ZN (n_4_134), .A (n_6_130), .B (n_6_129), .C1 (n_9_126), .C2 (n_4_130) );
AOI211_X1 g_6_133 (.ZN (n_6_133), .A (n_5_132), .B (n_7_131), .C1 (n_8_128), .C2 (n_5_128) );
AOI211_X1 g_5_135 (.ZN (n_5_135), .A (n_4_134), .B (n_8_129), .C1 (n_6_129), .C2 (n_7_127) );
AOI211_X1 g_3_136 (.ZN (n_3_136), .A (n_6_133), .B (n_6_130), .C1 (n_7_131), .C2 (n_9_126) );
AOI211_X1 g_2_138 (.ZN (n_2_138), .A (n_5_135), .B (n_5_132), .C1 (n_8_129), .C2 (n_8_128) );
AOI211_X1 g_1_140 (.ZN (n_1_140), .A (n_3_136), .B (n_4_134), .C1 (n_6_130), .C2 (n_6_129) );
AOI211_X1 g_3_139 (.ZN (n_3_139), .A (n_2_138), .B (n_6_133), .C1 (n_5_132), .C2 (n_7_131) );
AOI211_X1 g_4_137 (.ZN (n_4_137), .A (n_1_140), .B (n_5_135), .C1 (n_4_134), .C2 (n_8_129) );
AOI211_X1 g_6_136 (.ZN (n_6_136), .A (n_3_139), .B (n_3_136), .C1 (n_6_133), .C2 (n_6_130) );
AOI211_X1 g_4_135 (.ZN (n_4_135), .A (n_4_137), .B (n_2_138), .C1 (n_5_135), .C2 (n_5_132) );
AOI211_X1 g_3_137 (.ZN (n_3_137), .A (n_6_136), .B (n_1_140), .C1 (n_3_136), .C2 (n_4_134) );
AOI211_X1 g_5_138 (.ZN (n_5_138), .A (n_4_135), .B (n_3_139), .C1 (n_2_138), .C2 (n_6_133) );
AOI211_X1 g_7_137 (.ZN (n_7_137), .A (n_3_137), .B (n_4_137), .C1 (n_1_140), .C2 (n_5_135) );
AOI211_X1 g_5_136 (.ZN (n_5_136), .A (n_5_138), .B (n_6_136), .C1 (n_3_139), .C2 (n_3_136) );
AOI211_X1 g_6_134 (.ZN (n_6_134), .A (n_7_137), .B (n_4_135), .C1 (n_4_137), .C2 (n_2_138) );
AOI211_X1 g_8_133 (.ZN (n_8_133), .A (n_5_136), .B (n_3_137), .C1 (n_6_136), .C2 (n_1_140) );
AOI211_X1 g_7_135 (.ZN (n_7_135), .A (n_6_134), .B (n_5_138), .C1 (n_4_135), .C2 (n_3_139) );
AOI211_X1 g_6_137 (.ZN (n_6_137), .A (n_8_133), .B (n_7_137), .C1 (n_3_137), .C2 (n_4_137) );
AOI211_X1 g_4_138 (.ZN (n_4_138), .A (n_7_135), .B (n_5_136), .C1 (n_5_138), .C2 (n_6_136) );
AOI211_X1 g_3_140 (.ZN (n_3_140), .A (n_6_137), .B (n_6_134), .C1 (n_7_137), .C2 (n_4_135) );
AOI211_X1 g_5_139 (.ZN (n_5_139), .A (n_4_138), .B (n_8_133), .C1 (n_5_136), .C2 (n_3_137) );
AOI211_X1 g_4_141 (.ZN (n_4_141), .A (n_3_140), .B (n_7_135), .C1 (n_6_134), .C2 (n_5_138) );
AOI211_X1 g_2_142 (.ZN (n_2_142), .A (n_5_139), .B (n_6_137), .C1 (n_8_133), .C2 (n_7_137) );
AOI211_X1 g_1_144 (.ZN (n_1_144), .A (n_4_141), .B (n_4_138), .C1 (n_7_135), .C2 (n_5_136) );
AOI211_X1 g_3_143 (.ZN (n_3_143), .A (n_2_142), .B (n_3_140), .C1 (n_6_137), .C2 (n_6_134) );
AOI211_X1 g_5_142 (.ZN (n_5_142), .A (n_1_144), .B (n_5_139), .C1 (n_4_138), .C2 (n_8_133) );
AOI211_X1 g_3_141 (.ZN (n_3_141), .A (n_3_143), .B (n_4_141), .C1 (n_3_140), .C2 (n_7_135) );
AOI211_X1 g_4_139 (.ZN (n_4_139), .A (n_5_142), .B (n_2_142), .C1 (n_5_139), .C2 (n_6_137) );
AOI211_X1 g_5_137 (.ZN (n_5_137), .A (n_3_141), .B (n_1_144), .C1 (n_4_141), .C2 (n_4_138) );
AOI211_X1 g_6_135 (.ZN (n_6_135), .A (n_4_139), .B (n_3_143), .C1 (n_2_142), .C2 (n_3_140) );
AOI211_X1 g_5_133 (.ZN (n_5_133), .A (n_5_137), .B (n_5_142), .C1 (n_1_144), .C2 (n_5_139) );
AOI211_X1 g_6_131 (.ZN (n_6_131), .A (n_6_135), .B (n_3_141), .C1 (n_3_143), .C2 (n_4_141) );
AOI211_X1 g_7_133 (.ZN (n_7_133), .A (n_5_133), .B (n_4_139), .C1 (n_5_142), .C2 (n_2_142) );
AOI211_X1 g_8_131 (.ZN (n_8_131), .A (n_6_131), .B (n_5_137), .C1 (n_3_141), .C2 (n_1_144) );
AOI211_X1 g_9_129 (.ZN (n_9_129), .A (n_7_133), .B (n_6_135), .C1 (n_4_139), .C2 (n_3_143) );
AOI211_X1 g_10_127 (.ZN (n_10_127), .A (n_8_131), .B (n_5_133), .C1 (n_5_137), .C2 (n_5_142) );
AOI211_X1 g_12_126 (.ZN (n_12_126), .A (n_9_129), .B (n_6_131), .C1 (n_6_135), .C2 (n_3_141) );
AOI211_X1 g_14_125 (.ZN (n_14_125), .A (n_10_127), .B (n_7_133), .C1 (n_5_133), .C2 (n_4_139) );
AOI211_X1 g_16_124 (.ZN (n_16_124), .A (n_12_126), .B (n_8_131), .C1 (n_6_131), .C2 (n_5_137) );
AOI211_X1 g_18_123 (.ZN (n_18_123), .A (n_14_125), .B (n_9_129), .C1 (n_7_133), .C2 (n_6_135) );
AOI211_X1 g_17_125 (.ZN (n_17_125), .A (n_16_124), .B (n_10_127), .C1 (n_8_131), .C2 (n_5_133) );
AOI211_X1 g_15_126 (.ZN (n_15_126), .A (n_18_123), .B (n_12_126), .C1 (n_9_129), .C2 (n_6_131) );
AOI211_X1 g_13_127 (.ZN (n_13_127), .A (n_17_125), .B (n_14_125), .C1 (n_10_127), .C2 (n_7_133) );
AOI211_X1 g_11_128 (.ZN (n_11_128), .A (n_15_126), .B (n_16_124), .C1 (n_12_126), .C2 (n_8_131) );
AOI211_X1 g_10_130 (.ZN (n_10_130), .A (n_13_127), .B (n_18_123), .C1 (n_14_125), .C2 (n_9_129) );
AOI211_X1 g_9_128 (.ZN (n_9_128), .A (n_11_128), .B (n_17_125), .C1 (n_16_124), .C2 (n_10_127) );
AOI211_X1 g_11_127 (.ZN (n_11_127), .A (n_10_130), .B (n_15_126), .C1 (n_18_123), .C2 (n_12_126) );
AOI211_X1 g_13_126 (.ZN (n_13_126), .A (n_9_128), .B (n_13_127), .C1 (n_17_125), .C2 (n_14_125) );
AOI211_X1 g_12_128 (.ZN (n_12_128), .A (n_11_127), .B (n_11_128), .C1 (n_15_126), .C2 (n_16_124) );
AOI211_X1 g_14_127 (.ZN (n_14_127), .A (n_13_126), .B (n_10_130), .C1 (n_13_127), .C2 (n_18_123) );
AOI211_X1 g_16_126 (.ZN (n_16_126), .A (n_12_128), .B (n_9_128), .C1 (n_11_128), .C2 (n_17_125) );
AOI211_X1 g_18_125 (.ZN (n_18_125), .A (n_14_127), .B (n_11_127), .C1 (n_10_130), .C2 (n_15_126) );
AOI211_X1 g_20_124 (.ZN (n_20_124), .A (n_16_126), .B (n_13_126), .C1 (n_9_128), .C2 (n_13_127) );
AOI211_X1 g_19_126 (.ZN (n_19_126), .A (n_18_125), .B (n_12_128), .C1 (n_11_127), .C2 (n_11_128) );
AOI211_X1 g_21_125 (.ZN (n_21_125), .A (n_20_124), .B (n_14_127), .C1 (n_13_126), .C2 (n_10_130) );
AOI211_X1 g_23_124 (.ZN (n_23_124), .A (n_19_126), .B (n_16_126), .C1 (n_12_128), .C2 (n_9_128) );
AOI211_X1 g_24_122 (.ZN (n_24_122), .A (n_21_125), .B (n_18_125), .C1 (n_14_127), .C2 (n_11_127) );
AOI211_X1 g_26_121 (.ZN (n_26_121), .A (n_23_124), .B (n_20_124), .C1 (n_16_126), .C2 (n_13_126) );
AOI211_X1 g_27_119 (.ZN (n_27_119), .A (n_24_122), .B (n_19_126), .C1 (n_18_125), .C2 (n_12_128) );
AOI211_X1 g_29_118 (.ZN (n_29_118), .A (n_26_121), .B (n_21_125), .C1 (n_20_124), .C2 (n_14_127) );
AOI211_X1 g_31_117 (.ZN (n_31_117), .A (n_27_119), .B (n_23_124), .C1 (n_19_126), .C2 (n_16_126) );
AOI211_X1 g_30_119 (.ZN (n_30_119), .A (n_29_118), .B (n_24_122), .C1 (n_21_125), .C2 (n_18_125) );
AOI211_X1 g_28_120 (.ZN (n_28_120), .A (n_31_117), .B (n_26_121), .C1 (n_23_124), .C2 (n_20_124) );
AOI211_X1 g_27_122 (.ZN (n_27_122), .A (n_30_119), .B (n_27_119), .C1 (n_24_122), .C2 (n_19_126) );
AOI211_X1 g_26_120 (.ZN (n_26_120), .A (n_28_120), .B (n_29_118), .C1 (n_26_121), .C2 (n_21_125) );
AOI211_X1 g_28_119 (.ZN (n_28_119), .A (n_27_122), .B (n_31_117), .C1 (n_27_119), .C2 (n_23_124) );
AOI211_X1 g_29_121 (.ZN (n_29_121), .A (n_26_120), .B (n_30_119), .C1 (n_29_118), .C2 (n_24_122) );
AOI211_X1 g_31_120 (.ZN (n_31_120), .A (n_28_119), .B (n_28_120), .C1 (n_31_117), .C2 (n_26_121) );
AOI211_X1 g_32_118 (.ZN (n_32_118), .A (n_29_121), .B (n_27_122), .C1 (n_30_119), .C2 (n_27_119) );
AOI211_X1 g_34_117 (.ZN (n_34_117), .A (n_31_120), .B (n_26_120), .C1 (n_28_120), .C2 (n_29_118) );
AOI211_X1 g_36_116 (.ZN (n_36_116), .A (n_32_118), .B (n_28_119), .C1 (n_27_122), .C2 (n_31_117) );
AOI211_X1 g_38_115 (.ZN (n_38_115), .A (n_34_117), .B (n_29_121), .C1 (n_26_120), .C2 (n_30_119) );
AOI211_X1 g_40_114 (.ZN (n_40_114), .A (n_36_116), .B (n_31_120), .C1 (n_28_119), .C2 (n_28_120) );
AOI211_X1 g_42_113 (.ZN (n_42_113), .A (n_38_115), .B (n_32_118), .C1 (n_29_121), .C2 (n_27_122) );
AOI211_X1 g_44_112 (.ZN (n_44_112), .A (n_40_114), .B (n_34_117), .C1 (n_31_120), .C2 (n_26_120) );
AOI211_X1 g_46_111 (.ZN (n_46_111), .A (n_42_113), .B (n_36_116), .C1 (n_32_118), .C2 (n_28_119) );
AOI211_X1 g_48_110 (.ZN (n_48_110), .A (n_44_112), .B (n_38_115), .C1 (n_34_117), .C2 (n_29_121) );
AOI211_X1 g_50_109 (.ZN (n_50_109), .A (n_46_111), .B (n_40_114), .C1 (n_36_116), .C2 (n_31_120) );
AOI211_X1 g_52_108 (.ZN (n_52_108), .A (n_48_110), .B (n_42_113), .C1 (n_38_115), .C2 (n_32_118) );
AOI211_X1 g_54_107 (.ZN (n_54_107), .A (n_50_109), .B (n_44_112), .C1 (n_40_114), .C2 (n_34_117) );
AOI211_X1 g_56_106 (.ZN (n_56_106), .A (n_52_108), .B (n_46_111), .C1 (n_42_113), .C2 (n_36_116) );
AOI211_X1 g_58_105 (.ZN (n_58_105), .A (n_54_107), .B (n_48_110), .C1 (n_44_112), .C2 (n_38_115) );
AOI211_X1 g_60_104 (.ZN (n_60_104), .A (n_56_106), .B (n_50_109), .C1 (n_46_111), .C2 (n_40_114) );
AOI211_X1 g_62_103 (.ZN (n_62_103), .A (n_58_105), .B (n_52_108), .C1 (n_48_110), .C2 (n_42_113) );
AOI211_X1 g_64_102 (.ZN (n_64_102), .A (n_60_104), .B (n_54_107), .C1 (n_50_109), .C2 (n_44_112) );
AOI211_X1 g_66_101 (.ZN (n_66_101), .A (n_62_103), .B (n_56_106), .C1 (n_52_108), .C2 (n_46_111) );
AOI211_X1 g_68_100 (.ZN (n_68_100), .A (n_64_102), .B (n_58_105), .C1 (n_54_107), .C2 (n_48_110) );
AOI211_X1 g_67_102 (.ZN (n_67_102), .A (n_66_101), .B (n_60_104), .C1 (n_56_106), .C2 (n_50_109) );
AOI211_X1 g_69_101 (.ZN (n_69_101), .A (n_68_100), .B (n_62_103), .C1 (n_58_105), .C2 (n_52_108) );
AOI211_X1 g_71_100 (.ZN (n_71_100), .A (n_67_102), .B (n_64_102), .C1 (n_60_104), .C2 (n_54_107) );
AOI211_X1 g_73_99 (.ZN (n_73_99), .A (n_69_101), .B (n_66_101), .C1 (n_62_103), .C2 (n_56_106) );
AOI211_X1 g_75_98 (.ZN (n_75_98), .A (n_71_100), .B (n_68_100), .C1 (n_64_102), .C2 (n_58_105) );
AOI211_X1 g_77_97 (.ZN (n_77_97), .A (n_73_99), .B (n_67_102), .C1 (n_66_101), .C2 (n_60_104) );
AOI211_X1 g_76_95 (.ZN (n_76_95), .A (n_75_98), .B (n_69_101), .C1 (n_68_100), .C2 (n_62_103) );
AOI211_X1 g_78_94 (.ZN (n_78_94), .A (n_77_97), .B (n_71_100), .C1 (n_67_102), .C2 (n_64_102) );
AOI211_X1 g_80_93 (.ZN (n_80_93), .A (n_76_95), .B (n_73_99), .C1 (n_69_101), .C2 (n_66_101) );
AOI211_X1 g_82_92 (.ZN (n_82_92), .A (n_78_94), .B (n_75_98), .C1 (n_71_100), .C2 (n_68_100) );
AOI211_X1 g_84_91 (.ZN (n_84_91), .A (n_80_93), .B (n_77_97), .C1 (n_73_99), .C2 (n_67_102) );
AOI211_X1 g_83_93 (.ZN (n_83_93), .A (n_82_92), .B (n_76_95), .C1 (n_75_98), .C2 (n_69_101) );
AOI211_X1 g_85_92 (.ZN (n_85_92), .A (n_84_91), .B (n_78_94), .C1 (n_77_97), .C2 (n_71_100) );
AOI211_X1 g_87_91 (.ZN (n_87_91), .A (n_83_93), .B (n_80_93), .C1 (n_76_95), .C2 (n_73_99) );
AOI211_X1 g_89_90 (.ZN (n_89_90), .A (n_85_92), .B (n_82_92), .C1 (n_78_94), .C2 (n_75_98) );
AOI211_X1 g_91_89 (.ZN (n_91_89), .A (n_87_91), .B (n_84_91), .C1 (n_80_93), .C2 (n_77_97) );
AOI211_X1 g_93_88 (.ZN (n_93_88), .A (n_89_90), .B (n_83_93), .C1 (n_82_92), .C2 (n_76_95) );
AOI211_X1 g_95_87 (.ZN (n_95_87), .A (n_91_89), .B (n_85_92), .C1 (n_84_91), .C2 (n_78_94) );
AOI211_X1 g_94_89 (.ZN (n_94_89), .A (n_93_88), .B (n_87_91), .C1 (n_83_93), .C2 (n_80_93) );
AOI211_X1 g_93_87 (.ZN (n_93_87), .A (n_95_87), .B (n_89_90), .C1 (n_85_92), .C2 (n_82_92) );
AOI211_X1 g_95_86 (.ZN (n_95_86), .A (n_94_89), .B (n_91_89), .C1 (n_87_91), .C2 (n_84_91) );
AOI211_X1 g_97_85 (.ZN (n_97_85), .A (n_93_87), .B (n_93_88), .C1 (n_89_90), .C2 (n_83_93) );
AOI211_X1 g_96_87 (.ZN (n_96_87), .A (n_95_86), .B (n_95_87), .C1 (n_91_89), .C2 (n_85_92) );
AOI211_X1 g_98_86 (.ZN (n_98_86), .A (n_97_85), .B (n_94_89), .C1 (n_93_88), .C2 (n_87_91) );
AOI211_X1 g_100_85 (.ZN (n_100_85), .A (n_96_87), .B (n_93_87), .C1 (n_95_87), .C2 (n_89_90) );
AOI211_X1 g_102_84 (.ZN (n_102_84), .A (n_98_86), .B (n_95_86), .C1 (n_94_89), .C2 (n_91_89) );
AOI211_X1 g_104_83 (.ZN (n_104_83), .A (n_100_85), .B (n_97_85), .C1 (n_93_87), .C2 (n_93_88) );
AOI211_X1 g_106_82 (.ZN (n_106_82), .A (n_102_84), .B (n_96_87), .C1 (n_95_86), .C2 (n_95_87) );
AOI211_X1 g_108_81 (.ZN (n_108_81), .A (n_104_83), .B (n_98_86), .C1 (n_97_85), .C2 (n_94_89) );
AOI211_X1 g_110_80 (.ZN (n_110_80), .A (n_106_82), .B (n_100_85), .C1 (n_96_87), .C2 (n_93_87) );
AOI211_X1 g_112_79 (.ZN (n_112_79), .A (n_108_81), .B (n_102_84), .C1 (n_98_86), .C2 (n_95_86) );
AOI211_X1 g_114_78 (.ZN (n_114_78), .A (n_110_80), .B (n_104_83), .C1 (n_100_85), .C2 (n_97_85) );
AOI211_X1 g_116_77 (.ZN (n_116_77), .A (n_112_79), .B (n_106_82), .C1 (n_102_84), .C2 (n_96_87) );
AOI211_X1 g_118_76 (.ZN (n_118_76), .A (n_114_78), .B (n_108_81), .C1 (n_104_83), .C2 (n_98_86) );
AOI211_X1 g_120_77 (.ZN (n_120_77), .A (n_116_77), .B (n_110_80), .C1 (n_106_82), .C2 (n_100_85) );
AOI211_X1 g_118_78 (.ZN (n_118_78), .A (n_118_76), .B (n_112_79), .C1 (n_108_81), .C2 (n_102_84) );
AOI211_X1 g_116_79 (.ZN (n_116_79), .A (n_120_77), .B (n_114_78), .C1 (n_110_80), .C2 (n_104_83) );
AOI211_X1 g_117_77 (.ZN (n_117_77), .A (n_118_78), .B (n_116_77), .C1 (n_112_79), .C2 (n_106_82) );
AOI211_X1 g_115_78 (.ZN (n_115_78), .A (n_116_79), .B (n_118_76), .C1 (n_114_78), .C2 (n_108_81) );
AOI211_X1 g_113_79 (.ZN (n_113_79), .A (n_117_77), .B (n_120_77), .C1 (n_116_77), .C2 (n_110_80) );
AOI211_X1 g_111_80 (.ZN (n_111_80), .A (n_115_78), .B (n_118_78), .C1 (n_118_76), .C2 (n_112_79) );
AOI211_X1 g_109_81 (.ZN (n_109_81), .A (n_113_79), .B (n_116_79), .C1 (n_120_77), .C2 (n_114_78) );
AOI211_X1 g_107_82 (.ZN (n_107_82), .A (n_111_80), .B (n_117_77), .C1 (n_118_78), .C2 (n_116_77) );
AOI211_X1 g_105_83 (.ZN (n_105_83), .A (n_109_81), .B (n_115_78), .C1 (n_116_79), .C2 (n_118_76) );
AOI211_X1 g_103_84 (.ZN (n_103_84), .A (n_107_82), .B (n_113_79), .C1 (n_117_77), .C2 (n_120_77) );
AOI211_X1 g_101_85 (.ZN (n_101_85), .A (n_105_83), .B (n_111_80), .C1 (n_115_78), .C2 (n_118_78) );
AOI211_X1 g_99_86 (.ZN (n_99_86), .A (n_103_84), .B (n_109_81), .C1 (n_113_79), .C2 (n_116_79) );
AOI211_X1 g_97_87 (.ZN (n_97_87), .A (n_101_85), .B (n_107_82), .C1 (n_111_80), .C2 (n_117_77) );
AOI211_X1 g_95_88 (.ZN (n_95_88), .A (n_99_86), .B (n_105_83), .C1 (n_109_81), .C2 (n_115_78) );
AOI211_X1 g_93_89 (.ZN (n_93_89), .A (n_97_87), .B (n_103_84), .C1 (n_107_82), .C2 (n_113_79) );
AOI211_X1 g_91_88 (.ZN (n_91_88), .A (n_95_88), .B (n_101_85), .C1 (n_105_83), .C2 (n_111_80) );
AOI211_X1 g_89_89 (.ZN (n_89_89), .A (n_93_89), .B (n_99_86), .C1 (n_103_84), .C2 (n_109_81) );
AOI211_X1 g_87_90 (.ZN (n_87_90), .A (n_91_88), .B (n_97_87), .C1 (n_101_85), .C2 (n_107_82) );
AOI211_X1 g_85_91 (.ZN (n_85_91), .A (n_89_89), .B (n_95_88), .C1 (n_99_86), .C2 (n_105_83) );
AOI211_X1 g_84_93 (.ZN (n_84_93), .A (n_87_90), .B (n_93_89), .C1 (n_97_87), .C2 (n_103_84) );
AOI211_X1 g_86_92 (.ZN (n_86_92), .A (n_85_91), .B (n_91_88), .C1 (n_95_88), .C2 (n_101_85) );
AOI211_X1 g_88_91 (.ZN (n_88_91), .A (n_84_93), .B (n_89_89), .C1 (n_93_89), .C2 (n_99_86) );
AOI211_X1 g_90_90 (.ZN (n_90_90), .A (n_86_92), .B (n_87_90), .C1 (n_91_88), .C2 (n_97_87) );
AOI211_X1 g_92_89 (.ZN (n_92_89), .A (n_88_91), .B (n_85_91), .C1 (n_89_89), .C2 (n_95_88) );
AOI211_X1 g_94_88 (.ZN (n_94_88), .A (n_90_90), .B (n_84_93), .C1 (n_87_90), .C2 (n_93_89) );
AOI211_X1 g_93_90 (.ZN (n_93_90), .A (n_92_89), .B (n_86_92), .C1 (n_85_91), .C2 (n_91_88) );
AOI211_X1 g_95_89 (.ZN (n_95_89), .A (n_94_88), .B (n_88_91), .C1 (n_84_93), .C2 (n_89_89) );
AOI211_X1 g_97_88 (.ZN (n_97_88), .A (n_93_90), .B (n_90_90), .C1 (n_86_92), .C2 (n_87_90) );
AOI211_X1 g_99_87 (.ZN (n_99_87), .A (n_95_89), .B (n_92_89), .C1 (n_88_91), .C2 (n_85_91) );
AOI211_X1 g_101_86 (.ZN (n_101_86), .A (n_97_88), .B (n_94_88), .C1 (n_90_90), .C2 (n_84_93) );
AOI211_X1 g_103_85 (.ZN (n_103_85), .A (n_99_87), .B (n_93_90), .C1 (n_92_89), .C2 (n_86_92) );
AOI211_X1 g_105_84 (.ZN (n_105_84), .A (n_101_86), .B (n_95_89), .C1 (n_94_88), .C2 (n_88_91) );
AOI211_X1 g_107_83 (.ZN (n_107_83), .A (n_103_85), .B (n_97_88), .C1 (n_93_90), .C2 (n_90_90) );
AOI211_X1 g_109_82 (.ZN (n_109_82), .A (n_105_84), .B (n_99_87), .C1 (n_95_89), .C2 (n_92_89) );
AOI211_X1 g_111_81 (.ZN (n_111_81), .A (n_107_83), .B (n_101_86), .C1 (n_97_88), .C2 (n_94_88) );
AOI211_X1 g_113_80 (.ZN (n_113_80), .A (n_109_82), .B (n_103_85), .C1 (n_99_87), .C2 (n_93_90) );
AOI211_X1 g_115_79 (.ZN (n_115_79), .A (n_111_81), .B (n_105_84), .C1 (n_101_86), .C2 (n_95_89) );
AOI211_X1 g_117_78 (.ZN (n_117_78), .A (n_113_80), .B (n_107_83), .C1 (n_103_85), .C2 (n_97_88) );
AOI211_X1 g_119_77 (.ZN (n_119_77), .A (n_115_79), .B (n_109_82), .C1 (n_105_84), .C2 (n_99_87) );
AOI211_X1 g_121_76 (.ZN (n_121_76), .A (n_117_78), .B (n_111_81), .C1 (n_107_83), .C2 (n_101_86) );
AOI211_X1 g_123_75 (.ZN (n_123_75), .A (n_119_77), .B (n_113_80), .C1 (n_109_82), .C2 (n_103_85) );
AOI211_X1 g_124_77 (.ZN (n_124_77), .A (n_121_76), .B (n_115_79), .C1 (n_111_81), .C2 (n_105_84) );
AOI211_X1 g_122_78 (.ZN (n_122_78), .A (n_123_75), .B (n_117_78), .C1 (n_113_80), .C2 (n_107_83) );
AOI211_X1 g_120_79 (.ZN (n_120_79), .A (n_124_77), .B (n_119_77), .C1 (n_115_79), .C2 (n_109_82) );
AOI211_X1 g_121_77 (.ZN (n_121_77), .A (n_122_78), .B (n_121_76), .C1 (n_117_78), .C2 (n_111_81) );
AOI211_X1 g_119_78 (.ZN (n_119_78), .A (n_120_79), .B (n_123_75), .C1 (n_119_77), .C2 (n_113_80) );
AOI211_X1 g_117_79 (.ZN (n_117_79), .A (n_121_77), .B (n_124_77), .C1 (n_121_76), .C2 (n_115_79) );
AOI211_X1 g_115_80 (.ZN (n_115_80), .A (n_119_78), .B (n_122_78), .C1 (n_123_75), .C2 (n_117_78) );
AOI211_X1 g_116_78 (.ZN (n_116_78), .A (n_117_79), .B (n_120_79), .C1 (n_124_77), .C2 (n_119_77) );
AOI211_X1 g_114_79 (.ZN (n_114_79), .A (n_115_80), .B (n_121_77), .C1 (n_122_78), .C2 (n_121_76) );
AOI211_X1 g_112_80 (.ZN (n_112_80), .A (n_116_78), .B (n_119_78), .C1 (n_120_79), .C2 (n_123_75) );
AOI211_X1 g_110_81 (.ZN (n_110_81), .A (n_114_79), .B (n_117_79), .C1 (n_121_77), .C2 (n_124_77) );
AOI211_X1 g_108_82 (.ZN (n_108_82), .A (n_112_80), .B (n_115_80), .C1 (n_119_78), .C2 (n_122_78) );
AOI211_X1 g_106_83 (.ZN (n_106_83), .A (n_110_81), .B (n_116_78), .C1 (n_117_79), .C2 (n_120_79) );
AOI211_X1 g_104_84 (.ZN (n_104_84), .A (n_108_82), .B (n_114_79), .C1 (n_115_80), .C2 (n_121_77) );
AOI211_X1 g_102_85 (.ZN (n_102_85), .A (n_106_83), .B (n_112_80), .C1 (n_116_78), .C2 (n_119_78) );
AOI211_X1 g_100_86 (.ZN (n_100_86), .A (n_104_84), .B (n_110_81), .C1 (n_114_79), .C2 (n_117_79) );
AOI211_X1 g_98_87 (.ZN (n_98_87), .A (n_102_85), .B (n_108_82), .C1 (n_112_80), .C2 (n_115_80) );
AOI211_X1 g_96_88 (.ZN (n_96_88), .A (n_100_86), .B (n_106_83), .C1 (n_110_81), .C2 (n_116_78) );
AOI211_X1 g_95_90 (.ZN (n_95_90), .A (n_98_87), .B (n_104_84), .C1 (n_108_82), .C2 (n_114_79) );
AOI211_X1 g_97_89 (.ZN (n_97_89), .A (n_96_88), .B (n_102_85), .C1 (n_106_83), .C2 (n_112_80) );
AOI211_X1 g_99_88 (.ZN (n_99_88), .A (n_95_90), .B (n_100_86), .C1 (n_104_84), .C2 (n_110_81) );
AOI211_X1 g_101_87 (.ZN (n_101_87), .A (n_97_89), .B (n_98_87), .C1 (n_102_85), .C2 (n_108_82) );
AOI211_X1 g_103_86 (.ZN (n_103_86), .A (n_99_88), .B (n_96_88), .C1 (n_100_86), .C2 (n_106_83) );
AOI211_X1 g_105_85 (.ZN (n_105_85), .A (n_101_87), .B (n_95_90), .C1 (n_98_87), .C2 (n_104_84) );
AOI211_X1 g_107_84 (.ZN (n_107_84), .A (n_103_86), .B (n_97_89), .C1 (n_96_88), .C2 (n_102_85) );
AOI211_X1 g_109_83 (.ZN (n_109_83), .A (n_105_85), .B (n_99_88), .C1 (n_95_90), .C2 (n_100_86) );
AOI211_X1 g_111_82 (.ZN (n_111_82), .A (n_107_84), .B (n_101_87), .C1 (n_97_89), .C2 (n_98_87) );
AOI211_X1 g_113_81 (.ZN (n_113_81), .A (n_109_83), .B (n_103_86), .C1 (n_99_88), .C2 (n_96_88) );
AOI211_X1 g_112_83 (.ZN (n_112_83), .A (n_111_82), .B (n_105_85), .C1 (n_101_87), .C2 (n_95_90) );
AOI211_X1 g_110_82 (.ZN (n_110_82), .A (n_113_81), .B (n_107_84), .C1 (n_103_86), .C2 (n_97_89) );
AOI211_X1 g_112_81 (.ZN (n_112_81), .A (n_112_83), .B (n_109_83), .C1 (n_105_85), .C2 (n_99_88) );
AOI211_X1 g_114_80 (.ZN (n_114_80), .A (n_110_82), .B (n_111_82), .C1 (n_107_84), .C2 (n_101_87) );
AOI211_X1 g_113_82 (.ZN (n_113_82), .A (n_112_81), .B (n_113_81), .C1 (n_109_83), .C2 (n_103_86) );
AOI211_X1 g_115_81 (.ZN (n_115_81), .A (n_114_80), .B (n_112_83), .C1 (n_111_82), .C2 (n_105_85) );
AOI211_X1 g_117_80 (.ZN (n_117_80), .A (n_113_82), .B (n_110_82), .C1 (n_113_81), .C2 (n_107_84) );
AOI211_X1 g_119_79 (.ZN (n_119_79), .A (n_115_81), .B (n_112_81), .C1 (n_112_83), .C2 (n_109_83) );
AOI211_X1 g_121_78 (.ZN (n_121_78), .A (n_117_80), .B (n_114_80), .C1 (n_110_82), .C2 (n_111_82) );
AOI211_X1 g_123_77 (.ZN (n_123_77), .A (n_119_79), .B (n_113_82), .C1 (n_112_81), .C2 (n_113_81) );
AOI211_X1 g_125_76 (.ZN (n_125_76), .A (n_121_78), .B (n_115_81), .C1 (n_114_80), .C2 (n_112_83) );
AOI211_X1 g_127_75 (.ZN (n_127_75), .A (n_123_77), .B (n_117_80), .C1 (n_113_82), .C2 (n_110_82) );
AOI211_X1 g_129_76 (.ZN (n_129_76), .A (n_125_76), .B (n_119_79), .C1 (n_115_81), .C2 (n_112_81) );
AOI211_X1 g_127_77 (.ZN (n_127_77), .A (n_127_75), .B (n_121_78), .C1 (n_117_80), .C2 (n_114_80) );
AOI211_X1 g_128_75 (.ZN (n_128_75), .A (n_129_76), .B (n_123_77), .C1 (n_119_79), .C2 (n_113_82) );
AOI211_X1 g_130_76 (.ZN (n_130_76), .A (n_127_77), .B (n_125_76), .C1 (n_121_78), .C2 (n_115_81) );
AOI211_X1 g_132_75 (.ZN (n_132_75), .A (n_128_75), .B (n_127_75), .C1 (n_123_77), .C2 (n_117_80) );
AOI211_X1 g_134_74 (.ZN (n_134_74), .A (n_130_76), .B (n_129_76), .C1 (n_125_76), .C2 (n_119_79) );
AOI211_X1 g_136_73 (.ZN (n_136_73), .A (n_132_75), .B (n_127_77), .C1 (n_127_75), .C2 (n_121_78) );
AOI211_X1 g_135_75 (.ZN (n_135_75), .A (n_134_74), .B (n_128_75), .C1 (n_129_76), .C2 (n_123_77) );
AOI211_X1 g_133_74 (.ZN (n_133_74), .A (n_136_73), .B (n_130_76), .C1 (n_127_77), .C2 (n_125_76) );
AOI211_X1 g_135_73 (.ZN (n_135_73), .A (n_135_75), .B (n_132_75), .C1 (n_128_75), .C2 (n_127_75) );
AOI211_X1 g_137_72 (.ZN (n_137_72), .A (n_133_74), .B (n_134_74), .C1 (n_130_76), .C2 (n_129_76) );
AOI211_X1 g_139_71 (.ZN (n_139_71), .A (n_135_73), .B (n_136_73), .C1 (n_132_75), .C2 (n_127_77) );
AOI211_X1 g_141_70 (.ZN (n_141_70), .A (n_137_72), .B (n_135_75), .C1 (n_134_74), .C2 (n_128_75) );
AOI211_X1 g_143_69 (.ZN (n_143_69), .A (n_139_71), .B (n_133_74), .C1 (n_136_73), .C2 (n_130_76) );
AOI211_X1 g_145_68 (.ZN (n_145_68), .A (n_141_70), .B (n_135_73), .C1 (n_135_75), .C2 (n_132_75) );
AOI211_X1 g_147_69 (.ZN (n_147_69), .A (n_143_69), .B (n_137_72), .C1 (n_133_74), .C2 (n_134_74) );
AOI211_X1 g_145_70 (.ZN (n_145_70), .A (n_145_68), .B (n_139_71), .C1 (n_135_73), .C2 (n_136_73) );
AOI211_X1 g_143_71 (.ZN (n_143_71), .A (n_147_69), .B (n_141_70), .C1 (n_137_72), .C2 (n_135_75) );
AOI211_X1 g_142_69 (.ZN (n_142_69), .A (n_145_70), .B (n_143_69), .C1 (n_139_71), .C2 (n_133_74) );
AOI211_X1 g_140_70 (.ZN (n_140_70), .A (n_143_71), .B (n_145_68), .C1 (n_141_70), .C2 (n_135_73) );
AOI211_X1 g_141_72 (.ZN (n_141_72), .A (n_142_69), .B (n_147_69), .C1 (n_143_69), .C2 (n_137_72) );
AOI211_X1 g_139_73 (.ZN (n_139_73), .A (n_140_70), .B (n_145_70), .C1 (n_145_68), .C2 (n_139_71) );
AOI211_X1 g_137_74 (.ZN (n_137_74), .A (n_141_72), .B (n_143_71), .C1 (n_147_69), .C2 (n_141_70) );
AOI211_X1 g_136_72 (.ZN (n_136_72), .A (n_139_73), .B (n_142_69), .C1 (n_145_70), .C2 (n_143_69) );
AOI211_X1 g_134_73 (.ZN (n_134_73), .A (n_137_74), .B (n_140_70), .C1 (n_143_71), .C2 (n_145_68) );
AOI211_X1 g_132_74 (.ZN (n_132_74), .A (n_136_72), .B (n_141_72), .C1 (n_142_69), .C2 (n_147_69) );
AOI211_X1 g_130_75 (.ZN (n_130_75), .A (n_134_73), .B (n_139_73), .C1 (n_140_70), .C2 (n_145_70) );
AOI211_X1 g_128_76 (.ZN (n_128_76), .A (n_132_74), .B (n_137_74), .C1 (n_141_72), .C2 (n_143_71) );
AOI211_X1 g_126_75 (.ZN (n_126_75), .A (n_130_75), .B (n_136_72), .C1 (n_139_73), .C2 (n_142_69) );
AOI211_X1 g_124_76 (.ZN (n_124_76), .A (n_128_76), .B (n_134_73), .C1 (n_137_74), .C2 (n_140_70) );
AOI211_X1 g_122_77 (.ZN (n_122_77), .A (n_126_75), .B (n_132_74), .C1 (n_136_72), .C2 (n_141_72) );
AOI211_X1 g_120_78 (.ZN (n_120_78), .A (n_124_76), .B (n_130_75), .C1 (n_134_73), .C2 (n_139_73) );
AOI211_X1 g_118_79 (.ZN (n_118_79), .A (n_122_77), .B (n_128_76), .C1 (n_132_74), .C2 (n_137_74) );
AOI211_X1 g_116_80 (.ZN (n_116_80), .A (n_120_78), .B (n_126_75), .C1 (n_130_75), .C2 (n_136_72) );
AOI211_X1 g_114_81 (.ZN (n_114_81), .A (n_118_79), .B (n_124_76), .C1 (n_128_76), .C2 (n_134_73) );
AOI211_X1 g_112_82 (.ZN (n_112_82), .A (n_116_80), .B (n_122_77), .C1 (n_126_75), .C2 (n_132_74) );
AOI211_X1 g_110_83 (.ZN (n_110_83), .A (n_114_81), .B (n_120_78), .C1 (n_124_76), .C2 (n_130_75) );
AOI211_X1 g_108_84 (.ZN (n_108_84), .A (n_112_82), .B (n_118_79), .C1 (n_122_77), .C2 (n_128_76) );
AOI211_X1 g_106_85 (.ZN (n_106_85), .A (n_110_83), .B (n_116_80), .C1 (n_120_78), .C2 (n_126_75) );
AOI211_X1 g_104_86 (.ZN (n_104_86), .A (n_108_84), .B (n_114_81), .C1 (n_118_79), .C2 (n_124_76) );
AOI211_X1 g_102_87 (.ZN (n_102_87), .A (n_106_85), .B (n_112_82), .C1 (n_116_80), .C2 (n_122_77) );
AOI211_X1 g_100_88 (.ZN (n_100_88), .A (n_104_86), .B (n_110_83), .C1 (n_114_81), .C2 (n_120_78) );
AOI211_X1 g_98_89 (.ZN (n_98_89), .A (n_102_87), .B (n_108_84), .C1 (n_112_82), .C2 (n_118_79) );
AOI211_X1 g_96_90 (.ZN (n_96_90), .A (n_100_88), .B (n_106_85), .C1 (n_110_83), .C2 (n_116_80) );
AOI211_X1 g_94_91 (.ZN (n_94_91), .A (n_98_89), .B (n_104_86), .C1 (n_108_84), .C2 (n_114_81) );
AOI211_X1 g_92_90 (.ZN (n_92_90), .A (n_96_90), .B (n_102_87), .C1 (n_106_85), .C2 (n_112_82) );
AOI211_X1 g_90_91 (.ZN (n_90_91), .A (n_94_91), .B (n_100_88), .C1 (n_104_86), .C2 (n_110_83) );
AOI211_X1 g_88_92 (.ZN (n_88_92), .A (n_92_90), .B (n_98_89), .C1 (n_102_87), .C2 (n_108_84) );
AOI211_X1 g_86_93 (.ZN (n_86_93), .A (n_90_91), .B (n_96_90), .C1 (n_100_88), .C2 (n_106_85) );
AOI211_X1 g_84_94 (.ZN (n_84_94), .A (n_88_92), .B (n_94_91), .C1 (n_98_89), .C2 (n_104_86) );
AOI211_X1 g_82_95 (.ZN (n_82_95), .A (n_86_93), .B (n_92_90), .C1 (n_96_90), .C2 (n_102_87) );
AOI211_X1 g_80_96 (.ZN (n_80_96), .A (n_84_94), .B (n_90_91), .C1 (n_94_91), .C2 (n_100_88) );
AOI211_X1 g_81_94 (.ZN (n_81_94), .A (n_82_95), .B (n_88_92), .C1 (n_92_90), .C2 (n_98_89) );
AOI211_X1 g_79_95 (.ZN (n_79_95), .A (n_80_96), .B (n_86_93), .C1 (n_90_91), .C2 (n_96_90) );
AOI211_X1 g_77_96 (.ZN (n_77_96), .A (n_81_94), .B (n_84_94), .C1 (n_88_92), .C2 (n_94_91) );
AOI211_X1 g_75_97 (.ZN (n_75_97), .A (n_79_95), .B (n_82_95), .C1 (n_86_93), .C2 (n_92_90) );
AOI211_X1 g_73_98 (.ZN (n_73_98), .A (n_77_96), .B (n_80_96), .C1 (n_84_94), .C2 (n_90_91) );
AOI211_X1 g_72_100 (.ZN (n_72_100), .A (n_75_97), .B (n_81_94), .C1 (n_82_95), .C2 (n_88_92) );
AOI211_X1 g_74_99 (.ZN (n_74_99), .A (n_73_98), .B (n_79_95), .C1 (n_80_96), .C2 (n_86_93) );
AOI211_X1 g_76_98 (.ZN (n_76_98), .A (n_72_100), .B (n_77_96), .C1 (n_81_94), .C2 (n_84_94) );
AOI211_X1 g_78_97 (.ZN (n_78_97), .A (n_74_99), .B (n_75_97), .C1 (n_79_95), .C2 (n_82_95) );
AOI211_X1 g_77_99 (.ZN (n_77_99), .A (n_76_98), .B (n_73_98), .C1 (n_77_96), .C2 (n_80_96) );
AOI211_X1 g_75_100 (.ZN (n_75_100), .A (n_78_97), .B (n_72_100), .C1 (n_75_97), .C2 (n_81_94) );
AOI211_X1 g_73_101 (.ZN (n_73_101), .A (n_77_99), .B (n_74_99), .C1 (n_73_98), .C2 (n_79_95) );
AOI211_X1 g_71_102 (.ZN (n_71_102), .A (n_75_100), .B (n_76_98), .C1 (n_72_100), .C2 (n_77_96) );
AOI211_X1 g_69_103 (.ZN (n_69_103), .A (n_73_101), .B (n_78_97), .C1 (n_74_99), .C2 (n_75_97) );
AOI211_X1 g_70_101 (.ZN (n_70_101), .A (n_71_102), .B (n_77_99), .C1 (n_76_98), .C2 (n_73_98) );
AOI211_X1 g_68_102 (.ZN (n_68_102), .A (n_69_103), .B (n_75_100), .C1 (n_78_97), .C2 (n_72_100) );
AOI211_X1 g_69_100 (.ZN (n_69_100), .A (n_70_101), .B (n_73_101), .C1 (n_77_99), .C2 (n_74_99) );
AOI211_X1 g_67_101 (.ZN (n_67_101), .A (n_68_102), .B (n_71_102), .C1 (n_75_100), .C2 (n_76_98) );
AOI211_X1 g_65_102 (.ZN (n_65_102), .A (n_69_100), .B (n_69_103), .C1 (n_73_101), .C2 (n_78_97) );
AOI211_X1 g_63_103 (.ZN (n_63_103), .A (n_67_101), .B (n_70_101), .C1 (n_71_102), .C2 (n_77_99) );
AOI211_X1 g_61_104 (.ZN (n_61_104), .A (n_65_102), .B (n_68_102), .C1 (n_69_103), .C2 (n_75_100) );
AOI211_X1 g_59_105 (.ZN (n_59_105), .A (n_63_103), .B (n_69_100), .C1 (n_70_101), .C2 (n_73_101) );
AOI211_X1 g_57_106 (.ZN (n_57_106), .A (n_61_104), .B (n_67_101), .C1 (n_68_102), .C2 (n_71_102) );
AOI211_X1 g_55_107 (.ZN (n_55_107), .A (n_59_105), .B (n_65_102), .C1 (n_69_100), .C2 (n_69_103) );
AOI211_X1 g_53_108 (.ZN (n_53_108), .A (n_57_106), .B (n_63_103), .C1 (n_67_101), .C2 (n_70_101) );
AOI211_X1 g_51_109 (.ZN (n_51_109), .A (n_55_107), .B (n_61_104), .C1 (n_65_102), .C2 (n_68_102) );
AOI211_X1 g_49_110 (.ZN (n_49_110), .A (n_53_108), .B (n_59_105), .C1 (n_63_103), .C2 (n_69_100) );
AOI211_X1 g_47_111 (.ZN (n_47_111), .A (n_51_109), .B (n_57_106), .C1 (n_61_104), .C2 (n_67_101) );
AOI211_X1 g_45_112 (.ZN (n_45_112), .A (n_49_110), .B (n_55_107), .C1 (n_59_105), .C2 (n_65_102) );
AOI211_X1 g_43_113 (.ZN (n_43_113), .A (n_47_111), .B (n_53_108), .C1 (n_57_106), .C2 (n_63_103) );
AOI211_X1 g_41_114 (.ZN (n_41_114), .A (n_45_112), .B (n_51_109), .C1 (n_55_107), .C2 (n_61_104) );
AOI211_X1 g_39_115 (.ZN (n_39_115), .A (n_43_113), .B (n_49_110), .C1 (n_53_108), .C2 (n_59_105) );
AOI211_X1 g_37_116 (.ZN (n_37_116), .A (n_41_114), .B (n_47_111), .C1 (n_51_109), .C2 (n_57_106) );
AOI211_X1 g_35_117 (.ZN (n_35_117), .A (n_39_115), .B (n_45_112), .C1 (n_49_110), .C2 (n_55_107) );
AOI211_X1 g_33_118 (.ZN (n_33_118), .A (n_37_116), .B (n_43_113), .C1 (n_47_111), .C2 (n_53_108) );
AOI211_X1 g_31_119 (.ZN (n_31_119), .A (n_35_117), .B (n_41_114), .C1 (n_45_112), .C2 (n_51_109) );
AOI211_X1 g_29_120 (.ZN (n_29_120), .A (n_33_118), .B (n_39_115), .C1 (n_43_113), .C2 (n_49_110) );
AOI211_X1 g_27_121 (.ZN (n_27_121), .A (n_31_119), .B (n_37_116), .C1 (n_41_114), .C2 (n_47_111) );
AOI211_X1 g_25_122 (.ZN (n_25_122), .A (n_29_120), .B (n_35_117), .C1 (n_39_115), .C2 (n_45_112) );
AOI211_X1 g_23_123 (.ZN (n_23_123), .A (n_27_121), .B (n_33_118), .C1 (n_37_116), .C2 (n_43_113) );
AOI211_X1 g_24_121 (.ZN (n_24_121), .A (n_25_122), .B (n_31_119), .C1 (n_35_117), .C2 (n_41_114) );
AOI211_X1 g_22_122 (.ZN (n_22_122), .A (n_23_123), .B (n_29_120), .C1 (n_33_118), .C2 (n_39_115) );
AOI211_X1 g_21_124 (.ZN (n_21_124), .A (n_24_121), .B (n_27_121), .C1 (n_31_119), .C2 (n_37_116) );
AOI211_X1 g_19_125 (.ZN (n_19_125), .A (n_22_122), .B (n_25_122), .C1 (n_29_120), .C2 (n_35_117) );
AOI211_X1 g_17_126 (.ZN (n_17_126), .A (n_21_124), .B (n_23_123), .C1 (n_27_121), .C2 (n_33_118) );
AOI211_X1 g_15_127 (.ZN (n_15_127), .A (n_19_125), .B (n_24_121), .C1 (n_25_122), .C2 (n_31_119) );
AOI211_X1 g_13_128 (.ZN (n_13_128), .A (n_17_126), .B (n_22_122), .C1 (n_23_123), .C2 (n_29_120) );
AOI211_X1 g_11_129 (.ZN (n_11_129), .A (n_15_127), .B (n_21_124), .C1 (n_24_121), .C2 (n_27_121) );
AOI211_X1 g_12_127 (.ZN (n_12_127), .A (n_13_128), .B (n_19_125), .C1 (n_22_122), .C2 (n_25_122) );
AOI211_X1 g_10_128 (.ZN (n_10_128), .A (n_11_129), .B (n_17_126), .C1 (n_21_124), .C2 (n_23_123) );
AOI211_X1 g_9_130 (.ZN (n_9_130), .A (n_12_127), .B (n_15_127), .C1 (n_19_125), .C2 (n_24_121) );
AOI211_X1 g_8_132 (.ZN (n_8_132), .A (n_10_128), .B (n_13_128), .C1 (n_17_126), .C2 (n_22_122) );
AOI211_X1 g_7_134 (.ZN (n_7_134), .A (n_9_130), .B (n_11_129), .C1 (n_15_127), .C2 (n_21_124) );
AOI211_X1 g_8_136 (.ZN (n_8_136), .A (n_8_132), .B (n_12_127), .C1 (n_13_128), .C2 (n_19_125) );
AOI211_X1 g_9_134 (.ZN (n_9_134), .A (n_7_134), .B (n_10_128), .C1 (n_11_129), .C2 (n_17_126) );
AOI211_X1 g_10_132 (.ZN (n_10_132), .A (n_8_136), .B (n_9_130), .C1 (n_12_127), .C2 (n_15_127) );
AOI211_X1 g_11_130 (.ZN (n_11_130), .A (n_9_134), .B (n_8_132), .C1 (n_10_128), .C2 (n_13_128) );
AOI211_X1 g_13_129 (.ZN (n_13_129), .A (n_10_132), .B (n_7_134), .C1 (n_9_130), .C2 (n_11_129) );
AOI211_X1 g_15_128 (.ZN (n_15_128), .A (n_11_130), .B (n_8_136), .C1 (n_8_132), .C2 (n_12_127) );
AOI211_X1 g_17_127 (.ZN (n_17_127), .A (n_13_129), .B (n_9_134), .C1 (n_7_134), .C2 (n_10_128) );
AOI211_X1 g_16_129 (.ZN (n_16_129), .A (n_15_128), .B (n_10_132), .C1 (n_8_136), .C2 (n_9_130) );
AOI211_X1 g_14_128 (.ZN (n_14_128), .A (n_17_127), .B (n_11_130), .C1 (n_9_134), .C2 (n_8_132) );
AOI211_X1 g_12_129 (.ZN (n_12_129), .A (n_16_129), .B (n_13_129), .C1 (n_10_132), .C2 (n_7_134) );
AOI211_X1 g_14_130 (.ZN (n_14_130), .A (n_14_128), .B (n_15_128), .C1 (n_11_130), .C2 (n_8_136) );
AOI211_X1 g_12_131 (.ZN (n_12_131), .A (n_12_129), .B (n_17_127), .C1 (n_13_129), .C2 (n_9_134) );
AOI211_X1 g_11_133 (.ZN (n_11_133), .A (n_14_130), .B (n_16_129), .C1 (n_15_128), .C2 (n_10_132) );
AOI211_X1 g_10_131 (.ZN (n_10_131), .A (n_12_131), .B (n_14_128), .C1 (n_17_127), .C2 (n_11_130) );
AOI211_X1 g_8_130 (.ZN (n_8_130), .A (n_11_133), .B (n_12_129), .C1 (n_16_129), .C2 (n_13_129) );
AOI211_X1 g_10_129 (.ZN (n_10_129), .A (n_10_131), .B (n_14_130), .C1 (n_14_128), .C2 (n_15_128) );
AOI211_X1 g_9_131 (.ZN (n_9_131), .A (n_8_130), .B (n_12_131), .C1 (n_12_129), .C2 (n_17_127) );
AOI211_X1 g_7_132 (.ZN (n_7_132), .A (n_10_129), .B (n_11_133), .C1 (n_14_130), .C2 (n_16_129) );
AOI211_X1 g_9_133 (.ZN (n_9_133), .A (n_9_131), .B (n_10_131), .C1 (n_12_131), .C2 (n_14_128) );
AOI211_X1 g_8_135 (.ZN (n_8_135), .A (n_7_132), .B (n_8_130), .C1 (n_11_133), .C2 (n_12_129) );
AOI211_X1 g_10_134 (.ZN (n_10_134), .A (n_9_133), .B (n_10_129), .C1 (n_10_131), .C2 (n_14_130) );
AOI211_X1 g_9_132 (.ZN (n_9_132), .A (n_8_135), .B (n_9_131), .C1 (n_8_130), .C2 (n_12_131) );
AOI211_X1 g_11_131 (.ZN (n_11_131), .A (n_10_134), .B (n_7_132), .C1 (n_10_129), .C2 (n_11_133) );
AOI211_X1 g_13_130 (.ZN (n_13_130), .A (n_9_132), .B (n_9_133), .C1 (n_9_131), .C2 (n_10_131) );
AOI211_X1 g_15_129 (.ZN (n_15_129), .A (n_11_131), .B (n_8_135), .C1 (n_7_132), .C2 (n_8_130) );
AOI211_X1 g_16_127 (.ZN (n_16_127), .A (n_13_130), .B (n_10_134), .C1 (n_9_133), .C2 (n_10_129) );
AOI211_X1 g_18_126 (.ZN (n_18_126), .A (n_15_129), .B (n_9_132), .C1 (n_8_135), .C2 (n_9_131) );
AOI211_X1 g_20_125 (.ZN (n_20_125), .A (n_16_127), .B (n_11_131), .C1 (n_10_134), .C2 (n_7_132) );
AOI211_X1 g_22_124 (.ZN (n_22_124), .A (n_18_126), .B (n_13_130), .C1 (n_9_132), .C2 (n_9_133) );
AOI211_X1 g_24_123 (.ZN (n_24_123), .A (n_20_125), .B (n_15_129), .C1 (n_11_131), .C2 (n_8_135) );
AOI211_X1 g_26_122 (.ZN (n_26_122), .A (n_22_124), .B (n_16_127), .C1 (n_13_130), .C2 (n_10_134) );
AOI211_X1 g_28_121 (.ZN (n_28_121), .A (n_24_123), .B (n_18_126), .C1 (n_15_129), .C2 (n_9_132) );
AOI211_X1 g_30_120 (.ZN (n_30_120), .A (n_26_122), .B (n_20_125), .C1 (n_16_127), .C2 (n_11_131) );
AOI211_X1 g_32_119 (.ZN (n_32_119), .A (n_28_121), .B (n_22_124), .C1 (n_18_126), .C2 (n_13_130) );
AOI211_X1 g_34_118 (.ZN (n_34_118), .A (n_30_120), .B (n_24_123), .C1 (n_20_125), .C2 (n_15_129) );
AOI211_X1 g_36_117 (.ZN (n_36_117), .A (n_32_119), .B (n_26_122), .C1 (n_22_124), .C2 (n_16_127) );
AOI211_X1 g_38_116 (.ZN (n_38_116), .A (n_34_118), .B (n_28_121), .C1 (n_24_123), .C2 (n_18_126) );
AOI211_X1 g_40_115 (.ZN (n_40_115), .A (n_36_117), .B (n_30_120), .C1 (n_26_122), .C2 (n_20_125) );
AOI211_X1 g_39_117 (.ZN (n_39_117), .A (n_38_116), .B (n_32_119), .C1 (n_28_121), .C2 (n_22_124) );
AOI211_X1 g_41_116 (.ZN (n_41_116), .A (n_40_115), .B (n_34_118), .C1 (n_30_120), .C2 (n_24_123) );
AOI211_X1 g_43_115 (.ZN (n_43_115), .A (n_39_117), .B (n_36_117), .C1 (n_32_119), .C2 (n_26_122) );
AOI211_X1 g_45_114 (.ZN (n_45_114), .A (n_41_116), .B (n_38_116), .C1 (n_34_118), .C2 (n_28_121) );
AOI211_X1 g_47_113 (.ZN (n_47_113), .A (n_43_115), .B (n_40_115), .C1 (n_36_117), .C2 (n_30_120) );
AOI211_X1 g_49_112 (.ZN (n_49_112), .A (n_45_114), .B (n_39_117), .C1 (n_38_116), .C2 (n_32_119) );
AOI211_X1 g_51_111 (.ZN (n_51_111), .A (n_47_113), .B (n_41_116), .C1 (n_40_115), .C2 (n_34_118) );
AOI211_X1 g_53_110 (.ZN (n_53_110), .A (n_49_112), .B (n_43_115), .C1 (n_39_117), .C2 (n_36_117) );
AOI211_X1 g_55_109 (.ZN (n_55_109), .A (n_51_111), .B (n_45_114), .C1 (n_41_116), .C2 (n_38_116) );
AOI211_X1 g_57_108 (.ZN (n_57_108), .A (n_53_110), .B (n_47_113), .C1 (n_43_115), .C2 (n_40_115) );
AOI211_X1 g_59_107 (.ZN (n_59_107), .A (n_55_109), .B (n_49_112), .C1 (n_45_114), .C2 (n_39_117) );
AOI211_X1 g_61_106 (.ZN (n_61_106), .A (n_57_108), .B (n_51_111), .C1 (n_47_113), .C2 (n_41_116) );
AOI211_X1 g_63_105 (.ZN (n_63_105), .A (n_59_107), .B (n_53_110), .C1 (n_49_112), .C2 (n_43_115) );
AOI211_X1 g_65_104 (.ZN (n_65_104), .A (n_61_106), .B (n_55_109), .C1 (n_51_111), .C2 (n_45_114) );
AOI211_X1 g_67_103 (.ZN (n_67_103), .A (n_63_105), .B (n_57_108), .C1 (n_53_110), .C2 (n_47_113) );
AOI211_X1 g_69_102 (.ZN (n_69_102), .A (n_65_104), .B (n_59_107), .C1 (n_55_109), .C2 (n_49_112) );
AOI211_X1 g_71_101 (.ZN (n_71_101), .A (n_67_103), .B (n_61_106), .C1 (n_57_108), .C2 (n_51_111) );
AOI211_X1 g_73_100 (.ZN (n_73_100), .A (n_69_102), .B (n_63_105), .C1 (n_59_107), .C2 (n_53_110) );
AOI211_X1 g_75_99 (.ZN (n_75_99), .A (n_71_101), .B (n_65_104), .C1 (n_61_106), .C2 (n_55_109) );
AOI211_X1 g_77_98 (.ZN (n_77_98), .A (n_73_100), .B (n_67_103), .C1 (n_63_105), .C2 (n_57_108) );
AOI211_X1 g_78_96 (.ZN (n_78_96), .A (n_75_99), .B (n_69_102), .C1 (n_65_104), .C2 (n_59_107) );
AOI211_X1 g_80_95 (.ZN (n_80_95), .A (n_77_98), .B (n_71_101), .C1 (n_67_103), .C2 (n_61_106) );
AOI211_X1 g_82_94 (.ZN (n_82_94), .A (n_78_96), .B (n_73_100), .C1 (n_69_102), .C2 (n_63_105) );
AOI211_X1 g_81_96 (.ZN (n_81_96), .A (n_80_95), .B (n_75_99), .C1 (n_71_101), .C2 (n_65_104) );
AOI211_X1 g_79_97 (.ZN (n_79_97), .A (n_82_94), .B (n_77_98), .C1 (n_73_100), .C2 (n_67_103) );
AOI211_X1 g_78_99 (.ZN (n_78_99), .A (n_81_96), .B (n_78_96), .C1 (n_75_99), .C2 (n_69_102) );
AOI211_X1 g_76_100 (.ZN (n_76_100), .A (n_79_97), .B (n_80_95), .C1 (n_77_98), .C2 (n_71_101) );
AOI211_X1 g_74_101 (.ZN (n_74_101), .A (n_78_99), .B (n_82_94), .C1 (n_78_96), .C2 (n_73_100) );
AOI211_X1 g_72_102 (.ZN (n_72_102), .A (n_76_100), .B (n_81_96), .C1 (n_80_95), .C2 (n_75_99) );
AOI211_X1 g_70_103 (.ZN (n_70_103), .A (n_74_101), .B (n_79_97), .C1 (n_82_94), .C2 (n_77_98) );
AOI211_X1 g_68_104 (.ZN (n_68_104), .A (n_72_102), .B (n_78_99), .C1 (n_81_96), .C2 (n_78_96) );
AOI211_X1 g_66_103 (.ZN (n_66_103), .A (n_70_103), .B (n_76_100), .C1 (n_79_97), .C2 (n_80_95) );
AOI211_X1 g_64_104 (.ZN (n_64_104), .A (n_68_104), .B (n_74_101), .C1 (n_78_99), .C2 (n_82_94) );
AOI211_X1 g_62_105 (.ZN (n_62_105), .A (n_66_103), .B (n_72_102), .C1 (n_76_100), .C2 (n_81_96) );
AOI211_X1 g_60_106 (.ZN (n_60_106), .A (n_64_104), .B (n_70_103), .C1 (n_74_101), .C2 (n_79_97) );
AOI211_X1 g_58_107 (.ZN (n_58_107), .A (n_62_105), .B (n_68_104), .C1 (n_72_102), .C2 (n_78_99) );
AOI211_X1 g_56_108 (.ZN (n_56_108), .A (n_60_106), .B (n_66_103), .C1 (n_70_103), .C2 (n_76_100) );
AOI211_X1 g_54_109 (.ZN (n_54_109), .A (n_58_107), .B (n_64_104), .C1 (n_68_104), .C2 (n_74_101) );
AOI211_X1 g_52_110 (.ZN (n_52_110), .A (n_56_108), .B (n_62_105), .C1 (n_66_103), .C2 (n_72_102) );
AOI211_X1 g_50_111 (.ZN (n_50_111), .A (n_54_109), .B (n_60_106), .C1 (n_64_104), .C2 (n_70_103) );
AOI211_X1 g_48_112 (.ZN (n_48_112), .A (n_52_110), .B (n_58_107), .C1 (n_62_105), .C2 (n_68_104) );
AOI211_X1 g_46_113 (.ZN (n_46_113), .A (n_50_111), .B (n_56_108), .C1 (n_60_106), .C2 (n_66_103) );
AOI211_X1 g_44_114 (.ZN (n_44_114), .A (n_48_112), .B (n_54_109), .C1 (n_58_107), .C2 (n_64_104) );
AOI211_X1 g_42_115 (.ZN (n_42_115), .A (n_46_113), .B (n_52_110), .C1 (n_56_108), .C2 (n_62_105) );
AOI211_X1 g_40_116 (.ZN (n_40_116), .A (n_44_114), .B (n_50_111), .C1 (n_54_109), .C2 (n_60_106) );
AOI211_X1 g_38_117 (.ZN (n_38_117), .A (n_42_115), .B (n_48_112), .C1 (n_52_110), .C2 (n_58_107) );
AOI211_X1 g_36_118 (.ZN (n_36_118), .A (n_40_116), .B (n_46_113), .C1 (n_50_111), .C2 (n_56_108) );
AOI211_X1 g_34_119 (.ZN (n_34_119), .A (n_38_117), .B (n_44_114), .C1 (n_48_112), .C2 (n_54_109) );
AOI211_X1 g_32_120 (.ZN (n_32_120), .A (n_36_118), .B (n_42_115), .C1 (n_46_113), .C2 (n_52_110) );
AOI211_X1 g_30_121 (.ZN (n_30_121), .A (n_34_119), .B (n_40_116), .C1 (n_44_114), .C2 (n_50_111) );
AOI211_X1 g_28_122 (.ZN (n_28_122), .A (n_32_120), .B (n_38_117), .C1 (n_42_115), .C2 (n_48_112) );
AOI211_X1 g_26_123 (.ZN (n_26_123), .A (n_30_121), .B (n_36_118), .C1 (n_40_116), .C2 (n_46_113) );
AOI211_X1 g_24_124 (.ZN (n_24_124), .A (n_28_122), .B (n_34_119), .C1 (n_38_117), .C2 (n_44_114) );
AOI211_X1 g_22_125 (.ZN (n_22_125), .A (n_26_123), .B (n_32_120), .C1 (n_36_118), .C2 (n_42_115) );
AOI211_X1 g_20_126 (.ZN (n_20_126), .A (n_24_124), .B (n_30_121), .C1 (n_34_119), .C2 (n_40_116) );
AOI211_X1 g_18_127 (.ZN (n_18_127), .A (n_22_125), .B (n_28_122), .C1 (n_32_120), .C2 (n_38_117) );
AOI211_X1 g_16_128 (.ZN (n_16_128), .A (n_20_126), .B (n_26_123), .C1 (n_30_121), .C2 (n_36_118) );
AOI211_X1 g_14_129 (.ZN (n_14_129), .A (n_18_127), .B (n_24_124), .C1 (n_28_122), .C2 (n_34_119) );
AOI211_X1 g_12_130 (.ZN (n_12_130), .A (n_16_128), .B (n_22_125), .C1 (n_26_123), .C2 (n_32_120) );
AOI211_X1 g_11_132 (.ZN (n_11_132), .A (n_14_129), .B (n_20_126), .C1 (n_24_124), .C2 (n_30_121) );
AOI211_X1 g_13_131 (.ZN (n_13_131), .A (n_12_130), .B (n_18_127), .C1 (n_22_125), .C2 (n_28_122) );
AOI211_X1 g_15_130 (.ZN (n_15_130), .A (n_11_132), .B (n_16_128), .C1 (n_20_126), .C2 (n_26_123) );
AOI211_X1 g_17_129 (.ZN (n_17_129), .A (n_13_131), .B (n_14_129), .C1 (n_18_127), .C2 (n_24_124) );
AOI211_X1 g_19_128 (.ZN (n_19_128), .A (n_15_130), .B (n_12_130), .C1 (n_16_128), .C2 (n_22_125) );
AOI211_X1 g_21_127 (.ZN (n_21_127), .A (n_17_129), .B (n_11_132), .C1 (n_14_129), .C2 (n_20_126) );
AOI211_X1 g_23_126 (.ZN (n_23_126), .A (n_19_128), .B (n_13_131), .C1 (n_12_130), .C2 (n_18_127) );
AOI211_X1 g_25_125 (.ZN (n_25_125), .A (n_21_127), .B (n_15_130), .C1 (n_11_132), .C2 (n_16_128) );
AOI211_X1 g_27_124 (.ZN (n_27_124), .A (n_23_126), .B (n_17_129), .C1 (n_13_131), .C2 (n_14_129) );
AOI211_X1 g_25_123 (.ZN (n_25_123), .A (n_25_125), .B (n_19_128), .C1 (n_15_130), .C2 (n_12_130) );
AOI211_X1 g_24_125 (.ZN (n_24_125), .A (n_27_124), .B (n_21_127), .C1 (n_17_129), .C2 (n_11_132) );
AOI211_X1 g_26_124 (.ZN (n_26_124), .A (n_25_123), .B (n_23_126), .C1 (n_19_128), .C2 (n_13_131) );
AOI211_X1 g_28_123 (.ZN (n_28_123), .A (n_24_125), .B (n_25_125), .C1 (n_21_127), .C2 (n_15_130) );
AOI211_X1 g_30_122 (.ZN (n_30_122), .A (n_26_124), .B (n_27_124), .C1 (n_23_126), .C2 (n_17_129) );
AOI211_X1 g_32_121 (.ZN (n_32_121), .A (n_28_123), .B (n_25_123), .C1 (n_25_125), .C2 (n_19_128) );
AOI211_X1 g_33_119 (.ZN (n_33_119), .A (n_30_122), .B (n_24_125), .C1 (n_27_124), .C2 (n_21_127) );
AOI211_X1 g_35_118 (.ZN (n_35_118), .A (n_32_121), .B (n_26_124), .C1 (n_25_123), .C2 (n_23_126) );
AOI211_X1 g_37_117 (.ZN (n_37_117), .A (n_33_119), .B (n_28_123), .C1 (n_24_125), .C2 (n_25_125) );
AOI211_X1 g_39_116 (.ZN (n_39_116), .A (n_35_118), .B (n_30_122), .C1 (n_26_124), .C2 (n_27_124) );
AOI211_X1 g_41_115 (.ZN (n_41_115), .A (n_37_117), .B (n_32_121), .C1 (n_28_123), .C2 (n_25_123) );
AOI211_X1 g_43_114 (.ZN (n_43_114), .A (n_39_116), .B (n_33_119), .C1 (n_30_122), .C2 (n_24_125) );
AOI211_X1 g_45_113 (.ZN (n_45_113), .A (n_41_115), .B (n_35_118), .C1 (n_32_121), .C2 (n_26_124) );
AOI211_X1 g_47_112 (.ZN (n_47_112), .A (n_43_114), .B (n_37_117), .C1 (n_33_119), .C2 (n_28_123) );
AOI211_X1 g_49_111 (.ZN (n_49_111), .A (n_45_113), .B (n_39_116), .C1 (n_35_118), .C2 (n_30_122) );
AOI211_X1 g_51_110 (.ZN (n_51_110), .A (n_47_112), .B (n_41_115), .C1 (n_37_117), .C2 (n_32_121) );
AOI211_X1 g_53_109 (.ZN (n_53_109), .A (n_49_111), .B (n_43_114), .C1 (n_39_116), .C2 (n_33_119) );
AOI211_X1 g_55_108 (.ZN (n_55_108), .A (n_51_110), .B (n_45_113), .C1 (n_41_115), .C2 (n_35_118) );
AOI211_X1 g_57_107 (.ZN (n_57_107), .A (n_53_109), .B (n_47_112), .C1 (n_43_114), .C2 (n_37_117) );
AOI211_X1 g_59_106 (.ZN (n_59_106), .A (n_55_108), .B (n_49_111), .C1 (n_45_113), .C2 (n_39_116) );
AOI211_X1 g_61_105 (.ZN (n_61_105), .A (n_57_107), .B (n_51_110), .C1 (n_47_112), .C2 (n_41_115) );
AOI211_X1 g_63_104 (.ZN (n_63_104), .A (n_59_106), .B (n_53_109), .C1 (n_49_111), .C2 (n_43_114) );
AOI211_X1 g_65_103 (.ZN (n_65_103), .A (n_61_105), .B (n_55_108), .C1 (n_51_110), .C2 (n_45_113) );
AOI211_X1 g_66_105 (.ZN (n_66_105), .A (n_63_104), .B (n_57_107), .C1 (n_53_109), .C2 (n_47_112) );
AOI211_X1 g_64_106 (.ZN (n_64_106), .A (n_65_103), .B (n_59_106), .C1 (n_55_108), .C2 (n_49_111) );
AOI211_X1 g_62_107 (.ZN (n_62_107), .A (n_66_105), .B (n_61_105), .C1 (n_57_107), .C2 (n_51_110) );
AOI211_X1 g_60_108 (.ZN (n_60_108), .A (n_64_106), .B (n_63_104), .C1 (n_59_106), .C2 (n_53_109) );
AOI211_X1 g_58_109 (.ZN (n_58_109), .A (n_62_107), .B (n_65_103), .C1 (n_61_105), .C2 (n_55_108) );
AOI211_X1 g_56_110 (.ZN (n_56_110), .A (n_60_108), .B (n_66_105), .C1 (n_63_104), .C2 (n_57_107) );
AOI211_X1 g_54_111 (.ZN (n_54_111), .A (n_58_109), .B (n_64_106), .C1 (n_65_103), .C2 (n_59_106) );
AOI211_X1 g_52_112 (.ZN (n_52_112), .A (n_56_110), .B (n_62_107), .C1 (n_66_105), .C2 (n_61_105) );
AOI211_X1 g_50_113 (.ZN (n_50_113), .A (n_54_111), .B (n_60_108), .C1 (n_64_106), .C2 (n_63_104) );
AOI211_X1 g_48_114 (.ZN (n_48_114), .A (n_52_112), .B (n_58_109), .C1 (n_62_107), .C2 (n_65_103) );
AOI211_X1 g_46_115 (.ZN (n_46_115), .A (n_50_113), .B (n_56_110), .C1 (n_60_108), .C2 (n_66_105) );
AOI211_X1 g_44_116 (.ZN (n_44_116), .A (n_48_114), .B (n_54_111), .C1 (n_58_109), .C2 (n_64_106) );
AOI211_X1 g_42_117 (.ZN (n_42_117), .A (n_46_115), .B (n_52_112), .C1 (n_56_110), .C2 (n_62_107) );
AOI211_X1 g_40_118 (.ZN (n_40_118), .A (n_44_116), .B (n_50_113), .C1 (n_54_111), .C2 (n_60_108) );
AOI211_X1 g_38_119 (.ZN (n_38_119), .A (n_42_117), .B (n_48_114), .C1 (n_52_112), .C2 (n_58_109) );
AOI211_X1 g_36_120 (.ZN (n_36_120), .A (n_40_118), .B (n_46_115), .C1 (n_50_113), .C2 (n_56_110) );
AOI211_X1 g_37_118 (.ZN (n_37_118), .A (n_38_119), .B (n_44_116), .C1 (n_48_114), .C2 (n_54_111) );
AOI211_X1 g_35_119 (.ZN (n_35_119), .A (n_36_120), .B (n_42_117), .C1 (n_46_115), .C2 (n_52_112) );
AOI211_X1 g_33_120 (.ZN (n_33_120), .A (n_37_118), .B (n_40_118), .C1 (n_44_116), .C2 (n_50_113) );
AOI211_X1 g_31_121 (.ZN (n_31_121), .A (n_35_119), .B (n_38_119), .C1 (n_42_117), .C2 (n_48_114) );
AOI211_X1 g_29_122 (.ZN (n_29_122), .A (n_33_120), .B (n_36_120), .C1 (n_40_118), .C2 (n_46_115) );
AOI211_X1 g_27_123 (.ZN (n_27_123), .A (n_31_121), .B (n_37_118), .C1 (n_38_119), .C2 (n_44_116) );
AOI211_X1 g_25_124 (.ZN (n_25_124), .A (n_29_122), .B (n_35_119), .C1 (n_36_120), .C2 (n_42_117) );
AOI211_X1 g_23_125 (.ZN (n_23_125), .A (n_27_123), .B (n_33_120), .C1 (n_37_118), .C2 (n_40_118) );
AOI211_X1 g_21_126 (.ZN (n_21_126), .A (n_25_124), .B (n_31_121), .C1 (n_35_119), .C2 (n_38_119) );
AOI211_X1 g_19_127 (.ZN (n_19_127), .A (n_23_125), .B (n_29_122), .C1 (n_33_120), .C2 (n_36_120) );
AOI211_X1 g_17_128 (.ZN (n_17_128), .A (n_21_126), .B (n_27_123), .C1 (n_31_121), .C2 (n_37_118) );
AOI211_X1 g_16_130 (.ZN (n_16_130), .A (n_19_127), .B (n_25_124), .C1 (n_29_122), .C2 (n_35_119) );
AOI211_X1 g_18_129 (.ZN (n_18_129), .A (n_17_128), .B (n_23_125), .C1 (n_27_123), .C2 (n_33_120) );
AOI211_X1 g_20_128 (.ZN (n_20_128), .A (n_16_130), .B (n_21_126), .C1 (n_25_124), .C2 (n_31_121) );
AOI211_X1 g_22_127 (.ZN (n_22_127), .A (n_18_129), .B (n_19_127), .C1 (n_23_125), .C2 (n_29_122) );
AOI211_X1 g_24_126 (.ZN (n_24_126), .A (n_20_128), .B (n_17_128), .C1 (n_21_126), .C2 (n_27_123) );
AOI211_X1 g_26_125 (.ZN (n_26_125), .A (n_22_127), .B (n_16_130), .C1 (n_19_127), .C2 (n_25_124) );
AOI211_X1 g_28_124 (.ZN (n_28_124), .A (n_24_126), .B (n_18_129), .C1 (n_17_128), .C2 (n_23_125) );
AOI211_X1 g_30_123 (.ZN (n_30_123), .A (n_26_125), .B (n_20_128), .C1 (n_16_130), .C2 (n_21_126) );
AOI211_X1 g_32_122 (.ZN (n_32_122), .A (n_28_124), .B (n_22_127), .C1 (n_18_129), .C2 (n_19_127) );
AOI211_X1 g_34_121 (.ZN (n_34_121), .A (n_30_123), .B (n_24_126), .C1 (n_20_128), .C2 (n_17_128) );
AOI211_X1 g_33_123 (.ZN (n_33_123), .A (n_32_122), .B (n_26_125), .C1 (n_22_127), .C2 (n_16_130) );
AOI211_X1 g_31_122 (.ZN (n_31_122), .A (n_34_121), .B (n_28_124), .C1 (n_24_126), .C2 (n_18_129) );
AOI211_X1 g_29_123 (.ZN (n_29_123), .A (n_33_123), .B (n_30_123), .C1 (n_26_125), .C2 (n_20_128) );
AOI211_X1 g_31_124 (.ZN (n_31_124), .A (n_31_122), .B (n_32_122), .C1 (n_28_124), .C2 (n_22_127) );
AOI211_X1 g_29_125 (.ZN (n_29_125), .A (n_29_123), .B (n_34_121), .C1 (n_30_123), .C2 (n_24_126) );
AOI211_X1 g_27_126 (.ZN (n_27_126), .A (n_31_124), .B (n_33_123), .C1 (n_32_122), .C2 (n_26_125) );
AOI211_X1 g_25_127 (.ZN (n_25_127), .A (n_29_125), .B (n_31_122), .C1 (n_34_121), .C2 (n_28_124) );
AOI211_X1 g_23_128 (.ZN (n_23_128), .A (n_27_126), .B (n_29_123), .C1 (n_33_123), .C2 (n_30_123) );
AOI211_X1 g_22_126 (.ZN (n_22_126), .A (n_25_127), .B (n_31_124), .C1 (n_31_122), .C2 (n_32_122) );
AOI211_X1 g_20_127 (.ZN (n_20_127), .A (n_23_128), .B (n_29_125), .C1 (n_29_123), .C2 (n_34_121) );
AOI211_X1 g_18_128 (.ZN (n_18_128), .A (n_22_126), .B (n_27_126), .C1 (n_31_124), .C2 (n_33_123) );
AOI211_X1 g_17_130 (.ZN (n_17_130), .A (n_20_127), .B (n_25_127), .C1 (n_29_125), .C2 (n_31_122) );
AOI211_X1 g_19_129 (.ZN (n_19_129), .A (n_18_128), .B (n_23_128), .C1 (n_27_126), .C2 (n_29_123) );
AOI211_X1 g_21_128 (.ZN (n_21_128), .A (n_17_130), .B (n_22_126), .C1 (n_25_127), .C2 (n_31_124) );
AOI211_X1 g_23_127 (.ZN (n_23_127), .A (n_19_129), .B (n_20_127), .C1 (n_23_128), .C2 (n_29_125) );
AOI211_X1 g_25_126 (.ZN (n_25_126), .A (n_21_128), .B (n_18_128), .C1 (n_22_126), .C2 (n_27_126) );
AOI211_X1 g_27_125 (.ZN (n_27_125), .A (n_23_127), .B (n_17_130), .C1 (n_20_127), .C2 (n_25_127) );
AOI211_X1 g_29_124 (.ZN (n_29_124), .A (n_25_126), .B (n_19_129), .C1 (n_18_128), .C2 (n_23_128) );
AOI211_X1 g_31_123 (.ZN (n_31_123), .A (n_27_125), .B (n_21_128), .C1 (n_17_130), .C2 (n_22_126) );
AOI211_X1 g_33_122 (.ZN (n_33_122), .A (n_29_124), .B (n_23_127), .C1 (n_19_129), .C2 (n_20_127) );
AOI211_X1 g_34_120 (.ZN (n_34_120), .A (n_31_123), .B (n_25_126), .C1 (n_21_128), .C2 (n_18_128) );
AOI211_X1 g_36_119 (.ZN (n_36_119), .A (n_33_122), .B (n_27_125), .C1 (n_23_127), .C2 (n_17_130) );
AOI211_X1 g_38_118 (.ZN (n_38_118), .A (n_34_120), .B (n_29_124), .C1 (n_25_126), .C2 (n_19_129) );
AOI211_X1 g_40_117 (.ZN (n_40_117), .A (n_36_119), .B (n_31_123), .C1 (n_27_125), .C2 (n_21_128) );
AOI211_X1 g_42_116 (.ZN (n_42_116), .A (n_38_118), .B (n_33_122), .C1 (n_29_124), .C2 (n_23_127) );
AOI211_X1 g_44_115 (.ZN (n_44_115), .A (n_40_117), .B (n_34_120), .C1 (n_31_123), .C2 (n_25_126) );
AOI211_X1 g_46_114 (.ZN (n_46_114), .A (n_42_116), .B (n_36_119), .C1 (n_33_122), .C2 (n_27_125) );
AOI211_X1 g_48_113 (.ZN (n_48_113), .A (n_44_115), .B (n_38_118), .C1 (n_34_120), .C2 (n_29_124) );
AOI211_X1 g_50_112 (.ZN (n_50_112), .A (n_46_114), .B (n_40_117), .C1 (n_36_119), .C2 (n_31_123) );
AOI211_X1 g_52_111 (.ZN (n_52_111), .A (n_48_113), .B (n_42_116), .C1 (n_38_118), .C2 (n_33_122) );
AOI211_X1 g_54_110 (.ZN (n_54_110), .A (n_50_112), .B (n_44_115), .C1 (n_40_117), .C2 (n_34_120) );
AOI211_X1 g_56_109 (.ZN (n_56_109), .A (n_52_111), .B (n_46_114), .C1 (n_42_116), .C2 (n_36_119) );
AOI211_X1 g_58_108 (.ZN (n_58_108), .A (n_54_110), .B (n_48_113), .C1 (n_44_115), .C2 (n_38_118) );
AOI211_X1 g_60_107 (.ZN (n_60_107), .A (n_56_109), .B (n_50_112), .C1 (n_46_114), .C2 (n_40_117) );
AOI211_X1 g_62_106 (.ZN (n_62_106), .A (n_58_108), .B (n_52_111), .C1 (n_48_113), .C2 (n_42_116) );
AOI211_X1 g_64_105 (.ZN (n_64_105), .A (n_60_107), .B (n_54_110), .C1 (n_50_112), .C2 (n_44_115) );
AOI211_X1 g_66_104 (.ZN (n_66_104), .A (n_62_106), .B (n_56_109), .C1 (n_52_111), .C2 (n_46_114) );
AOI211_X1 g_68_103 (.ZN (n_68_103), .A (n_64_105), .B (n_58_108), .C1 (n_54_110), .C2 (n_48_113) );
AOI211_X1 g_70_102 (.ZN (n_70_102), .A (n_66_104), .B (n_60_107), .C1 (n_56_109), .C2 (n_50_112) );
AOI211_X1 g_72_101 (.ZN (n_72_101), .A (n_68_103), .B (n_62_106), .C1 (n_58_108), .C2 (n_52_111) );
AOI211_X1 g_74_100 (.ZN (n_74_100), .A (n_70_102), .B (n_64_105), .C1 (n_60_107), .C2 (n_54_110) );
AOI211_X1 g_76_99 (.ZN (n_76_99), .A (n_72_101), .B (n_66_104), .C1 (n_62_106), .C2 (n_56_109) );
AOI211_X1 g_78_98 (.ZN (n_78_98), .A (n_74_100), .B (n_68_103), .C1 (n_64_105), .C2 (n_58_108) );
AOI211_X1 g_79_96 (.ZN (n_79_96), .A (n_76_99), .B (n_70_102), .C1 (n_66_104), .C2 (n_60_107) );
AOI211_X1 g_81_95 (.ZN (n_81_95), .A (n_78_98), .B (n_72_101), .C1 (n_68_103), .C2 (n_62_106) );
AOI211_X1 g_83_94 (.ZN (n_83_94), .A (n_79_96), .B (n_74_100), .C1 (n_70_102), .C2 (n_64_105) );
AOI211_X1 g_85_93 (.ZN (n_85_93), .A (n_81_95), .B (n_76_99), .C1 (n_72_101), .C2 (n_66_104) );
AOI211_X1 g_87_92 (.ZN (n_87_92), .A (n_83_94), .B (n_78_98), .C1 (n_74_100), .C2 (n_68_103) );
AOI211_X1 g_89_91 (.ZN (n_89_91), .A (n_85_93), .B (n_79_96), .C1 (n_76_99), .C2 (n_70_102) );
AOI211_X1 g_91_90 (.ZN (n_91_90), .A (n_87_92), .B (n_81_95), .C1 (n_78_98), .C2 (n_72_101) );
AOI211_X1 g_92_92 (.ZN (n_92_92), .A (n_89_91), .B (n_83_94), .C1 (n_79_96), .C2 (n_74_100) );
AOI211_X1 g_90_93 (.ZN (n_90_93), .A (n_91_90), .B (n_85_93), .C1 (n_81_95), .C2 (n_76_99) );
AOI211_X1 g_91_91 (.ZN (n_91_91), .A (n_92_92), .B (n_87_92), .C1 (n_83_94), .C2 (n_78_98) );
AOI211_X1 g_89_92 (.ZN (n_89_92), .A (n_90_93), .B (n_89_91), .C1 (n_85_93), .C2 (n_79_96) );
AOI211_X1 g_87_93 (.ZN (n_87_93), .A (n_91_91), .B (n_91_90), .C1 (n_87_92), .C2 (n_81_95) );
AOI211_X1 g_85_94 (.ZN (n_85_94), .A (n_89_92), .B (n_92_92), .C1 (n_89_91), .C2 (n_83_94) );
AOI211_X1 g_83_95 (.ZN (n_83_95), .A (n_87_93), .B (n_90_93), .C1 (n_91_90), .C2 (n_85_93) );
AOI211_X1 g_82_97 (.ZN (n_82_97), .A (n_85_94), .B (n_91_91), .C1 (n_92_92), .C2 (n_87_92) );
AOI211_X1 g_80_98 (.ZN (n_80_98), .A (n_83_95), .B (n_89_92), .C1 (n_90_93), .C2 (n_89_91) );
AOI211_X1 g_79_100 (.ZN (n_79_100), .A (n_82_97), .B (n_87_93), .C1 (n_91_91), .C2 (n_91_90) );
AOI211_X1 g_77_101 (.ZN (n_77_101), .A (n_80_98), .B (n_85_94), .C1 (n_89_92), .C2 (n_92_92) );
AOI211_X1 g_75_102 (.ZN (n_75_102), .A (n_79_100), .B (n_83_95), .C1 (n_87_93), .C2 (n_90_93) );
AOI211_X1 g_73_103 (.ZN (n_73_103), .A (n_77_101), .B (n_82_97), .C1 (n_85_94), .C2 (n_91_91) );
AOI211_X1 g_71_104 (.ZN (n_71_104), .A (n_75_102), .B (n_80_98), .C1 (n_83_95), .C2 (n_89_92) );
AOI211_X1 g_69_105 (.ZN (n_69_105), .A (n_73_103), .B (n_79_100), .C1 (n_82_97), .C2 (n_87_93) );
AOI211_X1 g_67_104 (.ZN (n_67_104), .A (n_71_104), .B (n_77_101), .C1 (n_80_98), .C2 (n_85_94) );
AOI211_X1 g_65_105 (.ZN (n_65_105), .A (n_69_105), .B (n_75_102), .C1 (n_79_100), .C2 (n_83_95) );
AOI211_X1 g_63_106 (.ZN (n_63_106), .A (n_67_104), .B (n_73_103), .C1 (n_77_101), .C2 (n_82_97) );
AOI211_X1 g_61_107 (.ZN (n_61_107), .A (n_65_105), .B (n_71_104), .C1 (n_75_102), .C2 (n_80_98) );
AOI211_X1 g_59_108 (.ZN (n_59_108), .A (n_63_106), .B (n_69_105), .C1 (n_73_103), .C2 (n_79_100) );
AOI211_X1 g_57_109 (.ZN (n_57_109), .A (n_61_107), .B (n_67_104), .C1 (n_71_104), .C2 (n_77_101) );
AOI211_X1 g_55_110 (.ZN (n_55_110), .A (n_59_108), .B (n_65_105), .C1 (n_69_105), .C2 (n_75_102) );
AOI211_X1 g_53_111 (.ZN (n_53_111), .A (n_57_109), .B (n_63_106), .C1 (n_67_104), .C2 (n_73_103) );
AOI211_X1 g_51_112 (.ZN (n_51_112), .A (n_55_110), .B (n_61_107), .C1 (n_65_105), .C2 (n_71_104) );
AOI211_X1 g_49_113 (.ZN (n_49_113), .A (n_53_111), .B (n_59_108), .C1 (n_63_106), .C2 (n_69_105) );
AOI211_X1 g_47_114 (.ZN (n_47_114), .A (n_51_112), .B (n_57_109), .C1 (n_61_107), .C2 (n_67_104) );
AOI211_X1 g_45_115 (.ZN (n_45_115), .A (n_49_113), .B (n_55_110), .C1 (n_59_108), .C2 (n_65_105) );
AOI211_X1 g_43_116 (.ZN (n_43_116), .A (n_47_114), .B (n_53_111), .C1 (n_57_109), .C2 (n_63_106) );
AOI211_X1 g_41_117 (.ZN (n_41_117), .A (n_45_115), .B (n_51_112), .C1 (n_55_110), .C2 (n_61_107) );
AOI211_X1 g_39_118 (.ZN (n_39_118), .A (n_43_116), .B (n_49_113), .C1 (n_53_111), .C2 (n_59_108) );
AOI211_X1 g_37_119 (.ZN (n_37_119), .A (n_41_117), .B (n_47_114), .C1 (n_51_112), .C2 (n_57_109) );
AOI211_X1 g_35_120 (.ZN (n_35_120), .A (n_39_118), .B (n_45_115), .C1 (n_49_113), .C2 (n_55_110) );
AOI211_X1 g_33_121 (.ZN (n_33_121), .A (n_37_119), .B (n_43_116), .C1 (n_47_114), .C2 (n_53_111) );
AOI211_X1 g_35_122 (.ZN (n_35_122), .A (n_35_120), .B (n_41_117), .C1 (n_45_115), .C2 (n_51_112) );
AOI211_X1 g_37_121 (.ZN (n_37_121), .A (n_33_121), .B (n_39_118), .C1 (n_43_116), .C2 (n_49_113) );
AOI211_X1 g_39_120 (.ZN (n_39_120), .A (n_35_122), .B (n_37_119), .C1 (n_41_117), .C2 (n_47_114) );
AOI211_X1 g_41_119 (.ZN (n_41_119), .A (n_37_121), .B (n_35_120), .C1 (n_39_118), .C2 (n_45_115) );
AOI211_X1 g_43_118 (.ZN (n_43_118), .A (n_39_120), .B (n_33_121), .C1 (n_37_119), .C2 (n_43_116) );
AOI211_X1 g_45_117 (.ZN (n_45_117), .A (n_41_119), .B (n_35_122), .C1 (n_35_120), .C2 (n_41_117) );
AOI211_X1 g_47_116 (.ZN (n_47_116), .A (n_43_118), .B (n_37_121), .C1 (n_33_121), .C2 (n_39_118) );
AOI211_X1 g_49_115 (.ZN (n_49_115), .A (n_45_117), .B (n_39_120), .C1 (n_35_122), .C2 (n_37_119) );
AOI211_X1 g_51_114 (.ZN (n_51_114), .A (n_47_116), .B (n_41_119), .C1 (n_37_121), .C2 (n_35_120) );
AOI211_X1 g_53_113 (.ZN (n_53_113), .A (n_49_115), .B (n_43_118), .C1 (n_39_120), .C2 (n_33_121) );
AOI211_X1 g_55_112 (.ZN (n_55_112), .A (n_51_114), .B (n_45_117), .C1 (n_41_119), .C2 (n_35_122) );
AOI211_X1 g_57_111 (.ZN (n_57_111), .A (n_53_113), .B (n_47_116), .C1 (n_43_118), .C2 (n_37_121) );
AOI211_X1 g_59_110 (.ZN (n_59_110), .A (n_55_112), .B (n_49_115), .C1 (n_45_117), .C2 (n_39_120) );
AOI211_X1 g_61_109 (.ZN (n_61_109), .A (n_57_111), .B (n_51_114), .C1 (n_47_116), .C2 (n_41_119) );
AOI211_X1 g_63_108 (.ZN (n_63_108), .A (n_59_110), .B (n_53_113), .C1 (n_49_115), .C2 (n_43_118) );
AOI211_X1 g_65_107 (.ZN (n_65_107), .A (n_61_109), .B (n_55_112), .C1 (n_51_114), .C2 (n_45_117) );
AOI211_X1 g_67_106 (.ZN (n_67_106), .A (n_63_108), .B (n_57_111), .C1 (n_53_113), .C2 (n_47_116) );
AOI211_X1 g_66_108 (.ZN (n_66_108), .A (n_65_107), .B (n_59_110), .C1 (n_55_112), .C2 (n_49_115) );
AOI211_X1 g_65_106 (.ZN (n_65_106), .A (n_67_106), .B (n_61_109), .C1 (n_57_111), .C2 (n_51_114) );
AOI211_X1 g_67_105 (.ZN (n_67_105), .A (n_66_108), .B (n_63_108), .C1 (n_59_110), .C2 (n_53_113) );
AOI211_X1 g_69_104 (.ZN (n_69_104), .A (n_65_106), .B (n_65_107), .C1 (n_61_109), .C2 (n_55_112) );
AOI211_X1 g_71_103 (.ZN (n_71_103), .A (n_67_105), .B (n_67_106), .C1 (n_63_108), .C2 (n_57_111) );
AOI211_X1 g_73_102 (.ZN (n_73_102), .A (n_69_104), .B (n_66_108), .C1 (n_65_107), .C2 (n_59_110) );
AOI211_X1 g_75_101 (.ZN (n_75_101), .A (n_71_103), .B (n_65_106), .C1 (n_67_106), .C2 (n_61_109) );
AOI211_X1 g_77_100 (.ZN (n_77_100), .A (n_73_102), .B (n_67_105), .C1 (n_66_108), .C2 (n_63_108) );
AOI211_X1 g_79_99 (.ZN (n_79_99), .A (n_75_101), .B (n_69_104), .C1 (n_65_106), .C2 (n_65_107) );
AOI211_X1 g_80_97 (.ZN (n_80_97), .A (n_77_100), .B (n_71_103), .C1 (n_67_105), .C2 (n_67_106) );
AOI211_X1 g_82_96 (.ZN (n_82_96), .A (n_79_99), .B (n_73_102), .C1 (n_69_104), .C2 (n_66_108) );
AOI211_X1 g_84_95 (.ZN (n_84_95), .A (n_80_97), .B (n_75_101), .C1 (n_71_103), .C2 (n_65_106) );
AOI211_X1 g_86_94 (.ZN (n_86_94), .A (n_82_96), .B (n_77_100), .C1 (n_73_102), .C2 (n_67_105) );
AOI211_X1 g_88_93 (.ZN (n_88_93), .A (n_84_95), .B (n_79_99), .C1 (n_75_101), .C2 (n_69_104) );
AOI211_X1 g_90_92 (.ZN (n_90_92), .A (n_86_94), .B (n_80_97), .C1 (n_77_100), .C2 (n_71_103) );
AOI211_X1 g_92_91 (.ZN (n_92_91), .A (n_88_93), .B (n_82_96), .C1 (n_79_99), .C2 (n_73_102) );
AOI211_X1 g_94_90 (.ZN (n_94_90), .A (n_90_92), .B (n_84_95), .C1 (n_80_97), .C2 (n_75_101) );
AOI211_X1 g_96_89 (.ZN (n_96_89), .A (n_92_91), .B (n_86_94), .C1 (n_82_96), .C2 (n_77_100) );
AOI211_X1 g_98_88 (.ZN (n_98_88), .A (n_94_90), .B (n_88_93), .C1 (n_84_95), .C2 (n_79_99) );
AOI211_X1 g_100_87 (.ZN (n_100_87), .A (n_96_89), .B (n_90_92), .C1 (n_86_94), .C2 (n_80_97) );
AOI211_X1 g_102_86 (.ZN (n_102_86), .A (n_98_88), .B (n_92_91), .C1 (n_88_93), .C2 (n_82_96) );
AOI211_X1 g_104_85 (.ZN (n_104_85), .A (n_100_87), .B (n_94_90), .C1 (n_90_92), .C2 (n_84_95) );
AOI211_X1 g_106_84 (.ZN (n_106_84), .A (n_102_86), .B (n_96_89), .C1 (n_92_91), .C2 (n_86_94) );
AOI211_X1 g_108_83 (.ZN (n_108_83), .A (n_104_85), .B (n_98_88), .C1 (n_94_90), .C2 (n_88_93) );
AOI211_X1 g_110_84 (.ZN (n_110_84), .A (n_106_84), .B (n_100_87), .C1 (n_96_89), .C2 (n_90_92) );
AOI211_X1 g_108_85 (.ZN (n_108_85), .A (n_108_83), .B (n_102_86), .C1 (n_98_88), .C2 (n_92_91) );
AOI211_X1 g_106_86 (.ZN (n_106_86), .A (n_110_84), .B (n_104_85), .C1 (n_100_87), .C2 (n_94_90) );
AOI211_X1 g_104_87 (.ZN (n_104_87), .A (n_108_85), .B (n_106_84), .C1 (n_102_86), .C2 (n_96_89) );
AOI211_X1 g_102_88 (.ZN (n_102_88), .A (n_106_86), .B (n_108_83), .C1 (n_104_85), .C2 (n_98_88) );
AOI211_X1 g_100_89 (.ZN (n_100_89), .A (n_104_87), .B (n_110_84), .C1 (n_106_84), .C2 (n_100_87) );
AOI211_X1 g_98_90 (.ZN (n_98_90), .A (n_102_88), .B (n_108_85), .C1 (n_108_83), .C2 (n_102_86) );
AOI211_X1 g_96_91 (.ZN (n_96_91), .A (n_100_89), .B (n_106_86), .C1 (n_110_84), .C2 (n_104_85) );
AOI211_X1 g_94_92 (.ZN (n_94_92), .A (n_98_90), .B (n_104_87), .C1 (n_108_85), .C2 (n_106_84) );
AOI211_X1 g_92_93 (.ZN (n_92_93), .A (n_96_91), .B (n_102_88), .C1 (n_106_86), .C2 (n_108_83) );
AOI211_X1 g_93_91 (.ZN (n_93_91), .A (n_94_92), .B (n_100_89), .C1 (n_104_87), .C2 (n_110_84) );
AOI211_X1 g_91_92 (.ZN (n_91_92), .A (n_92_93), .B (n_98_90), .C1 (n_102_88), .C2 (n_108_85) );
AOI211_X1 g_89_93 (.ZN (n_89_93), .A (n_93_91), .B (n_96_91), .C1 (n_100_89), .C2 (n_106_86) );
AOI211_X1 g_87_94 (.ZN (n_87_94), .A (n_91_92), .B (n_94_92), .C1 (n_98_90), .C2 (n_104_87) );
AOI211_X1 g_85_95 (.ZN (n_85_95), .A (n_89_93), .B (n_92_93), .C1 (n_96_91), .C2 (n_102_88) );
AOI211_X1 g_83_96 (.ZN (n_83_96), .A (n_87_94), .B (n_93_91), .C1 (n_94_92), .C2 (n_100_89) );
AOI211_X1 g_81_97 (.ZN (n_81_97), .A (n_85_95), .B (n_91_92), .C1 (n_92_93), .C2 (n_98_90) );
AOI211_X1 g_79_98 (.ZN (n_79_98), .A (n_83_96), .B (n_89_93), .C1 (n_93_91), .C2 (n_96_91) );
AOI211_X1 g_81_99 (.ZN (n_81_99), .A (n_81_97), .B (n_87_94), .C1 (n_91_92), .C2 (n_94_92) );
AOI211_X1 g_83_98 (.ZN (n_83_98), .A (n_79_98), .B (n_85_95), .C1 (n_89_93), .C2 (n_92_93) );
AOI211_X1 g_84_96 (.ZN (n_84_96), .A (n_81_99), .B (n_83_96), .C1 (n_87_94), .C2 (n_93_91) );
AOI211_X1 g_86_95 (.ZN (n_86_95), .A (n_83_98), .B (n_81_97), .C1 (n_85_95), .C2 (n_91_92) );
AOI211_X1 g_88_94 (.ZN (n_88_94), .A (n_84_96), .B (n_79_98), .C1 (n_83_96), .C2 (n_89_93) );
AOI211_X1 g_87_96 (.ZN (n_87_96), .A (n_86_95), .B (n_81_99), .C1 (n_81_97), .C2 (n_87_94) );
AOI211_X1 g_85_97 (.ZN (n_85_97), .A (n_88_94), .B (n_83_98), .C1 (n_79_98), .C2 (n_85_95) );
AOI211_X1 g_84_99 (.ZN (n_84_99), .A (n_87_96), .B (n_84_96), .C1 (n_81_99), .C2 (n_83_96) );
AOI211_X1 g_83_97 (.ZN (n_83_97), .A (n_85_97), .B (n_86_95), .C1 (n_83_98), .C2 (n_81_97) );
AOI211_X1 g_81_98 (.ZN (n_81_98), .A (n_84_99), .B (n_88_94), .C1 (n_84_96), .C2 (n_79_98) );
AOI211_X1 g_80_100 (.ZN (n_80_100), .A (n_83_97), .B (n_87_96), .C1 (n_86_95), .C2 (n_81_99) );
AOI211_X1 g_82_99 (.ZN (n_82_99), .A (n_81_98), .B (n_85_97), .C1 (n_88_94), .C2 (n_83_98) );
AOI211_X1 g_84_98 (.ZN (n_84_98), .A (n_80_100), .B (n_84_99), .C1 (n_87_96), .C2 (n_84_96) );
AOI211_X1 g_85_96 (.ZN (n_85_96), .A (n_82_99), .B (n_83_97), .C1 (n_85_97), .C2 (n_86_95) );
AOI211_X1 g_87_95 (.ZN (n_87_95), .A (n_84_98), .B (n_81_98), .C1 (n_84_99), .C2 (n_88_94) );
AOI211_X1 g_89_94 (.ZN (n_89_94), .A (n_85_96), .B (n_80_100), .C1 (n_83_97), .C2 (n_87_96) );
AOI211_X1 g_91_93 (.ZN (n_91_93), .A (n_87_95), .B (n_82_99), .C1 (n_81_98), .C2 (n_85_97) );
AOI211_X1 g_93_92 (.ZN (n_93_92), .A (n_89_94), .B (n_84_98), .C1 (n_80_100), .C2 (n_84_99) );
AOI211_X1 g_95_91 (.ZN (n_95_91), .A (n_91_93), .B (n_85_96), .C1 (n_82_99), .C2 (n_83_97) );
AOI211_X1 g_97_90 (.ZN (n_97_90), .A (n_93_92), .B (n_87_95), .C1 (n_84_98), .C2 (n_81_98) );
AOI211_X1 g_99_89 (.ZN (n_99_89), .A (n_95_91), .B (n_89_94), .C1 (n_85_96), .C2 (n_80_100) );
AOI211_X1 g_101_88 (.ZN (n_101_88), .A (n_97_90), .B (n_91_93), .C1 (n_87_95), .C2 (n_82_99) );
AOI211_X1 g_103_87 (.ZN (n_103_87), .A (n_99_89), .B (n_93_92), .C1 (n_89_94), .C2 (n_84_98) );
AOI211_X1 g_105_86 (.ZN (n_105_86), .A (n_101_88), .B (n_95_91), .C1 (n_91_93), .C2 (n_85_96) );
AOI211_X1 g_107_85 (.ZN (n_107_85), .A (n_103_87), .B (n_97_90), .C1 (n_93_92), .C2 (n_87_95) );
AOI211_X1 g_109_84 (.ZN (n_109_84), .A (n_105_86), .B (n_99_89), .C1 (n_95_91), .C2 (n_89_94) );
AOI211_X1 g_111_83 (.ZN (n_111_83), .A (n_107_85), .B (n_101_88), .C1 (n_97_90), .C2 (n_91_93) );
AOI211_X1 g_110_85 (.ZN (n_110_85), .A (n_109_84), .B (n_103_87), .C1 (n_99_89), .C2 (n_93_92) );
AOI211_X1 g_112_84 (.ZN (n_112_84), .A (n_111_83), .B (n_105_86), .C1 (n_101_88), .C2 (n_95_91) );
AOI211_X1 g_114_83 (.ZN (n_114_83), .A (n_110_85), .B (n_107_85), .C1 (n_103_87), .C2 (n_97_90) );
AOI211_X1 g_116_82 (.ZN (n_116_82), .A (n_112_84), .B (n_109_84), .C1 (n_105_86), .C2 (n_99_89) );
AOI211_X1 g_118_81 (.ZN (n_118_81), .A (n_114_83), .B (n_111_83), .C1 (n_107_85), .C2 (n_101_88) );
AOI211_X1 g_120_80 (.ZN (n_120_80), .A (n_116_82), .B (n_110_85), .C1 (n_109_84), .C2 (n_103_87) );
AOI211_X1 g_122_79 (.ZN (n_122_79), .A (n_118_81), .B (n_112_84), .C1 (n_111_83), .C2 (n_105_86) );
AOI211_X1 g_124_78 (.ZN (n_124_78), .A (n_120_80), .B (n_114_83), .C1 (n_110_85), .C2 (n_107_85) );
AOI211_X1 g_126_77 (.ZN (n_126_77), .A (n_122_79), .B (n_116_82), .C1 (n_112_84), .C2 (n_109_84) );
AOI211_X1 g_128_78 (.ZN (n_128_78), .A (n_124_78), .B (n_118_81), .C1 (n_114_83), .C2 (n_111_83) );
AOI211_X1 g_130_77 (.ZN (n_130_77), .A (n_126_77), .B (n_120_80), .C1 (n_116_82), .C2 (n_110_85) );
AOI211_X1 g_132_76 (.ZN (n_132_76), .A (n_128_78), .B (n_122_79), .C1 (n_118_81), .C2 (n_112_84) );
AOI211_X1 g_134_75 (.ZN (n_134_75), .A (n_130_77), .B (n_124_78), .C1 (n_120_80), .C2 (n_114_83) );
AOI211_X1 g_136_74 (.ZN (n_136_74), .A (n_132_76), .B (n_126_77), .C1 (n_122_79), .C2 (n_116_82) );
AOI211_X1 g_138_73 (.ZN (n_138_73), .A (n_134_75), .B (n_128_78), .C1 (n_124_78), .C2 (n_118_81) );
AOI211_X1 g_140_72 (.ZN (n_140_72), .A (n_136_74), .B (n_130_77), .C1 (n_126_77), .C2 (n_120_80) );
AOI211_X1 g_142_71 (.ZN (n_142_71), .A (n_138_73), .B (n_132_76), .C1 (n_128_78), .C2 (n_122_79) );
AOI211_X1 g_144_70 (.ZN (n_144_70), .A (n_140_72), .B (n_134_75), .C1 (n_130_77), .C2 (n_124_78) );
AOI211_X1 g_146_71 (.ZN (n_146_71), .A (n_142_71), .B (n_136_74), .C1 (n_132_76), .C2 (n_126_77) );
AOI211_X1 g_144_72 (.ZN (n_144_72), .A (n_144_70), .B (n_138_73), .C1 (n_134_75), .C2 (n_128_78) );
AOI211_X1 g_142_73 (.ZN (n_142_73), .A (n_146_71), .B (n_140_72), .C1 (n_136_74), .C2 (n_130_77) );
AOI211_X1 g_141_71 (.ZN (n_141_71), .A (n_144_72), .B (n_142_71), .C1 (n_138_73), .C2 (n_132_76) );
AOI211_X1 g_139_72 (.ZN (n_139_72), .A (n_142_73), .B (n_144_70), .C1 (n_140_72), .C2 (n_134_75) );
AOI211_X1 g_137_73 (.ZN (n_137_73), .A (n_141_71), .B (n_146_71), .C1 (n_142_71), .C2 (n_136_74) );
AOI211_X1 g_135_74 (.ZN (n_135_74), .A (n_139_72), .B (n_144_72), .C1 (n_144_70), .C2 (n_138_73) );
AOI211_X1 g_133_75 (.ZN (n_133_75), .A (n_137_73), .B (n_142_73), .C1 (n_146_71), .C2 (n_140_72) );
AOI211_X1 g_131_76 (.ZN (n_131_76), .A (n_135_74), .B (n_141_71), .C1 (n_144_72), .C2 (n_142_71) );
AOI211_X1 g_129_77 (.ZN (n_129_77), .A (n_133_75), .B (n_139_72), .C1 (n_142_73), .C2 (n_144_70) );
AOI211_X1 g_127_78 (.ZN (n_127_78), .A (n_131_76), .B (n_137_73), .C1 (n_141_71), .C2 (n_146_71) );
AOI211_X1 g_125_77 (.ZN (n_125_77), .A (n_129_77), .B (n_135_74), .C1 (n_139_72), .C2 (n_144_72) );
AOI211_X1 g_123_78 (.ZN (n_123_78), .A (n_127_78), .B (n_133_75), .C1 (n_137_73), .C2 (n_142_73) );
AOI211_X1 g_121_79 (.ZN (n_121_79), .A (n_125_77), .B (n_131_76), .C1 (n_135_74), .C2 (n_141_71) );
AOI211_X1 g_119_80 (.ZN (n_119_80), .A (n_123_78), .B (n_129_77), .C1 (n_133_75), .C2 (n_139_72) );
AOI211_X1 g_117_81 (.ZN (n_117_81), .A (n_121_79), .B (n_127_78), .C1 (n_131_76), .C2 (n_137_73) );
AOI211_X1 g_115_82 (.ZN (n_115_82), .A (n_119_80), .B (n_125_77), .C1 (n_129_77), .C2 (n_135_74) );
AOI211_X1 g_113_83 (.ZN (n_113_83), .A (n_117_81), .B (n_123_78), .C1 (n_127_78), .C2 (n_133_75) );
AOI211_X1 g_111_84 (.ZN (n_111_84), .A (n_115_82), .B (n_121_79), .C1 (n_125_77), .C2 (n_131_76) );
AOI211_X1 g_109_85 (.ZN (n_109_85), .A (n_113_83), .B (n_119_80), .C1 (n_123_78), .C2 (n_129_77) );
AOI211_X1 g_107_86 (.ZN (n_107_86), .A (n_111_84), .B (n_117_81), .C1 (n_121_79), .C2 (n_127_78) );
AOI211_X1 g_105_87 (.ZN (n_105_87), .A (n_109_85), .B (n_115_82), .C1 (n_119_80), .C2 (n_125_77) );
AOI211_X1 g_103_88 (.ZN (n_103_88), .A (n_107_86), .B (n_113_83), .C1 (n_117_81), .C2 (n_123_78) );
AOI211_X1 g_101_89 (.ZN (n_101_89), .A (n_105_87), .B (n_111_84), .C1 (n_115_82), .C2 (n_121_79) );
AOI211_X1 g_99_90 (.ZN (n_99_90), .A (n_103_88), .B (n_109_85), .C1 (n_113_83), .C2 (n_119_80) );
AOI211_X1 g_97_91 (.ZN (n_97_91), .A (n_101_89), .B (n_107_86), .C1 (n_111_84), .C2 (n_117_81) );
AOI211_X1 g_95_92 (.ZN (n_95_92), .A (n_99_90), .B (n_105_87), .C1 (n_109_85), .C2 (n_115_82) );
AOI211_X1 g_93_93 (.ZN (n_93_93), .A (n_97_91), .B (n_103_88), .C1 (n_107_86), .C2 (n_113_83) );
AOI211_X1 g_91_94 (.ZN (n_91_94), .A (n_95_92), .B (n_101_89), .C1 (n_105_87), .C2 (n_111_84) );
AOI211_X1 g_89_95 (.ZN (n_89_95), .A (n_93_93), .B (n_99_90), .C1 (n_103_88), .C2 (n_109_85) );
AOI211_X1 g_88_97 (.ZN (n_88_97), .A (n_91_94), .B (n_97_91), .C1 (n_101_89), .C2 (n_107_86) );
AOI211_X1 g_86_96 (.ZN (n_86_96), .A (n_89_95), .B (n_95_92), .C1 (n_99_90), .C2 (n_105_87) );
AOI211_X1 g_88_95 (.ZN (n_88_95), .A (n_88_97), .B (n_93_93), .C1 (n_97_91), .C2 (n_103_88) );
AOI211_X1 g_90_94 (.ZN (n_90_94), .A (n_86_96), .B (n_91_94), .C1 (n_95_92), .C2 (n_101_89) );
AOI211_X1 g_89_96 (.ZN (n_89_96), .A (n_88_95), .B (n_89_95), .C1 (n_93_93), .C2 (n_99_90) );
AOI211_X1 g_91_95 (.ZN (n_91_95), .A (n_90_94), .B (n_88_97), .C1 (n_91_94), .C2 (n_97_91) );
AOI211_X1 g_93_94 (.ZN (n_93_94), .A (n_89_96), .B (n_86_96), .C1 (n_89_95), .C2 (n_95_92) );
AOI211_X1 g_95_93 (.ZN (n_95_93), .A (n_91_95), .B (n_88_95), .C1 (n_88_97), .C2 (n_93_93) );
AOI211_X1 g_97_92 (.ZN (n_97_92), .A (n_93_94), .B (n_90_94), .C1 (n_86_96), .C2 (n_91_94) );
AOI211_X1 g_99_91 (.ZN (n_99_91), .A (n_95_93), .B (n_89_96), .C1 (n_88_95), .C2 (n_89_95) );
AOI211_X1 g_101_90 (.ZN (n_101_90), .A (n_97_92), .B (n_91_95), .C1 (n_90_94), .C2 (n_88_97) );
AOI211_X1 g_103_89 (.ZN (n_103_89), .A (n_99_91), .B (n_93_94), .C1 (n_89_96), .C2 (n_86_96) );
AOI211_X1 g_105_88 (.ZN (n_105_88), .A (n_101_90), .B (n_95_93), .C1 (n_91_95), .C2 (n_88_95) );
AOI211_X1 g_107_87 (.ZN (n_107_87), .A (n_103_89), .B (n_97_92), .C1 (n_93_94), .C2 (n_90_94) );
AOI211_X1 g_109_86 (.ZN (n_109_86), .A (n_105_88), .B (n_99_91), .C1 (n_95_93), .C2 (n_89_96) );
AOI211_X1 g_111_85 (.ZN (n_111_85), .A (n_107_87), .B (n_101_90), .C1 (n_97_92), .C2 (n_91_95) );
AOI211_X1 g_113_84 (.ZN (n_113_84), .A (n_109_86), .B (n_103_89), .C1 (n_99_91), .C2 (n_93_94) );
AOI211_X1 g_114_82 (.ZN (n_114_82), .A (n_111_85), .B (n_105_88), .C1 (n_101_90), .C2 (n_95_93) );
AOI211_X1 g_116_81 (.ZN (n_116_81), .A (n_113_84), .B (n_107_87), .C1 (n_103_89), .C2 (n_97_92) );
AOI211_X1 g_118_80 (.ZN (n_118_80), .A (n_114_82), .B (n_109_86), .C1 (n_105_88), .C2 (n_99_91) );
AOI211_X1 g_117_82 (.ZN (n_117_82), .A (n_116_81), .B (n_111_85), .C1 (n_107_87), .C2 (n_101_90) );
AOI211_X1 g_115_83 (.ZN (n_115_83), .A (n_118_80), .B (n_113_84), .C1 (n_109_86), .C2 (n_103_89) );
AOI211_X1 g_114_85 (.ZN (n_114_85), .A (n_117_82), .B (n_114_82), .C1 (n_111_85), .C2 (n_105_88) );
AOI211_X1 g_116_84 (.ZN (n_116_84), .A (n_115_83), .B (n_116_81), .C1 (n_113_84), .C2 (n_107_87) );
AOI211_X1 g_118_83 (.ZN (n_118_83), .A (n_114_85), .B (n_118_80), .C1 (n_114_82), .C2 (n_109_86) );
AOI211_X1 g_119_81 (.ZN (n_119_81), .A (n_116_84), .B (n_117_82), .C1 (n_116_81), .C2 (n_111_85) );
AOI211_X1 g_121_80 (.ZN (n_121_80), .A (n_118_83), .B (n_115_83), .C1 (n_118_80), .C2 (n_113_84) );
AOI211_X1 g_123_79 (.ZN (n_123_79), .A (n_119_81), .B (n_114_85), .C1 (n_117_82), .C2 (n_114_82) );
AOI211_X1 g_125_78 (.ZN (n_125_78), .A (n_121_80), .B (n_116_84), .C1 (n_115_83), .C2 (n_116_81) );
AOI211_X1 g_124_80 (.ZN (n_124_80), .A (n_123_79), .B (n_118_83), .C1 (n_114_85), .C2 (n_118_80) );
AOI211_X1 g_126_79 (.ZN (n_126_79), .A (n_125_78), .B (n_119_81), .C1 (n_116_84), .C2 (n_117_82) );
AOI211_X1 g_128_80 (.ZN (n_128_80), .A (n_124_80), .B (n_121_80), .C1 (n_118_83), .C2 (n_115_83) );
AOI211_X1 g_129_78 (.ZN (n_129_78), .A (n_126_79), .B (n_123_79), .C1 (n_119_81), .C2 (n_114_85) );
AOI211_X1 g_131_77 (.ZN (n_131_77), .A (n_128_80), .B (n_125_78), .C1 (n_121_80), .C2 (n_116_84) );
AOI211_X1 g_133_76 (.ZN (n_133_76), .A (n_129_78), .B (n_124_80), .C1 (n_123_79), .C2 (n_118_83) );
AOI211_X1 g_132_78 (.ZN (n_132_78), .A (n_131_77), .B (n_126_79), .C1 (n_125_78), .C2 (n_119_81) );
AOI211_X1 g_130_79 (.ZN (n_130_79), .A (n_133_76), .B (n_128_80), .C1 (n_124_80), .C2 (n_121_80) );
AOI211_X1 g_129_81 (.ZN (n_129_81), .A (n_132_78), .B (n_129_78), .C1 (n_126_79), .C2 (n_123_79) );
AOI211_X1 g_128_79 (.ZN (n_128_79), .A (n_130_79), .B (n_131_77), .C1 (n_128_80), .C2 (n_125_78) );
AOI211_X1 g_126_78 (.ZN (n_126_78), .A (n_129_81), .B (n_133_76), .C1 (n_129_78), .C2 (n_124_80) );
AOI211_X1 g_128_77 (.ZN (n_128_77), .A (n_128_79), .B (n_132_78), .C1 (n_131_77), .C2 (n_126_79) );
AOI211_X1 g_127_79 (.ZN (n_127_79), .A (n_126_78), .B (n_130_79), .C1 (n_133_76), .C2 (n_128_80) );
AOI211_X1 g_125_80 (.ZN (n_125_80), .A (n_128_77), .B (n_129_81), .C1 (n_132_78), .C2 (n_129_78) );
AOI211_X1 g_123_81 (.ZN (n_123_81), .A (n_127_79), .B (n_128_79), .C1 (n_130_79), .C2 (n_131_77) );
AOI211_X1 g_124_79 (.ZN (n_124_79), .A (n_125_80), .B (n_126_78), .C1 (n_129_81), .C2 (n_133_76) );
AOI211_X1 g_122_80 (.ZN (n_122_80), .A (n_123_81), .B (n_128_77), .C1 (n_128_79), .C2 (n_132_78) );
AOI211_X1 g_120_81 (.ZN (n_120_81), .A (n_124_79), .B (n_127_79), .C1 (n_126_78), .C2 (n_130_79) );
AOI211_X1 g_118_82 (.ZN (n_118_82), .A (n_122_80), .B (n_125_80), .C1 (n_128_77), .C2 (n_129_81) );
AOI211_X1 g_116_83 (.ZN (n_116_83), .A (n_120_81), .B (n_123_81), .C1 (n_127_79), .C2 (n_128_79) );
AOI211_X1 g_114_84 (.ZN (n_114_84), .A (n_118_82), .B (n_124_79), .C1 (n_125_80), .C2 (n_126_78) );
AOI211_X1 g_112_85 (.ZN (n_112_85), .A (n_116_83), .B (n_122_80), .C1 (n_123_81), .C2 (n_128_77) );
AOI211_X1 g_110_86 (.ZN (n_110_86), .A (n_114_84), .B (n_120_81), .C1 (n_124_79), .C2 (n_127_79) );
AOI211_X1 g_108_87 (.ZN (n_108_87), .A (n_112_85), .B (n_118_82), .C1 (n_122_80), .C2 (n_125_80) );
AOI211_X1 g_106_88 (.ZN (n_106_88), .A (n_110_86), .B (n_116_83), .C1 (n_120_81), .C2 (n_123_81) );
AOI211_X1 g_104_89 (.ZN (n_104_89), .A (n_108_87), .B (n_114_84), .C1 (n_118_82), .C2 (n_124_79) );
AOI211_X1 g_102_90 (.ZN (n_102_90), .A (n_106_88), .B (n_112_85), .C1 (n_116_83), .C2 (n_122_80) );
AOI211_X1 g_100_91 (.ZN (n_100_91), .A (n_104_89), .B (n_110_86), .C1 (n_114_84), .C2 (n_120_81) );
AOI211_X1 g_98_92 (.ZN (n_98_92), .A (n_102_90), .B (n_108_87), .C1 (n_112_85), .C2 (n_118_82) );
AOI211_X1 g_96_93 (.ZN (n_96_93), .A (n_100_91), .B (n_106_88), .C1 (n_110_86), .C2 (n_116_83) );
AOI211_X1 g_94_94 (.ZN (n_94_94), .A (n_98_92), .B (n_104_89), .C1 (n_108_87), .C2 (n_114_84) );
AOI211_X1 g_92_95 (.ZN (n_92_95), .A (n_96_93), .B (n_102_90), .C1 (n_106_88), .C2 (n_112_85) );
AOI211_X1 g_90_96 (.ZN (n_90_96), .A (n_94_94), .B (n_100_91), .C1 (n_104_89), .C2 (n_110_86) );
AOI211_X1 g_92_97 (.ZN (n_92_97), .A (n_92_95), .B (n_98_92), .C1 (n_102_90), .C2 (n_108_87) );
AOI211_X1 g_94_96 (.ZN (n_94_96), .A (n_90_96), .B (n_96_93), .C1 (n_100_91), .C2 (n_106_88) );
AOI211_X1 g_96_95 (.ZN (n_96_95), .A (n_92_97), .B (n_94_94), .C1 (n_98_92), .C2 (n_104_89) );
AOI211_X1 g_98_94 (.ZN (n_98_94), .A (n_94_96), .B (n_92_95), .C1 (n_96_93), .C2 (n_102_90) );
AOI211_X1 g_100_93 (.ZN (n_100_93), .A (n_96_95), .B (n_90_96), .C1 (n_94_94), .C2 (n_100_91) );
AOI211_X1 g_102_92 (.ZN (n_102_92), .A (n_98_94), .B (n_92_97), .C1 (n_92_95), .C2 (n_98_92) );
AOI211_X1 g_104_91 (.ZN (n_104_91), .A (n_100_93), .B (n_94_96), .C1 (n_90_96), .C2 (n_96_93) );
AOI211_X1 g_106_90 (.ZN (n_106_90), .A (n_102_92), .B (n_96_95), .C1 (n_92_97), .C2 (n_94_94) );
AOI211_X1 g_108_89 (.ZN (n_108_89), .A (n_104_91), .B (n_98_94), .C1 (n_94_96), .C2 (n_92_95) );
AOI211_X1 g_109_87 (.ZN (n_109_87), .A (n_106_90), .B (n_100_93), .C1 (n_96_95), .C2 (n_90_96) );
AOI211_X1 g_111_86 (.ZN (n_111_86), .A (n_108_89), .B (n_102_92), .C1 (n_98_94), .C2 (n_92_97) );
AOI211_X1 g_113_85 (.ZN (n_113_85), .A (n_109_87), .B (n_104_91), .C1 (n_100_93), .C2 (n_94_96) );
AOI211_X1 g_115_84 (.ZN (n_115_84), .A (n_111_86), .B (n_106_90), .C1 (n_102_92), .C2 (n_96_95) );
AOI211_X1 g_117_83 (.ZN (n_117_83), .A (n_113_85), .B (n_108_89), .C1 (n_104_91), .C2 (n_98_94) );
AOI211_X1 g_119_82 (.ZN (n_119_82), .A (n_115_84), .B (n_109_87), .C1 (n_106_90), .C2 (n_100_93) );
AOI211_X1 g_121_81 (.ZN (n_121_81), .A (n_117_83), .B (n_111_86), .C1 (n_108_89), .C2 (n_102_92) );
AOI211_X1 g_123_80 (.ZN (n_123_80), .A (n_119_82), .B (n_113_85), .C1 (n_109_87), .C2 (n_104_91) );
AOI211_X1 g_125_79 (.ZN (n_125_79), .A (n_121_81), .B (n_115_84), .C1 (n_111_86), .C2 (n_106_90) );
AOI211_X1 g_126_81 (.ZN (n_126_81), .A (n_123_80), .B (n_117_83), .C1 (n_113_85), .C2 (n_108_89) );
AOI211_X1 g_124_82 (.ZN (n_124_82), .A (n_125_79), .B (n_119_82), .C1 (n_115_84), .C2 (n_109_87) );
AOI211_X1 g_122_81 (.ZN (n_122_81), .A (n_126_81), .B (n_121_81), .C1 (n_117_83), .C2 (n_111_86) );
AOI211_X1 g_120_82 (.ZN (n_120_82), .A (n_124_82), .B (n_123_80), .C1 (n_119_82), .C2 (n_113_85) );
AOI211_X1 g_122_83 (.ZN (n_122_83), .A (n_122_81), .B (n_125_79), .C1 (n_121_81), .C2 (n_115_84) );
AOI211_X1 g_120_84 (.ZN (n_120_84), .A (n_120_82), .B (n_126_81), .C1 (n_123_80), .C2 (n_117_83) );
AOI211_X1 g_121_82 (.ZN (n_121_82), .A (n_122_83), .B (n_124_82), .C1 (n_125_79), .C2 (n_119_82) );
AOI211_X1 g_119_83 (.ZN (n_119_83), .A (n_120_84), .B (n_122_81), .C1 (n_126_81), .C2 (n_121_81) );
AOI211_X1 g_117_84 (.ZN (n_117_84), .A (n_121_82), .B (n_120_82), .C1 (n_124_82), .C2 (n_123_80) );
AOI211_X1 g_115_85 (.ZN (n_115_85), .A (n_119_83), .B (n_122_83), .C1 (n_122_81), .C2 (n_125_79) );
AOI211_X1 g_113_86 (.ZN (n_113_86), .A (n_117_84), .B (n_120_84), .C1 (n_120_82), .C2 (n_126_81) );
AOI211_X1 g_111_87 (.ZN (n_111_87), .A (n_115_85), .B (n_121_82), .C1 (n_122_83), .C2 (n_124_82) );
AOI211_X1 g_109_88 (.ZN (n_109_88), .A (n_113_86), .B (n_119_83), .C1 (n_120_84), .C2 (n_122_81) );
AOI211_X1 g_108_86 (.ZN (n_108_86), .A (n_111_87), .B (n_117_84), .C1 (n_121_82), .C2 (n_120_82) );
AOI211_X1 g_107_88 (.ZN (n_107_88), .A (n_109_88), .B (n_115_85), .C1 (n_119_83), .C2 (n_122_83) );
AOI211_X1 g_105_89 (.ZN (n_105_89), .A (n_108_86), .B (n_113_86), .C1 (n_117_84), .C2 (n_120_84) );
AOI211_X1 g_106_87 (.ZN (n_106_87), .A (n_107_88), .B (n_111_87), .C1 (n_115_85), .C2 (n_121_82) );
AOI211_X1 g_104_88 (.ZN (n_104_88), .A (n_105_89), .B (n_109_88), .C1 (n_113_86), .C2 (n_119_83) );
AOI211_X1 g_103_90 (.ZN (n_103_90), .A (n_106_87), .B (n_108_86), .C1 (n_111_87), .C2 (n_117_84) );
AOI211_X1 g_101_91 (.ZN (n_101_91), .A (n_104_88), .B (n_107_88), .C1 (n_109_88), .C2 (n_115_85) );
AOI211_X1 g_102_89 (.ZN (n_102_89), .A (n_103_90), .B (n_105_89), .C1 (n_108_86), .C2 (n_113_86) );
AOI211_X1 g_100_90 (.ZN (n_100_90), .A (n_101_91), .B (n_106_87), .C1 (n_107_88), .C2 (n_111_87) );
AOI211_X1 g_99_92 (.ZN (n_99_92), .A (n_102_89), .B (n_104_88), .C1 (n_105_89), .C2 (n_109_88) );
AOI211_X1 g_97_93 (.ZN (n_97_93), .A (n_100_90), .B (n_103_90), .C1 (n_106_87), .C2 (n_108_86) );
AOI211_X1 g_98_91 (.ZN (n_98_91), .A (n_99_92), .B (n_101_91), .C1 (n_104_88), .C2 (n_107_88) );
AOI211_X1 g_96_92 (.ZN (n_96_92), .A (n_97_93), .B (n_102_89), .C1 (n_103_90), .C2 (n_105_89) );
AOI211_X1 g_95_94 (.ZN (n_95_94), .A (n_98_91), .B (n_100_90), .C1 (n_101_91), .C2 (n_106_87) );
AOI211_X1 g_93_95 (.ZN (n_93_95), .A (n_96_92), .B (n_99_92), .C1 (n_102_89), .C2 (n_104_88) );
AOI211_X1 g_94_93 (.ZN (n_94_93), .A (n_95_94), .B (n_97_93), .C1 (n_100_90), .C2 (n_103_90) );
AOI211_X1 g_92_94 (.ZN (n_92_94), .A (n_93_95), .B (n_98_91), .C1 (n_99_92), .C2 (n_101_91) );
AOI211_X1 g_90_95 (.ZN (n_90_95), .A (n_94_93), .B (n_96_92), .C1 (n_97_93), .C2 (n_102_89) );
AOI211_X1 g_88_96 (.ZN (n_88_96), .A (n_92_94), .B (n_95_94), .C1 (n_98_91), .C2 (n_100_90) );
AOI211_X1 g_86_97 (.ZN (n_86_97), .A (n_90_95), .B (n_93_95), .C1 (n_96_92), .C2 (n_99_92) );
AOI211_X1 g_88_98 (.ZN (n_88_98), .A (n_88_96), .B (n_94_93), .C1 (n_95_94), .C2 (n_97_93) );
AOI211_X1 g_90_97 (.ZN (n_90_97), .A (n_86_97), .B (n_92_94), .C1 (n_93_95), .C2 (n_98_91) );
AOI211_X1 g_92_96 (.ZN (n_92_96), .A (n_88_98), .B (n_90_95), .C1 (n_94_93), .C2 (n_96_92) );
AOI211_X1 g_94_95 (.ZN (n_94_95), .A (n_90_97), .B (n_88_96), .C1 (n_92_94), .C2 (n_95_94) );
AOI211_X1 g_96_94 (.ZN (n_96_94), .A (n_92_96), .B (n_86_97), .C1 (n_90_95), .C2 (n_93_95) );
AOI211_X1 g_98_93 (.ZN (n_98_93), .A (n_94_95), .B (n_88_98), .C1 (n_88_96), .C2 (n_94_93) );
AOI211_X1 g_100_92 (.ZN (n_100_92), .A (n_96_94), .B (n_90_97), .C1 (n_86_97), .C2 (n_92_94) );
AOI211_X1 g_102_91 (.ZN (n_102_91), .A (n_98_93), .B (n_92_96), .C1 (n_88_98), .C2 (n_90_95) );
AOI211_X1 g_104_90 (.ZN (n_104_90), .A (n_100_92), .B (n_94_95), .C1 (n_90_97), .C2 (n_88_96) );
AOI211_X1 g_106_89 (.ZN (n_106_89), .A (n_102_91), .B (n_96_94), .C1 (n_92_96), .C2 (n_86_97) );
AOI211_X1 g_108_88 (.ZN (n_108_88), .A (n_104_90), .B (n_98_93), .C1 (n_94_95), .C2 (n_88_98) );
AOI211_X1 g_110_87 (.ZN (n_110_87), .A (n_106_89), .B (n_100_92), .C1 (n_96_94), .C2 (n_90_97) );
AOI211_X1 g_112_86 (.ZN (n_112_86), .A (n_108_88), .B (n_102_91), .C1 (n_98_93), .C2 (n_92_96) );
AOI211_X1 g_111_88 (.ZN (n_111_88), .A (n_110_87), .B (n_104_90), .C1 (n_100_92), .C2 (n_94_95) );
AOI211_X1 g_113_87 (.ZN (n_113_87), .A (n_112_86), .B (n_106_89), .C1 (n_102_91), .C2 (n_96_94) );
AOI211_X1 g_115_86 (.ZN (n_115_86), .A (n_111_88), .B (n_108_88), .C1 (n_104_90), .C2 (n_98_93) );
AOI211_X1 g_117_85 (.ZN (n_117_85), .A (n_113_87), .B (n_110_87), .C1 (n_106_89), .C2 (n_100_92) );
AOI211_X1 g_119_84 (.ZN (n_119_84), .A (n_115_86), .B (n_112_86), .C1 (n_108_88), .C2 (n_102_91) );
AOI211_X1 g_121_83 (.ZN (n_121_83), .A (n_117_85), .B (n_111_88), .C1 (n_110_87), .C2 (n_104_90) );
AOI211_X1 g_123_82 (.ZN (n_123_82), .A (n_119_84), .B (n_113_87), .C1 (n_112_86), .C2 (n_106_89) );
AOI211_X1 g_125_81 (.ZN (n_125_81), .A (n_121_83), .B (n_115_86), .C1 (n_111_88), .C2 (n_108_88) );
AOI211_X1 g_127_80 (.ZN (n_127_80), .A (n_123_82), .B (n_117_85), .C1 (n_113_87), .C2 (n_110_87) );
AOI211_X1 g_129_79 (.ZN (n_129_79), .A (n_125_81), .B (n_119_84), .C1 (n_115_86), .C2 (n_112_86) );
AOI211_X1 g_131_78 (.ZN (n_131_78), .A (n_127_80), .B (n_121_83), .C1 (n_117_85), .C2 (n_111_88) );
AOI211_X1 g_133_77 (.ZN (n_133_77), .A (n_129_79), .B (n_123_82), .C1 (n_119_84), .C2 (n_113_87) );
AOI211_X1 g_135_76 (.ZN (n_135_76), .A (n_131_78), .B (n_125_81), .C1 (n_121_83), .C2 (n_115_86) );
AOI211_X1 g_137_75 (.ZN (n_137_75), .A (n_133_77), .B (n_127_80), .C1 (n_123_82), .C2 (n_117_85) );
AOI211_X1 g_139_74 (.ZN (n_139_74), .A (n_135_76), .B (n_129_79), .C1 (n_125_81), .C2 (n_119_84) );
AOI211_X1 g_141_73 (.ZN (n_141_73), .A (n_137_75), .B (n_131_78), .C1 (n_127_80), .C2 (n_121_83) );
AOI211_X1 g_143_72 (.ZN (n_143_72), .A (n_139_74), .B (n_133_77), .C1 (n_129_79), .C2 (n_123_82) );
AOI211_X1 g_144_74 (.ZN (n_144_74), .A (n_141_73), .B (n_135_76), .C1 (n_131_78), .C2 (n_125_81) );
AOI211_X1 g_145_72 (.ZN (n_145_72), .A (n_143_72), .B (n_137_75), .C1 (n_133_77), .C2 (n_127_80) );
AOI211_X1 g_146_70 (.ZN (n_146_70), .A (n_144_74), .B (n_139_74), .C1 (n_135_76), .C2 (n_129_79) );
AOI211_X1 g_147_72 (.ZN (n_147_72), .A (n_145_72), .B (n_141_73), .C1 (n_137_75), .C2 (n_131_78) );
AOI211_X1 g_149_73 (.ZN (n_149_73), .A (n_146_70), .B (n_143_72), .C1 (n_139_74), .C2 (n_133_77) );
AOI211_X1 g_148_71 (.ZN (n_148_71), .A (n_147_72), .B (n_144_74), .C1 (n_141_73), .C2 (n_135_76) );
AOI211_X1 g_147_73 (.ZN (n_147_73), .A (n_149_73), .B (n_145_72), .C1 (n_143_72), .C2 (n_137_75) );
AOI211_X1 g_146_75 (.ZN (n_146_75), .A (n_148_71), .B (n_146_70), .C1 (n_144_74), .C2 (n_139_74) );
AOI211_X1 g_145_73 (.ZN (n_145_73), .A (n_147_73), .B (n_147_72), .C1 (n_145_72), .C2 (n_141_73) );
AOI211_X1 g_144_71 (.ZN (n_144_71), .A (n_146_75), .B (n_149_73), .C1 (n_146_70), .C2 (n_143_72) );
AOI211_X1 g_146_72 (.ZN (n_146_72), .A (n_145_73), .B (n_148_71), .C1 (n_147_72), .C2 (n_144_74) );
AOI211_X1 g_147_74 (.ZN (n_147_74), .A (n_144_71), .B (n_147_73), .C1 (n_149_73), .C2 (n_145_72) );
AOI211_X1 g_145_75 (.ZN (n_145_75), .A (n_146_72), .B (n_146_75), .C1 (n_148_71), .C2 (n_146_70) );
AOI211_X1 g_144_73 (.ZN (n_144_73), .A (n_147_74), .B (n_145_73), .C1 (n_147_73), .C2 (n_147_72) );
AOI211_X1 g_142_72 (.ZN (n_142_72), .A (n_145_75), .B (n_144_71), .C1 (n_146_75), .C2 (n_149_73) );
AOI211_X1 g_143_74 (.ZN (n_143_74), .A (n_144_73), .B (n_146_72), .C1 (n_145_73), .C2 (n_148_71) );
AOI211_X1 g_141_75 (.ZN (n_141_75), .A (n_142_72), .B (n_147_74), .C1 (n_144_71), .C2 (n_147_73) );
AOI211_X1 g_140_73 (.ZN (n_140_73), .A (n_143_74), .B (n_145_75), .C1 (n_146_72), .C2 (n_146_75) );
AOI211_X1 g_138_74 (.ZN (n_138_74), .A (n_141_75), .B (n_144_73), .C1 (n_147_74), .C2 (n_145_73) );
AOI211_X1 g_136_75 (.ZN (n_136_75), .A (n_140_73), .B (n_142_72), .C1 (n_145_75), .C2 (n_144_71) );
AOI211_X1 g_134_76 (.ZN (n_134_76), .A (n_138_74), .B (n_143_74), .C1 (n_144_73), .C2 (n_146_72) );
AOI211_X1 g_132_77 (.ZN (n_132_77), .A (n_136_75), .B (n_141_75), .C1 (n_142_72), .C2 (n_147_74) );
AOI211_X1 g_130_78 (.ZN (n_130_78), .A (n_134_76), .B (n_140_73), .C1 (n_143_74), .C2 (n_145_75) );
AOI211_X1 g_131_80 (.ZN (n_131_80), .A (n_132_77), .B (n_138_74), .C1 (n_141_75), .C2 (n_144_73) );
AOI211_X1 g_133_79 (.ZN (n_133_79), .A (n_130_78), .B (n_136_75), .C1 (n_140_73), .C2 (n_142_72) );
AOI211_X1 g_134_77 (.ZN (n_134_77), .A (n_131_80), .B (n_134_76), .C1 (n_138_74), .C2 (n_143_74) );
AOI211_X1 g_136_76 (.ZN (n_136_76), .A (n_133_79), .B (n_132_77), .C1 (n_136_75), .C2 (n_141_75) );
AOI211_X1 g_138_75 (.ZN (n_138_75), .A (n_134_77), .B (n_130_78), .C1 (n_134_76), .C2 (n_140_73) );
AOI211_X1 g_140_74 (.ZN (n_140_74), .A (n_136_76), .B (n_131_80), .C1 (n_132_77), .C2 (n_138_74) );
AOI211_X1 g_139_76 (.ZN (n_139_76), .A (n_138_75), .B (n_133_79), .C1 (n_130_78), .C2 (n_136_75) );
AOI211_X1 g_137_77 (.ZN (n_137_77), .A (n_140_74), .B (n_134_77), .C1 (n_131_80), .C2 (n_134_76) );
AOI211_X1 g_135_78 (.ZN (n_135_78), .A (n_139_76), .B (n_136_76), .C1 (n_133_79), .C2 (n_132_77) );
AOI211_X1 g_134_80 (.ZN (n_134_80), .A (n_137_77), .B (n_138_75), .C1 (n_134_77), .C2 (n_130_78) );
AOI211_X1 g_133_78 (.ZN (n_133_78), .A (n_135_78), .B (n_140_74), .C1 (n_136_76), .C2 (n_131_80) );
AOI211_X1 g_135_77 (.ZN (n_135_77), .A (n_134_80), .B (n_139_76), .C1 (n_138_75), .C2 (n_133_79) );
AOI211_X1 g_137_76 (.ZN (n_137_76), .A (n_133_78), .B (n_137_77), .C1 (n_140_74), .C2 (n_134_77) );
AOI211_X1 g_139_75 (.ZN (n_139_75), .A (n_135_77), .B (n_135_78), .C1 (n_139_76), .C2 (n_136_76) );
AOI211_X1 g_141_74 (.ZN (n_141_74), .A (n_137_76), .B (n_134_80), .C1 (n_137_77), .C2 (n_138_75) );
AOI211_X1 g_143_73 (.ZN (n_143_73), .A (n_139_75), .B (n_133_78), .C1 (n_135_78), .C2 (n_140_74) );
AOI211_X1 g_145_74 (.ZN (n_145_74), .A (n_141_74), .B (n_135_77), .C1 (n_134_80), .C2 (n_139_76) );
AOI211_X1 g_143_75 (.ZN (n_143_75), .A (n_143_73), .B (n_137_76), .C1 (n_133_78), .C2 (n_137_77) );
AOI211_X1 g_141_76 (.ZN (n_141_76), .A (n_145_74), .B (n_139_75), .C1 (n_135_77), .C2 (n_135_78) );
AOI211_X1 g_142_74 (.ZN (n_142_74), .A (n_143_75), .B (n_141_74), .C1 (n_137_76), .C2 (n_134_80) );
AOI211_X1 g_140_75 (.ZN (n_140_75), .A (n_141_76), .B (n_143_73), .C1 (n_139_75), .C2 (n_133_78) );
AOI211_X1 g_138_76 (.ZN (n_138_76), .A (n_142_74), .B (n_145_74), .C1 (n_141_74), .C2 (n_135_77) );
AOI211_X1 g_136_77 (.ZN (n_136_77), .A (n_140_75), .B (n_143_75), .C1 (n_143_73), .C2 (n_137_76) );
AOI211_X1 g_134_78 (.ZN (n_134_78), .A (n_138_76), .B (n_141_76), .C1 (n_145_74), .C2 (n_139_75) );
AOI211_X1 g_132_79 (.ZN (n_132_79), .A (n_136_77), .B (n_142_74), .C1 (n_143_75), .C2 (n_141_74) );
AOI211_X1 g_130_80 (.ZN (n_130_80), .A (n_134_78), .B (n_140_75), .C1 (n_141_76), .C2 (n_143_73) );
AOI211_X1 g_128_81 (.ZN (n_128_81), .A (n_132_79), .B (n_138_76), .C1 (n_142_74), .C2 (n_145_74) );
AOI211_X1 g_126_80 (.ZN (n_126_80), .A (n_130_80), .B (n_136_77), .C1 (n_140_75), .C2 (n_143_75) );
AOI211_X1 g_124_81 (.ZN (n_124_81), .A (n_128_81), .B (n_134_78), .C1 (n_138_76), .C2 (n_141_76) );
AOI211_X1 g_122_82 (.ZN (n_122_82), .A (n_126_80), .B (n_132_79), .C1 (n_136_77), .C2 (n_142_74) );
AOI211_X1 g_120_83 (.ZN (n_120_83), .A (n_124_81), .B (n_130_80), .C1 (n_134_78), .C2 (n_140_75) );
AOI211_X1 g_118_84 (.ZN (n_118_84), .A (n_122_82), .B (n_128_81), .C1 (n_132_79), .C2 (n_138_76) );
AOI211_X1 g_116_85 (.ZN (n_116_85), .A (n_120_83), .B (n_126_80), .C1 (n_130_80), .C2 (n_136_77) );
AOI211_X1 g_114_86 (.ZN (n_114_86), .A (n_118_84), .B (n_124_81), .C1 (n_128_81), .C2 (n_134_78) );
AOI211_X1 g_112_87 (.ZN (n_112_87), .A (n_116_85), .B (n_122_82), .C1 (n_126_80), .C2 (n_132_79) );
AOI211_X1 g_110_88 (.ZN (n_110_88), .A (n_114_86), .B (n_120_83), .C1 (n_124_81), .C2 (n_130_80) );
AOI211_X1 g_112_89 (.ZN (n_112_89), .A (n_112_87), .B (n_118_84), .C1 (n_122_82), .C2 (n_128_81) );
AOI211_X1 g_114_88 (.ZN (n_114_88), .A (n_110_88), .B (n_116_85), .C1 (n_120_83), .C2 (n_126_80) );
AOI211_X1 g_116_87 (.ZN (n_116_87), .A (n_112_89), .B (n_114_86), .C1 (n_118_84), .C2 (n_124_81) );
AOI211_X1 g_118_86 (.ZN (n_118_86), .A (n_114_88), .B (n_112_87), .C1 (n_116_85), .C2 (n_122_82) );
AOI211_X1 g_120_85 (.ZN (n_120_85), .A (n_116_87), .B (n_110_88), .C1 (n_114_86), .C2 (n_120_83) );
AOI211_X1 g_122_84 (.ZN (n_122_84), .A (n_118_86), .B (n_112_89), .C1 (n_112_87), .C2 (n_118_84) );
AOI211_X1 g_124_83 (.ZN (n_124_83), .A (n_120_85), .B (n_114_88), .C1 (n_110_88), .C2 (n_116_85) );
AOI211_X1 g_126_82 (.ZN (n_126_82), .A (n_122_84), .B (n_116_87), .C1 (n_112_89), .C2 (n_114_86) );
AOI211_X1 g_125_84 (.ZN (n_125_84), .A (n_124_83), .B (n_118_86), .C1 (n_114_88), .C2 (n_112_87) );
AOI211_X1 g_123_83 (.ZN (n_123_83), .A (n_126_82), .B (n_120_85), .C1 (n_116_87), .C2 (n_110_88) );
AOI211_X1 g_125_82 (.ZN (n_125_82), .A (n_125_84), .B (n_122_84), .C1 (n_118_86), .C2 (n_112_89) );
AOI211_X1 g_127_81 (.ZN (n_127_81), .A (n_123_83), .B (n_124_83), .C1 (n_120_85), .C2 (n_114_88) );
AOI211_X1 g_129_80 (.ZN (n_129_80), .A (n_125_82), .B (n_126_82), .C1 (n_122_84), .C2 (n_116_87) );
AOI211_X1 g_131_79 (.ZN (n_131_79), .A (n_127_81), .B (n_125_84), .C1 (n_124_83), .C2 (n_118_86) );
AOI211_X1 g_132_81 (.ZN (n_132_81), .A (n_129_80), .B (n_123_83), .C1 (n_126_82), .C2 (n_120_85) );
AOI211_X1 g_130_82 (.ZN (n_130_82), .A (n_131_79), .B (n_125_82), .C1 (n_125_84), .C2 (n_122_84) );
AOI211_X1 g_128_83 (.ZN (n_128_83), .A (n_132_81), .B (n_127_81), .C1 (n_123_83), .C2 (n_124_83) );
AOI211_X1 g_126_84 (.ZN (n_126_84), .A (n_130_82), .B (n_129_80), .C1 (n_125_82), .C2 (n_126_82) );
AOI211_X1 g_127_82 (.ZN (n_127_82), .A (n_128_83), .B (n_131_79), .C1 (n_127_81), .C2 (n_125_84) );
AOI211_X1 g_125_83 (.ZN (n_125_83), .A (n_126_84), .B (n_132_81), .C1 (n_129_80), .C2 (n_123_83) );
AOI211_X1 g_123_84 (.ZN (n_123_84), .A (n_127_82), .B (n_130_82), .C1 (n_131_79), .C2 (n_125_82) );
AOI211_X1 g_121_85 (.ZN (n_121_85), .A (n_125_83), .B (n_128_83), .C1 (n_132_81), .C2 (n_127_81) );
AOI211_X1 g_119_86 (.ZN (n_119_86), .A (n_123_84), .B (n_126_84), .C1 (n_130_82), .C2 (n_129_80) );
AOI211_X1 g_117_87 (.ZN (n_117_87), .A (n_121_85), .B (n_127_82), .C1 (n_128_83), .C2 (n_131_79) );
AOI211_X1 g_118_85 (.ZN (n_118_85), .A (n_119_86), .B (n_125_83), .C1 (n_126_84), .C2 (n_132_81) );
AOI211_X1 g_116_86 (.ZN (n_116_86), .A (n_117_87), .B (n_123_84), .C1 (n_127_82), .C2 (n_130_82) );
AOI211_X1 g_114_87 (.ZN (n_114_87), .A (n_118_85), .B (n_121_85), .C1 (n_125_83), .C2 (n_128_83) );
AOI211_X1 g_112_88 (.ZN (n_112_88), .A (n_116_86), .B (n_119_86), .C1 (n_123_84), .C2 (n_126_84) );
AOI211_X1 g_110_89 (.ZN (n_110_89), .A (n_114_87), .B (n_117_87), .C1 (n_121_85), .C2 (n_127_82) );
AOI211_X1 g_108_90 (.ZN (n_108_90), .A (n_112_88), .B (n_118_85), .C1 (n_119_86), .C2 (n_125_83) );
AOI211_X1 g_106_91 (.ZN (n_106_91), .A (n_110_89), .B (n_116_86), .C1 (n_117_87), .C2 (n_123_84) );
AOI211_X1 g_107_89 (.ZN (n_107_89), .A (n_108_90), .B (n_114_87), .C1 (n_118_85), .C2 (n_121_85) );
AOI211_X1 g_105_90 (.ZN (n_105_90), .A (n_106_91), .B (n_112_88), .C1 (n_116_86), .C2 (n_119_86) );
AOI211_X1 g_103_91 (.ZN (n_103_91), .A (n_107_89), .B (n_110_89), .C1 (n_114_87), .C2 (n_117_87) );
AOI211_X1 g_101_92 (.ZN (n_101_92), .A (n_105_90), .B (n_108_90), .C1 (n_112_88), .C2 (n_118_85) );
AOI211_X1 g_99_93 (.ZN (n_99_93), .A (n_103_91), .B (n_106_91), .C1 (n_110_89), .C2 (n_116_86) );
AOI211_X1 g_97_94 (.ZN (n_97_94), .A (n_101_92), .B (n_107_89), .C1 (n_108_90), .C2 (n_114_87) );
AOI211_X1 g_95_95 (.ZN (n_95_95), .A (n_99_93), .B (n_105_90), .C1 (n_106_91), .C2 (n_112_88) );
AOI211_X1 g_93_96 (.ZN (n_93_96), .A (n_97_94), .B (n_103_91), .C1 (n_107_89), .C2 (n_110_89) );
AOI211_X1 g_91_97 (.ZN (n_91_97), .A (n_95_95), .B (n_101_92), .C1 (n_105_90), .C2 (n_108_90) );
AOI211_X1 g_89_98 (.ZN (n_89_98), .A (n_93_96), .B (n_99_93), .C1 (n_103_91), .C2 (n_106_91) );
AOI211_X1 g_87_97 (.ZN (n_87_97), .A (n_91_97), .B (n_97_94), .C1 (n_101_92), .C2 (n_107_89) );
AOI211_X1 g_85_98 (.ZN (n_85_98), .A (n_89_98), .B (n_95_95), .C1 (n_99_93), .C2 (n_105_90) );
AOI211_X1 g_87_99 (.ZN (n_87_99), .A (n_87_97), .B (n_93_96), .C1 (n_97_94), .C2 (n_103_91) );
AOI211_X1 g_85_100 (.ZN (n_85_100), .A (n_85_98), .B (n_91_97), .C1 (n_95_95), .C2 (n_101_92) );
AOI211_X1 g_86_98 (.ZN (n_86_98), .A (n_87_99), .B (n_89_98), .C1 (n_93_96), .C2 (n_99_93) );
AOI211_X1 g_84_97 (.ZN (n_84_97), .A (n_85_100), .B (n_87_97), .C1 (n_91_97), .C2 (n_97_94) );
AOI211_X1 g_82_98 (.ZN (n_82_98), .A (n_86_98), .B (n_85_98), .C1 (n_89_98), .C2 (n_95_95) );
AOI211_X1 g_80_99 (.ZN (n_80_99), .A (n_84_97), .B (n_87_99), .C1 (n_87_97), .C2 (n_93_96) );
AOI211_X1 g_78_100 (.ZN (n_78_100), .A (n_82_98), .B (n_85_100), .C1 (n_85_98), .C2 (n_91_97) );
AOI211_X1 g_76_101 (.ZN (n_76_101), .A (n_80_99), .B (n_86_98), .C1 (n_87_99), .C2 (n_89_98) );
AOI211_X1 g_74_102 (.ZN (n_74_102), .A (n_78_100), .B (n_84_97), .C1 (n_85_100), .C2 (n_87_97) );
AOI211_X1 g_72_103 (.ZN (n_72_103), .A (n_76_101), .B (n_82_98), .C1 (n_86_98), .C2 (n_85_98) );
AOI211_X1 g_70_104 (.ZN (n_70_104), .A (n_74_102), .B (n_80_99), .C1 (n_84_97), .C2 (n_87_99) );
AOI211_X1 g_68_105 (.ZN (n_68_105), .A (n_72_103), .B (n_78_100), .C1 (n_82_98), .C2 (n_85_100) );
AOI211_X1 g_66_106 (.ZN (n_66_106), .A (n_70_104), .B (n_76_101), .C1 (n_80_99), .C2 (n_86_98) );
AOI211_X1 g_64_107 (.ZN (n_64_107), .A (n_68_105), .B (n_74_102), .C1 (n_78_100), .C2 (n_84_97) );
AOI211_X1 g_62_108 (.ZN (n_62_108), .A (n_66_106), .B (n_72_103), .C1 (n_76_101), .C2 (n_82_98) );
AOI211_X1 g_60_109 (.ZN (n_60_109), .A (n_64_107), .B (n_70_104), .C1 (n_74_102), .C2 (n_80_99) );
AOI211_X1 g_58_110 (.ZN (n_58_110), .A (n_62_108), .B (n_68_105), .C1 (n_72_103), .C2 (n_78_100) );
AOI211_X1 g_56_111 (.ZN (n_56_111), .A (n_60_109), .B (n_66_106), .C1 (n_70_104), .C2 (n_76_101) );
AOI211_X1 g_54_112 (.ZN (n_54_112), .A (n_58_110), .B (n_64_107), .C1 (n_68_105), .C2 (n_74_102) );
AOI211_X1 g_52_113 (.ZN (n_52_113), .A (n_56_111), .B (n_62_108), .C1 (n_66_106), .C2 (n_72_103) );
AOI211_X1 g_50_114 (.ZN (n_50_114), .A (n_54_112), .B (n_60_109), .C1 (n_64_107), .C2 (n_70_104) );
AOI211_X1 g_48_115 (.ZN (n_48_115), .A (n_52_113), .B (n_58_110), .C1 (n_62_108), .C2 (n_68_105) );
AOI211_X1 g_46_116 (.ZN (n_46_116), .A (n_50_114), .B (n_56_111), .C1 (n_60_109), .C2 (n_66_106) );
AOI211_X1 g_44_117 (.ZN (n_44_117), .A (n_48_115), .B (n_54_112), .C1 (n_58_110), .C2 (n_64_107) );
AOI211_X1 g_42_118 (.ZN (n_42_118), .A (n_46_116), .B (n_52_113), .C1 (n_56_111), .C2 (n_62_108) );
AOI211_X1 g_40_119 (.ZN (n_40_119), .A (n_44_117), .B (n_50_114), .C1 (n_54_112), .C2 (n_60_109) );
AOI211_X1 g_38_120 (.ZN (n_38_120), .A (n_42_118), .B (n_48_115), .C1 (n_52_113), .C2 (n_58_110) );
AOI211_X1 g_36_121 (.ZN (n_36_121), .A (n_40_119), .B (n_46_116), .C1 (n_50_114), .C2 (n_56_111) );
AOI211_X1 g_34_122 (.ZN (n_34_122), .A (n_38_120), .B (n_44_117), .C1 (n_48_115), .C2 (n_54_112) );
AOI211_X1 g_32_123 (.ZN (n_32_123), .A (n_36_121), .B (n_42_118), .C1 (n_46_116), .C2 (n_52_113) );
AOI211_X1 g_30_124 (.ZN (n_30_124), .A (n_34_122), .B (n_40_119), .C1 (n_44_117), .C2 (n_50_114) );
AOI211_X1 g_28_125 (.ZN (n_28_125), .A (n_32_123), .B (n_38_120), .C1 (n_42_118), .C2 (n_48_115) );
AOI211_X1 g_26_126 (.ZN (n_26_126), .A (n_30_124), .B (n_36_121), .C1 (n_40_119), .C2 (n_46_116) );
AOI211_X1 g_24_127 (.ZN (n_24_127), .A (n_28_125), .B (n_34_122), .C1 (n_38_120), .C2 (n_44_117) );
AOI211_X1 g_22_128 (.ZN (n_22_128), .A (n_26_126), .B (n_32_123), .C1 (n_36_121), .C2 (n_42_118) );
AOI211_X1 g_20_129 (.ZN (n_20_129), .A (n_24_127), .B (n_30_124), .C1 (n_34_122), .C2 (n_40_119) );
AOI211_X1 g_18_130 (.ZN (n_18_130), .A (n_22_128), .B (n_28_125), .C1 (n_32_123), .C2 (n_38_120) );
AOI211_X1 g_16_131 (.ZN (n_16_131), .A (n_20_129), .B (n_26_126), .C1 (n_30_124), .C2 (n_36_121) );
AOI211_X1 g_14_132 (.ZN (n_14_132), .A (n_18_130), .B (n_24_127), .C1 (n_28_125), .C2 (n_34_122) );
AOI211_X1 g_12_133 (.ZN (n_12_133), .A (n_16_131), .B (n_22_128), .C1 (n_26_126), .C2 (n_32_123) );
AOI211_X1 g_11_135 (.ZN (n_11_135), .A (n_14_132), .B (n_20_129), .C1 (n_24_127), .C2 (n_30_124) );
AOI211_X1 g_10_133 (.ZN (n_10_133), .A (n_12_133), .B (n_18_130), .C1 (n_22_128), .C2 (n_28_125) );
AOI211_X1 g_8_134 (.ZN (n_8_134), .A (n_11_135), .B (n_16_131), .C1 (n_20_129), .C2 (n_26_126) );
AOI211_X1 g_9_136 (.ZN (n_9_136), .A (n_10_133), .B (n_14_132), .C1 (n_18_130), .C2 (n_24_127) );
AOI211_X1 g_8_138 (.ZN (n_8_138), .A (n_8_134), .B (n_12_133), .C1 (n_16_131), .C2 (n_22_128) );
AOI211_X1 g_7_136 (.ZN (n_7_136), .A (n_9_136), .B (n_11_135), .C1 (n_14_132), .C2 (n_20_129) );
AOI211_X1 g_9_135 (.ZN (n_9_135), .A (n_8_138), .B (n_10_133), .C1 (n_12_133), .C2 (n_18_130) );
AOI211_X1 g_10_137 (.ZN (n_10_137), .A (n_7_136), .B (n_8_134), .C1 (n_11_135), .C2 (n_16_131) );
AOI211_X1 g_12_136 (.ZN (n_12_136), .A (n_9_135), .B (n_9_136), .C1 (n_10_133), .C2 (n_14_132) );
AOI211_X1 g_10_135 (.ZN (n_10_135), .A (n_10_137), .B (n_8_138), .C1 (n_8_134), .C2 (n_12_133) );
AOI211_X1 g_12_134 (.ZN (n_12_134), .A (n_12_136), .B (n_7_136), .C1 (n_9_136), .C2 (n_11_135) );
AOI211_X1 g_13_132 (.ZN (n_13_132), .A (n_10_135), .B (n_9_135), .C1 (n_8_138), .C2 (n_10_133) );
AOI211_X1 g_15_131 (.ZN (n_15_131), .A (n_12_134), .B (n_10_137), .C1 (n_7_136), .C2 (n_8_134) );
AOI211_X1 g_14_133 (.ZN (n_14_133), .A (n_13_132), .B (n_12_136), .C1 (n_9_135), .C2 (n_9_136) );
AOI211_X1 g_12_132 (.ZN (n_12_132), .A (n_15_131), .B (n_10_135), .C1 (n_10_137), .C2 (n_8_138) );
AOI211_X1 g_14_131 (.ZN (n_14_131), .A (n_14_133), .B (n_12_134), .C1 (n_12_136), .C2 (n_7_136) );
AOI211_X1 g_16_132 (.ZN (n_16_132), .A (n_12_132), .B (n_13_132), .C1 (n_10_135), .C2 (n_9_135) );
AOI211_X1 g_18_131 (.ZN (n_18_131), .A (n_14_131), .B (n_15_131), .C1 (n_12_134), .C2 (n_10_137) );
AOI211_X1 g_20_130 (.ZN (n_20_130), .A (n_16_132), .B (n_14_133), .C1 (n_13_132), .C2 (n_12_136) );
AOI211_X1 g_22_129 (.ZN (n_22_129), .A (n_18_131), .B (n_12_132), .C1 (n_15_131), .C2 (n_10_135) );
AOI211_X1 g_24_128 (.ZN (n_24_128), .A (n_20_130), .B (n_14_131), .C1 (n_14_133), .C2 (n_12_134) );
AOI211_X1 g_26_127 (.ZN (n_26_127), .A (n_22_129), .B (n_16_132), .C1 (n_12_132), .C2 (n_13_132) );
AOI211_X1 g_28_126 (.ZN (n_28_126), .A (n_24_128), .B (n_18_131), .C1 (n_14_131), .C2 (n_15_131) );
AOI211_X1 g_30_125 (.ZN (n_30_125), .A (n_26_127), .B (n_20_130), .C1 (n_16_132), .C2 (n_14_133) );
AOI211_X1 g_32_124 (.ZN (n_32_124), .A (n_28_126), .B (n_22_129), .C1 (n_18_131), .C2 (n_12_132) );
AOI211_X1 g_34_123 (.ZN (n_34_123), .A (n_30_125), .B (n_24_128), .C1 (n_20_130), .C2 (n_14_131) );
AOI211_X1 g_35_121 (.ZN (n_35_121), .A (n_32_124), .B (n_26_127), .C1 (n_22_129), .C2 (n_16_132) );
AOI211_X1 g_37_120 (.ZN (n_37_120), .A (n_34_123), .B (n_28_126), .C1 (n_24_128), .C2 (n_18_131) );
AOI211_X1 g_39_119 (.ZN (n_39_119), .A (n_35_121), .B (n_30_125), .C1 (n_26_127), .C2 (n_20_130) );
AOI211_X1 g_41_118 (.ZN (n_41_118), .A (n_37_120), .B (n_32_124), .C1 (n_28_126), .C2 (n_22_129) );
AOI211_X1 g_43_117 (.ZN (n_43_117), .A (n_39_119), .B (n_34_123), .C1 (n_30_125), .C2 (n_24_128) );
AOI211_X1 g_45_116 (.ZN (n_45_116), .A (n_41_118), .B (n_35_121), .C1 (n_32_124), .C2 (n_26_127) );
AOI211_X1 g_47_115 (.ZN (n_47_115), .A (n_43_117), .B (n_37_120), .C1 (n_34_123), .C2 (n_28_126) );
AOI211_X1 g_49_114 (.ZN (n_49_114), .A (n_45_116), .B (n_39_119), .C1 (n_35_121), .C2 (n_30_125) );
AOI211_X1 g_51_113 (.ZN (n_51_113), .A (n_47_115), .B (n_41_118), .C1 (n_37_120), .C2 (n_32_124) );
AOI211_X1 g_53_112 (.ZN (n_53_112), .A (n_49_114), .B (n_43_117), .C1 (n_39_119), .C2 (n_34_123) );
AOI211_X1 g_55_111 (.ZN (n_55_111), .A (n_51_113), .B (n_45_116), .C1 (n_41_118), .C2 (n_35_121) );
AOI211_X1 g_57_110 (.ZN (n_57_110), .A (n_53_112), .B (n_47_115), .C1 (n_43_117), .C2 (n_37_120) );
AOI211_X1 g_59_109 (.ZN (n_59_109), .A (n_55_111), .B (n_49_114), .C1 (n_45_116), .C2 (n_39_119) );
AOI211_X1 g_61_108 (.ZN (n_61_108), .A (n_57_110), .B (n_51_113), .C1 (n_47_115), .C2 (n_41_118) );
AOI211_X1 g_63_107 (.ZN (n_63_107), .A (n_59_109), .B (n_53_112), .C1 (n_49_114), .C2 (n_43_117) );
AOI211_X1 g_64_109 (.ZN (n_64_109), .A (n_61_108), .B (n_55_111), .C1 (n_51_113), .C2 (n_45_116) );
AOI211_X1 g_62_110 (.ZN (n_62_110), .A (n_63_107), .B (n_57_110), .C1 (n_53_112), .C2 (n_47_115) );
AOI211_X1 g_60_111 (.ZN (n_60_111), .A (n_64_109), .B (n_59_109), .C1 (n_55_111), .C2 (n_49_114) );
AOI211_X1 g_58_112 (.ZN (n_58_112), .A (n_62_110), .B (n_61_108), .C1 (n_57_110), .C2 (n_51_113) );
AOI211_X1 g_56_113 (.ZN (n_56_113), .A (n_60_111), .B (n_63_107), .C1 (n_59_109), .C2 (n_53_112) );
AOI211_X1 g_54_114 (.ZN (n_54_114), .A (n_58_112), .B (n_64_109), .C1 (n_61_108), .C2 (n_55_111) );
AOI211_X1 g_52_115 (.ZN (n_52_115), .A (n_56_113), .B (n_62_110), .C1 (n_63_107), .C2 (n_57_110) );
AOI211_X1 g_50_116 (.ZN (n_50_116), .A (n_54_114), .B (n_60_111), .C1 (n_64_109), .C2 (n_59_109) );
AOI211_X1 g_48_117 (.ZN (n_48_117), .A (n_52_115), .B (n_58_112), .C1 (n_62_110), .C2 (n_61_108) );
AOI211_X1 g_46_118 (.ZN (n_46_118), .A (n_50_116), .B (n_56_113), .C1 (n_60_111), .C2 (n_63_107) );
AOI211_X1 g_44_119 (.ZN (n_44_119), .A (n_48_117), .B (n_54_114), .C1 (n_58_112), .C2 (n_64_109) );
AOI211_X1 g_42_120 (.ZN (n_42_120), .A (n_46_118), .B (n_52_115), .C1 (n_56_113), .C2 (n_62_110) );
AOI211_X1 g_40_121 (.ZN (n_40_121), .A (n_44_119), .B (n_50_116), .C1 (n_54_114), .C2 (n_60_111) );
AOI211_X1 g_38_122 (.ZN (n_38_122), .A (n_42_120), .B (n_48_117), .C1 (n_52_115), .C2 (n_58_112) );
AOI211_X1 g_36_123 (.ZN (n_36_123), .A (n_40_121), .B (n_46_118), .C1 (n_50_116), .C2 (n_56_113) );
AOI211_X1 g_34_124 (.ZN (n_34_124), .A (n_38_122), .B (n_44_119), .C1 (n_48_117), .C2 (n_54_114) );
AOI211_X1 g_32_125 (.ZN (n_32_125), .A (n_36_123), .B (n_42_120), .C1 (n_46_118), .C2 (n_52_115) );
AOI211_X1 g_30_126 (.ZN (n_30_126), .A (n_34_124), .B (n_40_121), .C1 (n_44_119), .C2 (n_50_116) );
AOI211_X1 g_28_127 (.ZN (n_28_127), .A (n_32_125), .B (n_38_122), .C1 (n_42_120), .C2 (n_48_117) );
AOI211_X1 g_26_128 (.ZN (n_26_128), .A (n_30_126), .B (n_36_123), .C1 (n_40_121), .C2 (n_46_118) );
AOI211_X1 g_24_129 (.ZN (n_24_129), .A (n_28_127), .B (n_34_124), .C1 (n_38_122), .C2 (n_44_119) );
AOI211_X1 g_22_130 (.ZN (n_22_130), .A (n_26_128), .B (n_32_125), .C1 (n_36_123), .C2 (n_42_120) );
AOI211_X1 g_20_131 (.ZN (n_20_131), .A (n_24_129), .B (n_30_126), .C1 (n_34_124), .C2 (n_40_121) );
AOI211_X1 g_21_129 (.ZN (n_21_129), .A (n_22_130), .B (n_28_127), .C1 (n_32_125), .C2 (n_38_122) );
AOI211_X1 g_19_130 (.ZN (n_19_130), .A (n_20_131), .B (n_26_128), .C1 (n_30_126), .C2 (n_36_123) );
AOI211_X1 g_17_131 (.ZN (n_17_131), .A (n_21_129), .B (n_24_129), .C1 (n_28_127), .C2 (n_34_124) );
AOI211_X1 g_15_132 (.ZN (n_15_132), .A (n_19_130), .B (n_22_130), .C1 (n_26_128), .C2 (n_32_125) );
AOI211_X1 g_13_133 (.ZN (n_13_133), .A (n_17_131), .B (n_20_131), .C1 (n_24_129), .C2 (n_30_126) );
AOI211_X1 g_11_134 (.ZN (n_11_134), .A (n_15_132), .B (n_21_129), .C1 (n_22_130), .C2 (n_28_127) );
AOI211_X1 g_10_136 (.ZN (n_10_136), .A (n_13_133), .B (n_19_130), .C1 (n_20_131), .C2 (n_26_128) );
AOI211_X1 g_12_135 (.ZN (n_12_135), .A (n_11_134), .B (n_17_131), .C1 (n_21_129), .C2 (n_24_129) );
AOI211_X1 g_14_134 (.ZN (n_14_134), .A (n_10_136), .B (n_15_132), .C1 (n_19_130), .C2 (n_22_130) );
AOI211_X1 g_16_133 (.ZN (n_16_133), .A (n_12_135), .B (n_13_133), .C1 (n_17_131), .C2 (n_20_131) );
AOI211_X1 g_18_132 (.ZN (n_18_132), .A (n_14_134), .B (n_11_134), .C1 (n_15_132), .C2 (n_21_129) );
AOI211_X1 g_17_134 (.ZN (n_17_134), .A (n_16_133), .B (n_10_136), .C1 (n_13_133), .C2 (n_19_130) );
AOI211_X1 g_15_133 (.ZN (n_15_133), .A (n_18_132), .B (n_12_135), .C1 (n_11_134), .C2 (n_17_131) );
AOI211_X1 g_13_134 (.ZN (n_13_134), .A (n_17_134), .B (n_14_134), .C1 (n_10_136), .C2 (n_15_132) );
AOI211_X1 g_15_135 (.ZN (n_15_135), .A (n_15_133), .B (n_16_133), .C1 (n_12_135), .C2 (n_13_133) );
AOI211_X1 g_13_136 (.ZN (n_13_136), .A (n_13_134), .B (n_18_132), .C1 (n_14_134), .C2 (n_11_134) );
AOI211_X1 g_11_137 (.ZN (n_11_137), .A (n_15_135), .B (n_17_134), .C1 (n_16_133), .C2 (n_10_136) );
AOI211_X1 g_9_138 (.ZN (n_9_138), .A (n_13_136), .B (n_15_133), .C1 (n_18_132), .C2 (n_12_135) );
AOI211_X1 g_7_139 (.ZN (n_7_139), .A (n_11_137), .B (n_13_134), .C1 (n_17_134), .C2 (n_14_134) );
AOI211_X1 g_8_137 (.ZN (n_8_137), .A (n_9_138), .B (n_15_135), .C1 (n_15_133), .C2 (n_16_133) );
AOI211_X1 g_6_138 (.ZN (n_6_138), .A (n_7_139), .B (n_13_136), .C1 (n_13_134), .C2 (n_18_132) );
AOI211_X1 g_5_140 (.ZN (n_5_140), .A (n_8_137), .B (n_11_137), .C1 (n_15_135), .C2 (n_17_134) );
AOI211_X1 g_4_142 (.ZN (n_4_142), .A (n_6_138), .B (n_9_138), .C1 (n_13_136), .C2 (n_15_133) );
AOI211_X1 g_6_141 (.ZN (n_6_141), .A (n_5_140), .B (n_7_139), .C1 (n_11_137), .C2 (n_13_134) );
AOI211_X1 g_5_143 (.ZN (n_5_143), .A (n_4_142), .B (n_8_137), .C1 (n_9_138), .C2 (n_15_135) );
AOI211_X1 g_3_144 (.ZN (n_3_144), .A (n_6_141), .B (n_6_138), .C1 (n_7_139), .C2 (n_13_136) );
AOI211_X1 g_2_146 (.ZN (n_2_146), .A (n_5_143), .B (n_5_140), .C1 (n_8_137), .C2 (n_11_137) );
AOI211_X1 g_1_148 (.ZN (n_1_148), .A (n_3_144), .B (n_4_142), .C1 (n_6_138), .C2 (n_9_138) );
AOI211_X1 g_2_150 (.ZN (n_2_150), .A (n_2_146), .B (n_6_141), .C1 (n_5_140), .C2 (n_7_139) );
AOI211_X1 g_3_148 (.ZN (n_3_148), .A (n_1_148), .B (n_5_143), .C1 (n_4_142), .C2 (n_8_137) );
AOI211_X1 g_4_146 (.ZN (n_4_146), .A (n_2_150), .B (n_3_144), .C1 (n_6_141), .C2 (n_6_138) );
AOI211_X1 g_5_148 (.ZN (n_5_148), .A (n_3_148), .B (n_2_146), .C1 (n_5_143), .C2 (n_5_140) );
AOI211_X1 g_3_147 (.ZN (n_3_147), .A (n_4_146), .B (n_1_148), .C1 (n_3_144), .C2 (n_4_142) );
AOI211_X1 g_4_145 (.ZN (n_4_145), .A (n_5_148), .B (n_2_150), .C1 (n_2_146), .C2 (n_6_141) );
AOI211_X1 g_5_147 (.ZN (n_5_147), .A (n_3_147), .B (n_3_148), .C1 (n_1_148), .C2 (n_5_143) );
AOI211_X1 g_4_149 (.ZN (n_4_149), .A (n_4_145), .B (n_4_146), .C1 (n_2_150), .C2 (n_3_144) );
AOI211_X1 g_6_150 (.ZN (n_6_150), .A (n_5_147), .B (n_5_148), .C1 (n_3_148), .C2 (n_2_146) );
AOI211_X1 g_7_148 (.ZN (n_7_148), .A (n_4_149), .B (n_3_147), .C1 (n_4_146), .C2 (n_1_148) );
AOI211_X1 g_6_146 (.ZN (n_6_146), .A (n_6_150), .B (n_4_145), .C1 (n_5_148), .C2 (n_2_150) );
AOI211_X1 g_4_147 (.ZN (n_4_147), .A (n_7_148), .B (n_5_147), .C1 (n_3_147), .C2 (n_3_148) );
AOI211_X1 g_3_145 (.ZN (n_3_145), .A (n_6_146), .B (n_4_149), .C1 (n_4_145), .C2 (n_4_146) );
AOI211_X1 g_5_144 (.ZN (n_5_144), .A (n_4_147), .B (n_6_150), .C1 (n_5_147), .C2 (n_5_148) );
AOI211_X1 g_7_143 (.ZN (n_7_143), .A (n_3_145), .B (n_7_148), .C1 (n_4_149), .C2 (n_3_147) );
AOI211_X1 g_6_145 (.ZN (n_6_145), .A (n_5_144), .B (n_6_146), .C1 (n_6_150), .C2 (n_4_145) );
AOI211_X1 g_7_147 (.ZN (n_7_147), .A (n_7_143), .B (n_4_147), .C1 (n_7_148), .C2 (n_5_147) );
AOI211_X1 g_5_146 (.ZN (n_5_146), .A (n_6_145), .B (n_3_145), .C1 (n_6_146), .C2 (n_4_149) );
AOI211_X1 g_6_148 (.ZN (n_6_148), .A (n_7_147), .B (n_5_144), .C1 (n_4_147), .C2 (n_6_150) );
AOI211_X1 g_8_149 (.ZN (n_8_149), .A (n_5_146), .B (n_7_143), .C1 (n_3_145), .C2 (n_7_148) );
AOI211_X1 g_10_150 (.ZN (n_10_150), .A (n_6_148), .B (n_6_145), .C1 (n_5_144), .C2 (n_6_146) );
AOI211_X1 g_9_148 (.ZN (n_9_148), .A (n_8_149), .B (n_7_147), .C1 (n_7_143), .C2 (n_4_147) );
AOI211_X1 g_8_146 (.ZN (n_8_146), .A (n_10_150), .B (n_5_146), .C1 (n_6_145), .C2 (n_3_145) );
AOI211_X1 g_6_147 (.ZN (n_6_147), .A (n_9_148), .B (n_6_148), .C1 (n_7_147), .C2 (n_5_144) );
AOI211_X1 g_8_148 (.ZN (n_8_148), .A (n_8_146), .B (n_8_149), .C1 (n_5_146), .C2 (n_7_143) );
AOI211_X1 g_10_147 (.ZN (n_10_147), .A (n_6_147), .B (n_10_150), .C1 (n_6_148), .C2 (n_6_145) );
AOI211_X1 g_12_148 (.ZN (n_12_148), .A (n_8_148), .B (n_9_148), .C1 (n_8_149), .C2 (n_7_147) );
AOI211_X1 g_14_147 (.ZN (n_14_147), .A (n_10_147), .B (n_8_146), .C1 (n_10_150), .C2 (n_5_146) );
AOI211_X1 g_16_148 (.ZN (n_16_148), .A (n_12_148), .B (n_6_147), .C1 (n_9_148), .C2 (n_6_148) );
AOI211_X1 g_18_147 (.ZN (n_18_147), .A (n_14_147), .B (n_8_148), .C1 (n_8_146), .C2 (n_8_149) );
AOI211_X1 g_20_148 (.ZN (n_20_148), .A (n_16_148), .B (n_10_147), .C1 (n_6_147), .C2 (n_10_150) );
AOI211_X1 g_22_147 (.ZN (n_22_147), .A (n_18_147), .B (n_12_148), .C1 (n_8_148), .C2 (n_9_148) );
AOI211_X1 g_24_148 (.ZN (n_24_148), .A (n_20_148), .B (n_14_147), .C1 (n_10_147), .C2 (n_8_146) );
AOI211_X1 g_26_147 (.ZN (n_26_147), .A (n_22_147), .B (n_16_148), .C1 (n_12_148), .C2 (n_6_147) );
AOI211_X1 g_28_148 (.ZN (n_28_148), .A (n_24_148), .B (n_18_147), .C1 (n_14_147), .C2 (n_8_148) );
AOI211_X1 g_30_147 (.ZN (n_30_147), .A (n_26_147), .B (n_20_148), .C1 (n_16_148), .C2 (n_10_147) );
AOI211_X1 g_32_148 (.ZN (n_32_148), .A (n_28_148), .B (n_22_147), .C1 (n_18_147), .C2 (n_12_148) );
AOI211_X1 g_34_147 (.ZN (n_34_147), .A (n_30_147), .B (n_24_148), .C1 (n_20_148), .C2 (n_14_147) );
AOI211_X1 g_36_148 (.ZN (n_36_148), .A (n_32_148), .B (n_26_147), .C1 (n_22_147), .C2 (n_16_148) );
AOI211_X1 g_38_147 (.ZN (n_38_147), .A (n_34_147), .B (n_28_148), .C1 (n_24_148), .C2 (n_18_147) );
AOI211_X1 g_40_148 (.ZN (n_40_148), .A (n_36_148), .B (n_30_147), .C1 (n_26_147), .C2 (n_20_148) );
AOI211_X1 g_42_147 (.ZN (n_42_147), .A (n_38_147), .B (n_32_148), .C1 (n_28_148), .C2 (n_22_147) );
AOI211_X1 g_44_148 (.ZN (n_44_148), .A (n_40_148), .B (n_34_147), .C1 (n_30_147), .C2 (n_24_148) );
AOI211_X1 g_46_147 (.ZN (n_46_147), .A (n_42_147), .B (n_36_148), .C1 (n_32_148), .C2 (n_26_147) );
AOI211_X1 g_48_148 (.ZN (n_48_148), .A (n_44_148), .B (n_38_147), .C1 (n_34_147), .C2 (n_28_148) );
AOI211_X1 g_50_147 (.ZN (n_50_147), .A (n_46_147), .B (n_40_148), .C1 (n_36_148), .C2 (n_30_147) );
AOI211_X1 g_52_148 (.ZN (n_52_148), .A (n_48_148), .B (n_42_147), .C1 (n_38_147), .C2 (n_32_148) );
AOI211_X1 g_54_147 (.ZN (n_54_147), .A (n_50_147), .B (n_44_148), .C1 (n_40_148), .C2 (n_34_147) );
AOI211_X1 g_56_148 (.ZN (n_56_148), .A (n_52_148), .B (n_46_147), .C1 (n_42_147), .C2 (n_36_148) );
AOI211_X1 g_58_147 (.ZN (n_58_147), .A (n_54_147), .B (n_48_148), .C1 (n_44_148), .C2 (n_38_147) );
AOI211_X1 g_60_148 (.ZN (n_60_148), .A (n_56_148), .B (n_50_147), .C1 (n_46_147), .C2 (n_40_148) );
AOI211_X1 g_62_147 (.ZN (n_62_147), .A (n_58_147), .B (n_52_148), .C1 (n_48_148), .C2 (n_42_147) );
AOI211_X1 g_64_148 (.ZN (n_64_148), .A (n_60_148), .B (n_54_147), .C1 (n_50_147), .C2 (n_44_148) );
AOI211_X1 g_66_147 (.ZN (n_66_147), .A (n_62_147), .B (n_56_148), .C1 (n_52_148), .C2 (n_46_147) );
AOI211_X1 g_68_148 (.ZN (n_68_148), .A (n_64_148), .B (n_58_147), .C1 (n_54_147), .C2 (n_48_148) );
AOI211_X1 g_70_147 (.ZN (n_70_147), .A (n_66_147), .B (n_60_148), .C1 (n_56_148), .C2 (n_50_147) );
AOI211_X1 g_72_148 (.ZN (n_72_148), .A (n_68_148), .B (n_62_147), .C1 (n_58_147), .C2 (n_52_148) );
AOI211_X1 g_74_147 (.ZN (n_74_147), .A (n_70_147), .B (n_64_148), .C1 (n_60_148), .C2 (n_54_147) );
AOI211_X1 g_76_148 (.ZN (n_76_148), .A (n_72_148), .B (n_66_147), .C1 (n_62_147), .C2 (n_56_148) );
AOI211_X1 g_78_147 (.ZN (n_78_147), .A (n_74_147), .B (n_68_148), .C1 (n_64_148), .C2 (n_58_147) );
AOI211_X1 g_80_148 (.ZN (n_80_148), .A (n_76_148), .B (n_70_147), .C1 (n_66_147), .C2 (n_60_148) );
AOI211_X1 g_82_147 (.ZN (n_82_147), .A (n_78_147), .B (n_72_148), .C1 (n_68_148), .C2 (n_62_147) );
AOI211_X1 g_84_148 (.ZN (n_84_148), .A (n_80_148), .B (n_74_147), .C1 (n_70_147), .C2 (n_64_148) );
AOI211_X1 g_86_147 (.ZN (n_86_147), .A (n_82_147), .B (n_76_148), .C1 (n_72_148), .C2 (n_66_147) );
AOI211_X1 g_88_148 (.ZN (n_88_148), .A (n_84_148), .B (n_78_147), .C1 (n_74_147), .C2 (n_68_148) );
AOI211_X1 g_90_147 (.ZN (n_90_147), .A (n_86_147), .B (n_80_148), .C1 (n_76_148), .C2 (n_70_147) );
AOI211_X1 g_92_148 (.ZN (n_92_148), .A (n_88_148), .B (n_82_147), .C1 (n_78_147), .C2 (n_72_148) );
AOI211_X1 g_94_147 (.ZN (n_94_147), .A (n_90_147), .B (n_84_148), .C1 (n_80_148), .C2 (n_74_147) );
AOI211_X1 g_96_148 (.ZN (n_96_148), .A (n_92_148), .B (n_86_147), .C1 (n_82_147), .C2 (n_76_148) );
AOI211_X1 g_98_147 (.ZN (n_98_147), .A (n_94_147), .B (n_88_148), .C1 (n_84_148), .C2 (n_78_147) );
AOI211_X1 g_100_148 (.ZN (n_100_148), .A (n_96_148), .B (n_90_147), .C1 (n_86_147), .C2 (n_80_148) );
AOI211_X1 g_102_147 (.ZN (n_102_147), .A (n_98_147), .B (n_92_148), .C1 (n_88_148), .C2 (n_82_147) );
AOI211_X1 g_104_148 (.ZN (n_104_148), .A (n_100_148), .B (n_94_147), .C1 (n_90_147), .C2 (n_84_148) );
AOI211_X1 g_106_147 (.ZN (n_106_147), .A (n_102_147), .B (n_96_148), .C1 (n_92_148), .C2 (n_86_147) );
AOI211_X1 g_108_148 (.ZN (n_108_148), .A (n_104_148), .B (n_98_147), .C1 (n_94_147), .C2 (n_88_148) );
AOI211_X1 g_110_147 (.ZN (n_110_147), .A (n_106_147), .B (n_100_148), .C1 (n_96_148), .C2 (n_90_147) );
AOI211_X1 g_112_148 (.ZN (n_112_148), .A (n_108_148), .B (n_102_147), .C1 (n_98_147), .C2 (n_92_148) );
AOI211_X1 g_114_147 (.ZN (n_114_147), .A (n_110_147), .B (n_104_148), .C1 (n_100_148), .C2 (n_94_147) );
AOI211_X1 g_116_148 (.ZN (n_116_148), .A (n_112_148), .B (n_106_147), .C1 (n_102_147), .C2 (n_96_148) );
AOI211_X1 g_118_147 (.ZN (n_118_147), .A (n_114_147), .B (n_108_148), .C1 (n_104_148), .C2 (n_98_147) );
AOI211_X1 g_120_148 (.ZN (n_120_148), .A (n_116_148), .B (n_110_147), .C1 (n_106_147), .C2 (n_100_148) );
AOI211_X1 g_122_147 (.ZN (n_122_147), .A (n_118_147), .B (n_112_148), .C1 (n_108_148), .C2 (n_102_147) );
AOI211_X1 g_124_148 (.ZN (n_124_148), .A (n_120_148), .B (n_114_147), .C1 (n_110_147), .C2 (n_104_148) );
AOI211_X1 g_126_147 (.ZN (n_126_147), .A (n_122_147), .B (n_116_148), .C1 (n_112_148), .C2 (n_106_147) );
AOI211_X1 g_128_148 (.ZN (n_128_148), .A (n_124_148), .B (n_118_147), .C1 (n_114_147), .C2 (n_108_148) );
AOI211_X1 g_130_147 (.ZN (n_130_147), .A (n_126_147), .B (n_120_148), .C1 (n_116_148), .C2 (n_110_147) );
AOI211_X1 g_132_148 (.ZN (n_132_148), .A (n_128_148), .B (n_122_147), .C1 (n_118_147), .C2 (n_112_148) );
AOI211_X1 g_134_147 (.ZN (n_134_147), .A (n_130_147), .B (n_124_148), .C1 (n_120_148), .C2 (n_114_147) );
AOI211_X1 g_136_148 (.ZN (n_136_148), .A (n_132_148), .B (n_126_147), .C1 (n_122_147), .C2 (n_116_148) );
AOI211_X1 g_138_147 (.ZN (n_138_147), .A (n_134_147), .B (n_128_148), .C1 (n_124_148), .C2 (n_118_147) );
AOI211_X1 g_140_146 (.ZN (n_140_146), .A (n_136_148), .B (n_130_147), .C1 (n_126_147), .C2 (n_120_148) );
AOI211_X1 g_141_148 (.ZN (n_141_148), .A (n_138_147), .B (n_132_148), .C1 (n_128_148), .C2 (n_122_147) );
AOI211_X1 g_143_147 (.ZN (n_143_147), .A (n_140_146), .B (n_134_147), .C1 (n_130_147), .C2 (n_124_148) );
AOI211_X1 g_145_146 (.ZN (n_145_146), .A (n_141_148), .B (n_136_148), .C1 (n_132_148), .C2 (n_126_147) );
AOI211_X1 g_147_145 (.ZN (n_147_145), .A (n_143_147), .B (n_138_147), .C1 (n_134_147), .C2 (n_128_148) );
AOI211_X1 g_148_143 (.ZN (n_148_143), .A (n_145_146), .B (n_140_146), .C1 (n_136_148), .C2 (n_130_147) );
AOI211_X1 g_149_141 (.ZN (n_149_141), .A (n_147_145), .B (n_141_148), .C1 (n_138_147), .C2 (n_132_148) );
AOI211_X1 g_150_139 (.ZN (n_150_139), .A (n_148_143), .B (n_143_147), .C1 (n_140_146), .C2 (n_134_147) );
AOI211_X1 g_148_138 (.ZN (n_148_138), .A (n_149_141), .B (n_145_146), .C1 (n_141_148), .C2 (n_136_148) );
AOI211_X1 g_147_136 (.ZN (n_147_136), .A (n_150_139), .B (n_147_145), .C1 (n_143_147), .C2 (n_138_147) );
AOI211_X1 g_149_137 (.ZN (n_149_137), .A (n_148_138), .B (n_148_143), .C1 (n_145_146), .C2 (n_140_146) );
AOI211_X1 g_148_139 (.ZN (n_148_139), .A (n_147_136), .B (n_149_141), .C1 (n_147_145), .C2 (n_141_148) );
AOI211_X1 g_147_141 (.ZN (n_147_141), .A (n_149_137), .B (n_150_139), .C1 (n_148_143), .C2 (n_143_147) );
AOI211_X1 g_146_143 (.ZN (n_146_143), .A (n_148_139), .B (n_148_138), .C1 (n_149_141), .C2 (n_145_146) );
AOI211_X1 g_148_142 (.ZN (n_148_142), .A (n_147_141), .B (n_147_136), .C1 (n_150_139), .C2 (n_147_145) );
AOI211_X1 g_147_140 (.ZN (n_147_140), .A (n_146_143), .B (n_149_137), .C1 (n_148_138), .C2 (n_148_143) );
AOI211_X1 g_146_138 (.ZN (n_146_138), .A (n_148_142), .B (n_148_139), .C1 (n_147_136), .C2 (n_149_141) );
AOI211_X1 g_145_140 (.ZN (n_145_140), .A (n_147_140), .B (n_147_141), .C1 (n_149_137), .C2 (n_150_139) );
AOI211_X1 g_146_142 (.ZN (n_146_142), .A (n_146_138), .B (n_146_143), .C1 (n_148_139), .C2 (n_148_138) );
AOI211_X1 g_147_144 (.ZN (n_147_144), .A (n_145_140), .B (n_148_142), .C1 (n_147_141), .C2 (n_147_136) );
AOI211_X1 g_146_146 (.ZN (n_146_146), .A (n_146_142), .B (n_147_140), .C1 (n_146_143), .C2 (n_149_137) );
AOI211_X1 g_145_144 (.ZN (n_145_144), .A (n_147_144), .B (n_146_138), .C1 (n_148_142), .C2 (n_148_139) );
AOI211_X1 g_144_142 (.ZN (n_144_142), .A (n_146_146), .B (n_145_140), .C1 (n_147_140), .C2 (n_147_141) );
AOI211_X1 g_146_141 (.ZN (n_146_141), .A (n_145_144), .B (n_146_142), .C1 (n_146_138), .C2 (n_146_143) );
AOI211_X1 g_148_140 (.ZN (n_148_140), .A (n_144_142), .B (n_147_144), .C1 (n_145_140), .C2 (n_148_142) );
AOI211_X1 g_147_138 (.ZN (n_147_138), .A (n_146_141), .B (n_146_146), .C1 (n_146_142), .C2 (n_147_140) );
AOI211_X1 g_145_139 (.ZN (n_145_139), .A (n_148_140), .B (n_145_144), .C1 (n_147_144), .C2 (n_146_138) );
AOI211_X1 g_144_137 (.ZN (n_144_137), .A (n_147_138), .B (n_144_142), .C1 (n_146_146), .C2 (n_145_140) );
AOI211_X1 g_145_135 (.ZN (n_145_135), .A (n_145_139), .B (n_146_141), .C1 (n_145_144), .C2 (n_146_142) );
AOI211_X1 g_147_134 (.ZN (n_147_134), .A (n_144_137), .B (n_148_140), .C1 (n_144_142), .C2 (n_147_144) );
AOI211_X1 g_149_133 (.ZN (n_149_133), .A (n_145_135), .B (n_147_138), .C1 (n_146_141), .C2 (n_146_146) );
AOI211_X1 g_147_132 (.ZN (n_147_132), .A (n_147_134), .B (n_145_139), .C1 (n_148_140), .C2 (n_145_144) );
AOI211_X1 g_145_131 (.ZN (n_145_131), .A (n_149_133), .B (n_144_137), .C1 (n_147_138), .C2 (n_144_142) );
AOI211_X1 g_147_130 (.ZN (n_147_130), .A (n_147_132), .B (n_145_135), .C1 (n_145_139), .C2 (n_146_141) );
AOI211_X1 g_149_129 (.ZN (n_149_129), .A (n_145_131), .B (n_147_134), .C1 (n_144_137), .C2 (n_148_140) );
AOI211_X1 g_147_128 (.ZN (n_147_128), .A (n_147_130), .B (n_149_133), .C1 (n_145_135), .C2 (n_147_138) );
AOI211_X1 g_145_127 (.ZN (n_145_127), .A (n_149_129), .B (n_147_132), .C1 (n_147_134), .C2 (n_145_139) );
AOI211_X1 g_147_126 (.ZN (n_147_126), .A (n_147_128), .B (n_145_131), .C1 (n_149_133), .C2 (n_144_137) );
AOI211_X1 g_149_125 (.ZN (n_149_125), .A (n_145_127), .B (n_147_130), .C1 (n_147_132), .C2 (n_145_135) );
AOI211_X1 g_147_124 (.ZN (n_147_124), .A (n_147_126), .B (n_149_129), .C1 (n_145_131), .C2 (n_147_134) );
AOI211_X1 g_145_123 (.ZN (n_145_123), .A (n_149_125), .B (n_147_128), .C1 (n_147_130), .C2 (n_149_133) );
AOI211_X1 g_147_122 (.ZN (n_147_122), .A (n_147_124), .B (n_145_127), .C1 (n_149_129), .C2 (n_147_132) );
AOI211_X1 g_149_121 (.ZN (n_149_121), .A (n_145_123), .B (n_147_126), .C1 (n_147_128), .C2 (n_145_131) );
AOI211_X1 g_147_120 (.ZN (n_147_120), .A (n_147_122), .B (n_149_125), .C1 (n_145_127), .C2 (n_147_130) );
AOI211_X1 g_145_119 (.ZN (n_145_119), .A (n_149_121), .B (n_147_124), .C1 (n_147_126), .C2 (n_149_129) );
AOI211_X1 g_147_118 (.ZN (n_147_118), .A (n_147_120), .B (n_145_123), .C1 (n_149_125), .C2 (n_147_128) );
AOI211_X1 g_149_117 (.ZN (n_149_117), .A (n_145_119), .B (n_147_122), .C1 (n_147_124), .C2 (n_145_127) );
AOI211_X1 g_147_116 (.ZN (n_147_116), .A (n_147_118), .B (n_149_121), .C1 (n_145_123), .C2 (n_147_126) );
AOI211_X1 g_145_115 (.ZN (n_145_115), .A (n_149_117), .B (n_147_120), .C1 (n_147_122), .C2 (n_149_125) );
AOI211_X1 g_147_114 (.ZN (n_147_114), .A (n_147_116), .B (n_145_119), .C1 (n_149_121), .C2 (n_147_124) );
AOI211_X1 g_149_113 (.ZN (n_149_113), .A (n_145_115), .B (n_147_118), .C1 (n_147_120), .C2 (n_145_123) );
AOI211_X1 g_147_112 (.ZN (n_147_112), .A (n_147_114), .B (n_149_117), .C1 (n_145_119), .C2 (n_147_122) );
AOI211_X1 g_145_111 (.ZN (n_145_111), .A (n_149_113), .B (n_147_116), .C1 (n_147_118), .C2 (n_149_121) );
AOI211_X1 g_147_110 (.ZN (n_147_110), .A (n_147_112), .B (n_145_115), .C1 (n_149_117), .C2 (n_147_120) );
AOI211_X1 g_149_109 (.ZN (n_149_109), .A (n_145_111), .B (n_147_114), .C1 (n_147_116), .C2 (n_145_119) );
AOI211_X1 g_147_108 (.ZN (n_147_108), .A (n_147_110), .B (n_149_113), .C1 (n_145_115), .C2 (n_147_118) );
AOI211_X1 g_145_107 (.ZN (n_145_107), .A (n_149_109), .B (n_147_112), .C1 (n_147_114), .C2 (n_149_117) );
AOI211_X1 g_147_106 (.ZN (n_147_106), .A (n_147_108), .B (n_145_111), .C1 (n_149_113), .C2 (n_147_116) );
AOI211_X1 g_149_105 (.ZN (n_149_105), .A (n_145_107), .B (n_147_110), .C1 (n_147_112), .C2 (n_145_115) );
AOI211_X1 g_147_104 (.ZN (n_147_104), .A (n_147_106), .B (n_149_109), .C1 (n_145_111), .C2 (n_147_114) );
AOI211_X1 g_145_103 (.ZN (n_145_103), .A (n_149_105), .B (n_147_108), .C1 (n_147_110), .C2 (n_149_113) );
AOI211_X1 g_147_102 (.ZN (n_147_102), .A (n_147_104), .B (n_145_107), .C1 (n_149_109), .C2 (n_147_112) );
AOI211_X1 g_149_101 (.ZN (n_149_101), .A (n_145_103), .B (n_147_106), .C1 (n_147_108), .C2 (n_145_111) );
AOI211_X1 g_147_100 (.ZN (n_147_100), .A (n_147_102), .B (n_149_105), .C1 (n_145_107), .C2 (n_147_110) );
AOI211_X1 g_145_99 (.ZN (n_145_99), .A (n_149_101), .B (n_147_104), .C1 (n_147_106), .C2 (n_149_109) );
AOI211_X1 g_147_98 (.ZN (n_147_98), .A (n_147_100), .B (n_145_103), .C1 (n_149_105), .C2 (n_147_108) );
AOI211_X1 g_149_97 (.ZN (n_149_97), .A (n_145_99), .B (n_147_102), .C1 (n_147_104), .C2 (n_145_107) );
AOI211_X1 g_147_96 (.ZN (n_147_96), .A (n_147_98), .B (n_149_101), .C1 (n_145_103), .C2 (n_147_106) );
AOI211_X1 g_145_95 (.ZN (n_145_95), .A (n_149_97), .B (n_147_100), .C1 (n_147_102), .C2 (n_149_105) );
AOI211_X1 g_147_94 (.ZN (n_147_94), .A (n_147_96), .B (n_145_99), .C1 (n_149_101), .C2 (n_147_104) );
AOI211_X1 g_149_93 (.ZN (n_149_93), .A (n_145_95), .B (n_147_98), .C1 (n_147_100), .C2 (n_145_103) );
AOI211_X1 g_147_92 (.ZN (n_147_92), .A (n_147_94), .B (n_149_97), .C1 (n_145_99), .C2 (n_147_102) );
AOI211_X1 g_145_91 (.ZN (n_145_91), .A (n_149_93), .B (n_147_96), .C1 (n_147_98), .C2 (n_149_101) );
AOI211_X1 g_147_90 (.ZN (n_147_90), .A (n_147_92), .B (n_145_95), .C1 (n_149_97), .C2 (n_147_100) );
AOI211_X1 g_149_89 (.ZN (n_149_89), .A (n_145_91), .B (n_147_94), .C1 (n_147_96), .C2 (n_145_99) );
AOI211_X1 g_147_88 (.ZN (n_147_88), .A (n_147_90), .B (n_149_93), .C1 (n_145_95), .C2 (n_147_98) );
AOI211_X1 g_145_87 (.ZN (n_145_87), .A (n_149_89), .B (n_147_92), .C1 (n_147_94), .C2 (n_149_97) );
AOI211_X1 g_147_86 (.ZN (n_147_86), .A (n_147_88), .B (n_145_91), .C1 (n_149_93), .C2 (n_147_96) );
AOI211_X1 g_149_85 (.ZN (n_149_85), .A (n_145_87), .B (n_147_90), .C1 (n_147_92), .C2 (n_145_95) );
AOI211_X1 g_147_84 (.ZN (n_147_84), .A (n_147_86), .B (n_149_89), .C1 (n_145_91), .C2 (n_147_94) );
AOI211_X1 g_145_83 (.ZN (n_145_83), .A (n_149_85), .B (n_147_88), .C1 (n_147_90), .C2 (n_149_93) );
AOI211_X1 g_147_82 (.ZN (n_147_82), .A (n_147_84), .B (n_145_87), .C1 (n_149_89), .C2 (n_147_92) );
AOI211_X1 g_149_81 (.ZN (n_149_81), .A (n_145_83), .B (n_147_86), .C1 (n_147_88), .C2 (n_145_91) );
AOI211_X1 g_147_80 (.ZN (n_147_80), .A (n_147_82), .B (n_149_85), .C1 (n_145_87), .C2 (n_147_90) );
AOI211_X1 g_145_79 (.ZN (n_145_79), .A (n_149_81), .B (n_147_84), .C1 (n_147_86), .C2 (n_149_89) );
AOI211_X1 g_147_78 (.ZN (n_147_78), .A (n_147_80), .B (n_145_83), .C1 (n_149_85), .C2 (n_147_88) );
AOI211_X1 g_149_77 (.ZN (n_149_77), .A (n_145_79), .B (n_147_82), .C1 (n_147_84), .C2 (n_145_87) );
AOI211_X1 g_148_75 (.ZN (n_148_75), .A (n_147_78), .B (n_149_81), .C1 (n_145_83), .C2 (n_147_86) );
AOI211_X1 g_146_74 (.ZN (n_146_74), .A (n_149_77), .B (n_147_80), .C1 (n_147_82), .C2 (n_149_85) );
AOI211_X1 g_147_76 (.ZN (n_147_76), .A (n_148_75), .B (n_145_79), .C1 (n_149_81), .C2 (n_147_84) );
AOI211_X1 g_145_77 (.ZN (n_145_77), .A (n_146_74), .B (n_147_78), .C1 (n_147_80), .C2 (n_145_83) );
AOI211_X1 g_144_75 (.ZN (n_144_75), .A (n_147_76), .B (n_149_77), .C1 (n_145_79), .C2 (n_147_82) );
AOI211_X1 g_146_76 (.ZN (n_146_76), .A (n_145_77), .B (n_148_75), .C1 (n_147_78), .C2 (n_149_81) );
AOI211_X1 g_144_77 (.ZN (n_144_77), .A (n_144_75), .B (n_146_74), .C1 (n_149_77), .C2 (n_147_80) );
AOI211_X1 g_142_76 (.ZN (n_142_76), .A (n_146_76), .B (n_147_76), .C1 (n_148_75), .C2 (n_145_79) );
AOI211_X1 g_140_77 (.ZN (n_140_77), .A (n_144_77), .B (n_145_77), .C1 (n_146_74), .C2 (n_147_78) );
AOI211_X1 g_138_78 (.ZN (n_138_78), .A (n_142_76), .B (n_144_75), .C1 (n_147_76), .C2 (n_149_77) );
AOI211_X1 g_136_79 (.ZN (n_136_79), .A (n_140_77), .B (n_146_76), .C1 (n_145_77), .C2 (n_148_75) );
AOI211_X1 g_135_81 (.ZN (n_135_81), .A (n_138_78), .B (n_144_77), .C1 (n_144_75), .C2 (n_146_74) );
AOI211_X1 g_134_79 (.ZN (n_134_79), .A (n_136_79), .B (n_142_76), .C1 (n_146_76), .C2 (n_147_76) );
AOI211_X1 g_136_78 (.ZN (n_136_78), .A (n_135_81), .B (n_140_77), .C1 (n_144_77), .C2 (n_145_77) );
AOI211_X1 g_138_77 (.ZN (n_138_77), .A (n_134_79), .B (n_138_78), .C1 (n_142_76), .C2 (n_144_75) );
AOI211_X1 g_140_76 (.ZN (n_140_76), .A (n_136_78), .B (n_136_79), .C1 (n_140_77), .C2 (n_146_76) );
AOI211_X1 g_142_75 (.ZN (n_142_75), .A (n_138_77), .B (n_135_81), .C1 (n_138_78), .C2 (n_144_77) );
AOI211_X1 g_144_76 (.ZN (n_144_76), .A (n_140_76), .B (n_134_79), .C1 (n_136_79), .C2 (n_142_76) );
AOI211_X1 g_142_77 (.ZN (n_142_77), .A (n_142_75), .B (n_136_78), .C1 (n_135_81), .C2 (n_140_77) );
AOI211_X1 g_140_78 (.ZN (n_140_78), .A (n_144_76), .B (n_138_77), .C1 (n_134_79), .C2 (n_138_78) );
AOI211_X1 g_138_79 (.ZN (n_138_79), .A (n_142_77), .B (n_140_76), .C1 (n_136_78), .C2 (n_136_79) );
AOI211_X1 g_139_77 (.ZN (n_139_77), .A (n_140_78), .B (n_142_75), .C1 (n_138_77), .C2 (n_135_81) );
AOI211_X1 g_137_78 (.ZN (n_137_78), .A (n_138_79), .B (n_144_76), .C1 (n_140_76), .C2 (n_134_79) );
AOI211_X1 g_135_79 (.ZN (n_135_79), .A (n_139_77), .B (n_142_77), .C1 (n_142_75), .C2 (n_136_78) );
AOI211_X1 g_133_80 (.ZN (n_133_80), .A (n_137_78), .B (n_140_78), .C1 (n_144_76), .C2 (n_138_77) );
AOI211_X1 g_131_81 (.ZN (n_131_81), .A (n_135_79), .B (n_138_79), .C1 (n_142_77), .C2 (n_140_76) );
AOI211_X1 g_129_82 (.ZN (n_129_82), .A (n_133_80), .B (n_139_77), .C1 (n_140_78), .C2 (n_142_75) );
AOI211_X1 g_127_83 (.ZN (n_127_83), .A (n_131_81), .B (n_137_78), .C1 (n_138_79), .C2 (n_144_76) );
AOI211_X1 g_126_85 (.ZN (n_126_85), .A (n_129_82), .B (n_135_79), .C1 (n_139_77), .C2 (n_142_77) );
AOI211_X1 g_124_84 (.ZN (n_124_84), .A (n_127_83), .B (n_133_80), .C1 (n_137_78), .C2 (n_140_78) );
AOI211_X1 g_126_83 (.ZN (n_126_83), .A (n_126_85), .B (n_131_81), .C1 (n_135_79), .C2 (n_138_79) );
AOI211_X1 g_128_82 (.ZN (n_128_82), .A (n_124_84), .B (n_129_82), .C1 (n_133_80), .C2 (n_139_77) );
AOI211_X1 g_130_81 (.ZN (n_130_81), .A (n_126_83), .B (n_127_83), .C1 (n_131_81), .C2 (n_137_78) );
AOI211_X1 g_132_80 (.ZN (n_132_80), .A (n_128_82), .B (n_126_85), .C1 (n_129_82), .C2 (n_135_79) );
AOI211_X1 g_133_82 (.ZN (n_133_82), .A (n_130_81), .B (n_124_84), .C1 (n_127_83), .C2 (n_133_80) );
AOI211_X1 g_131_83 (.ZN (n_131_83), .A (n_132_80), .B (n_126_83), .C1 (n_126_85), .C2 (n_131_81) );
AOI211_X1 g_129_84 (.ZN (n_129_84), .A (n_133_82), .B (n_128_82), .C1 (n_124_84), .C2 (n_129_82) );
AOI211_X1 g_127_85 (.ZN (n_127_85), .A (n_131_83), .B (n_130_81), .C1 (n_126_83), .C2 (n_127_83) );
AOI211_X1 g_125_86 (.ZN (n_125_86), .A (n_129_84), .B (n_132_80), .C1 (n_128_82), .C2 (n_126_85) );
AOI211_X1 g_123_85 (.ZN (n_123_85), .A (n_127_85), .B (n_133_82), .C1 (n_130_81), .C2 (n_124_84) );
AOI211_X1 g_121_84 (.ZN (n_121_84), .A (n_125_86), .B (n_131_83), .C1 (n_132_80), .C2 (n_126_83) );
AOI211_X1 g_119_85 (.ZN (n_119_85), .A (n_123_85), .B (n_129_84), .C1 (n_133_82), .C2 (n_128_82) );
AOI211_X1 g_117_86 (.ZN (n_117_86), .A (n_121_84), .B (n_127_85), .C1 (n_131_83), .C2 (n_130_81) );
AOI211_X1 g_115_87 (.ZN (n_115_87), .A (n_119_85), .B (n_125_86), .C1 (n_129_84), .C2 (n_132_80) );
AOI211_X1 g_113_88 (.ZN (n_113_88), .A (n_117_86), .B (n_123_85), .C1 (n_127_85), .C2 (n_133_82) );
AOI211_X1 g_111_89 (.ZN (n_111_89), .A (n_115_87), .B (n_121_84), .C1 (n_125_86), .C2 (n_131_83) );
AOI211_X1 g_109_90 (.ZN (n_109_90), .A (n_113_88), .B (n_119_85), .C1 (n_123_85), .C2 (n_129_84) );
AOI211_X1 g_107_91 (.ZN (n_107_91), .A (n_111_89), .B (n_117_86), .C1 (n_121_84), .C2 (n_127_85) );
AOI211_X1 g_105_92 (.ZN (n_105_92), .A (n_109_90), .B (n_115_87), .C1 (n_119_85), .C2 (n_125_86) );
AOI211_X1 g_103_93 (.ZN (n_103_93), .A (n_107_91), .B (n_113_88), .C1 (n_117_86), .C2 (n_123_85) );
AOI211_X1 g_101_94 (.ZN (n_101_94), .A (n_105_92), .B (n_111_89), .C1 (n_115_87), .C2 (n_121_84) );
AOI211_X1 g_99_95 (.ZN (n_99_95), .A (n_103_93), .B (n_109_90), .C1 (n_113_88), .C2 (n_119_85) );
AOI211_X1 g_97_96 (.ZN (n_97_96), .A (n_101_94), .B (n_107_91), .C1 (n_111_89), .C2 (n_117_86) );
AOI211_X1 g_95_97 (.ZN (n_95_97), .A (n_99_95), .B (n_105_92), .C1 (n_109_90), .C2 (n_115_87) );
AOI211_X1 g_93_98 (.ZN (n_93_98), .A (n_97_96), .B (n_103_93), .C1 (n_107_91), .C2 (n_113_88) );
AOI211_X1 g_91_99 (.ZN (n_91_99), .A (n_95_97), .B (n_101_94), .C1 (n_105_92), .C2 (n_111_89) );
AOI211_X1 g_89_100 (.ZN (n_89_100), .A (n_93_98), .B (n_99_95), .C1 (n_103_93), .C2 (n_109_90) );
AOI211_X1 g_90_98 (.ZN (n_90_98), .A (n_91_99), .B (n_97_96), .C1 (n_101_94), .C2 (n_107_91) );
AOI211_X1 g_91_96 (.ZN (n_91_96), .A (n_89_100), .B (n_95_97), .C1 (n_99_95), .C2 (n_105_92) );
AOI211_X1 g_89_97 (.ZN (n_89_97), .A (n_90_98), .B (n_93_98), .C1 (n_97_96), .C2 (n_103_93) );
AOI211_X1 g_87_98 (.ZN (n_87_98), .A (n_91_96), .B (n_91_99), .C1 (n_95_97), .C2 (n_101_94) );
AOI211_X1 g_85_99 (.ZN (n_85_99), .A (n_89_97), .B (n_89_100), .C1 (n_93_98), .C2 (n_99_95) );
AOI211_X1 g_83_100 (.ZN (n_83_100), .A (n_87_98), .B (n_90_98), .C1 (n_91_99), .C2 (n_97_96) );
AOI211_X1 g_81_101 (.ZN (n_81_101), .A (n_85_99), .B (n_91_96), .C1 (n_89_100), .C2 (n_95_97) );
AOI211_X1 g_79_102 (.ZN (n_79_102), .A (n_83_100), .B (n_89_97), .C1 (n_90_98), .C2 (n_93_98) );
AOI211_X1 g_77_103 (.ZN (n_77_103), .A (n_81_101), .B (n_87_98), .C1 (n_91_96), .C2 (n_91_99) );
AOI211_X1 g_78_101 (.ZN (n_78_101), .A (n_79_102), .B (n_85_99), .C1 (n_89_97), .C2 (n_89_100) );
AOI211_X1 g_76_102 (.ZN (n_76_102), .A (n_77_103), .B (n_83_100), .C1 (n_87_98), .C2 (n_90_98) );
AOI211_X1 g_74_103 (.ZN (n_74_103), .A (n_78_101), .B (n_81_101), .C1 (n_85_99), .C2 (n_91_96) );
AOI211_X1 g_72_104 (.ZN (n_72_104), .A (n_76_102), .B (n_79_102), .C1 (n_83_100), .C2 (n_89_97) );
AOI211_X1 g_70_105 (.ZN (n_70_105), .A (n_74_103), .B (n_77_103), .C1 (n_81_101), .C2 (n_87_98) );
AOI211_X1 g_68_106 (.ZN (n_68_106), .A (n_72_104), .B (n_78_101), .C1 (n_79_102), .C2 (n_85_99) );
AOI211_X1 g_66_107 (.ZN (n_66_107), .A (n_70_105), .B (n_76_102), .C1 (n_77_103), .C2 (n_83_100) );
AOI211_X1 g_64_108 (.ZN (n_64_108), .A (n_68_106), .B (n_74_103), .C1 (n_78_101), .C2 (n_81_101) );
AOI211_X1 g_62_109 (.ZN (n_62_109), .A (n_66_107), .B (n_72_104), .C1 (n_76_102), .C2 (n_79_102) );
AOI211_X1 g_60_110 (.ZN (n_60_110), .A (n_64_108), .B (n_70_105), .C1 (n_74_103), .C2 (n_77_103) );
AOI211_X1 g_58_111 (.ZN (n_58_111), .A (n_62_109), .B (n_68_106), .C1 (n_72_104), .C2 (n_78_101) );
AOI211_X1 g_56_112 (.ZN (n_56_112), .A (n_60_110), .B (n_66_107), .C1 (n_70_105), .C2 (n_76_102) );
AOI211_X1 g_54_113 (.ZN (n_54_113), .A (n_58_111), .B (n_64_108), .C1 (n_68_106), .C2 (n_74_103) );
AOI211_X1 g_52_114 (.ZN (n_52_114), .A (n_56_112), .B (n_62_109), .C1 (n_66_107), .C2 (n_72_104) );
AOI211_X1 g_50_115 (.ZN (n_50_115), .A (n_54_113), .B (n_60_110), .C1 (n_64_108), .C2 (n_70_105) );
AOI211_X1 g_48_116 (.ZN (n_48_116), .A (n_52_114), .B (n_58_111), .C1 (n_62_109), .C2 (n_68_106) );
AOI211_X1 g_46_117 (.ZN (n_46_117), .A (n_50_115), .B (n_56_112), .C1 (n_60_110), .C2 (n_66_107) );
AOI211_X1 g_44_118 (.ZN (n_44_118), .A (n_48_116), .B (n_54_113), .C1 (n_58_111), .C2 (n_64_108) );
AOI211_X1 g_42_119 (.ZN (n_42_119), .A (n_46_117), .B (n_52_114), .C1 (n_56_112), .C2 (n_62_109) );
AOI211_X1 g_40_120 (.ZN (n_40_120), .A (n_44_118), .B (n_50_115), .C1 (n_54_113), .C2 (n_60_110) );
AOI211_X1 g_38_121 (.ZN (n_38_121), .A (n_42_119), .B (n_48_116), .C1 (n_52_114), .C2 (n_58_111) );
AOI211_X1 g_36_122 (.ZN (n_36_122), .A (n_40_120), .B (n_46_117), .C1 (n_50_115), .C2 (n_56_112) );
AOI211_X1 g_35_124 (.ZN (n_35_124), .A (n_38_121), .B (n_44_118), .C1 (n_48_116), .C2 (n_54_113) );
AOI211_X1 g_37_123 (.ZN (n_37_123), .A (n_36_122), .B (n_42_119), .C1 (n_46_117), .C2 (n_52_114) );
AOI211_X1 g_39_122 (.ZN (n_39_122), .A (n_35_124), .B (n_40_120), .C1 (n_44_118), .C2 (n_50_115) );
AOI211_X1 g_41_121 (.ZN (n_41_121), .A (n_37_123), .B (n_38_121), .C1 (n_42_119), .C2 (n_48_116) );
AOI211_X1 g_43_120 (.ZN (n_43_120), .A (n_39_122), .B (n_36_122), .C1 (n_40_120), .C2 (n_46_117) );
AOI211_X1 g_45_119 (.ZN (n_45_119), .A (n_41_121), .B (n_35_124), .C1 (n_38_121), .C2 (n_44_118) );
AOI211_X1 g_47_118 (.ZN (n_47_118), .A (n_43_120), .B (n_37_123), .C1 (n_36_122), .C2 (n_42_119) );
AOI211_X1 g_49_117 (.ZN (n_49_117), .A (n_45_119), .B (n_39_122), .C1 (n_35_124), .C2 (n_40_120) );
AOI211_X1 g_51_116 (.ZN (n_51_116), .A (n_47_118), .B (n_41_121), .C1 (n_37_123), .C2 (n_38_121) );
AOI211_X1 g_53_115 (.ZN (n_53_115), .A (n_49_117), .B (n_43_120), .C1 (n_39_122), .C2 (n_36_122) );
AOI211_X1 g_55_114 (.ZN (n_55_114), .A (n_51_116), .B (n_45_119), .C1 (n_41_121), .C2 (n_35_124) );
AOI211_X1 g_57_113 (.ZN (n_57_113), .A (n_53_115), .B (n_47_118), .C1 (n_43_120), .C2 (n_37_123) );
AOI211_X1 g_59_112 (.ZN (n_59_112), .A (n_55_114), .B (n_49_117), .C1 (n_45_119), .C2 (n_39_122) );
AOI211_X1 g_61_111 (.ZN (n_61_111), .A (n_57_113), .B (n_51_116), .C1 (n_47_118), .C2 (n_41_121) );
AOI211_X1 g_63_110 (.ZN (n_63_110), .A (n_59_112), .B (n_53_115), .C1 (n_49_117), .C2 (n_43_120) );
AOI211_X1 g_65_109 (.ZN (n_65_109), .A (n_61_111), .B (n_55_114), .C1 (n_51_116), .C2 (n_45_119) );
AOI211_X1 g_67_108 (.ZN (n_67_108), .A (n_63_110), .B (n_57_113), .C1 (n_53_115), .C2 (n_47_118) );
AOI211_X1 g_69_107 (.ZN (n_69_107), .A (n_65_109), .B (n_59_112), .C1 (n_55_114), .C2 (n_49_117) );
AOI211_X1 g_71_106 (.ZN (n_71_106), .A (n_67_108), .B (n_61_111), .C1 (n_57_113), .C2 (n_51_116) );
AOI211_X1 g_73_105 (.ZN (n_73_105), .A (n_69_107), .B (n_63_110), .C1 (n_59_112), .C2 (n_53_115) );
AOI211_X1 g_75_104 (.ZN (n_75_104), .A (n_71_106), .B (n_65_109), .C1 (n_61_111), .C2 (n_55_114) );
AOI211_X1 g_74_106 (.ZN (n_74_106), .A (n_73_105), .B (n_67_108), .C1 (n_63_110), .C2 (n_57_113) );
AOI211_X1 g_73_104 (.ZN (n_73_104), .A (n_75_104), .B (n_69_107), .C1 (n_65_109), .C2 (n_59_112) );
AOI211_X1 g_75_103 (.ZN (n_75_103), .A (n_74_106), .B (n_71_106), .C1 (n_67_108), .C2 (n_61_111) );
AOI211_X1 g_77_102 (.ZN (n_77_102), .A (n_73_104), .B (n_73_105), .C1 (n_69_107), .C2 (n_63_110) );
AOI211_X1 g_79_101 (.ZN (n_79_101), .A (n_75_103), .B (n_75_104), .C1 (n_71_106), .C2 (n_65_109) );
AOI211_X1 g_81_100 (.ZN (n_81_100), .A (n_77_102), .B (n_74_106), .C1 (n_73_105), .C2 (n_67_108) );
AOI211_X1 g_83_99 (.ZN (n_83_99), .A (n_79_101), .B (n_73_104), .C1 (n_75_104), .C2 (n_69_107) );
AOI211_X1 g_82_101 (.ZN (n_82_101), .A (n_81_100), .B (n_75_103), .C1 (n_74_106), .C2 (n_71_106) );
AOI211_X1 g_84_100 (.ZN (n_84_100), .A (n_83_99), .B (n_77_102), .C1 (n_73_104), .C2 (n_73_105) );
AOI211_X1 g_86_99 (.ZN (n_86_99), .A (n_82_101), .B (n_79_101), .C1 (n_75_103), .C2 (n_75_104) );
AOI211_X1 g_85_101 (.ZN (n_85_101), .A (n_84_100), .B (n_81_100), .C1 (n_77_102), .C2 (n_74_106) );
AOI211_X1 g_87_100 (.ZN (n_87_100), .A (n_86_99), .B (n_83_99), .C1 (n_79_101), .C2 (n_73_104) );
AOI211_X1 g_89_99 (.ZN (n_89_99), .A (n_85_101), .B (n_82_101), .C1 (n_81_100), .C2 (n_75_103) );
AOI211_X1 g_91_98 (.ZN (n_91_98), .A (n_87_100), .B (n_84_100), .C1 (n_83_99), .C2 (n_77_102) );
AOI211_X1 g_93_97 (.ZN (n_93_97), .A (n_89_99), .B (n_86_99), .C1 (n_82_101), .C2 (n_79_101) );
AOI211_X1 g_95_96 (.ZN (n_95_96), .A (n_91_98), .B (n_85_101), .C1 (n_84_100), .C2 (n_81_100) );
AOI211_X1 g_97_95 (.ZN (n_97_95), .A (n_93_97), .B (n_87_100), .C1 (n_86_99), .C2 (n_83_99) );
AOI211_X1 g_99_94 (.ZN (n_99_94), .A (n_95_96), .B (n_89_99), .C1 (n_85_101), .C2 (n_82_101) );
AOI211_X1 g_101_93 (.ZN (n_101_93), .A (n_97_95), .B (n_91_98), .C1 (n_87_100), .C2 (n_84_100) );
AOI211_X1 g_103_92 (.ZN (n_103_92), .A (n_99_94), .B (n_93_97), .C1 (n_89_99), .C2 (n_86_99) );
AOI211_X1 g_105_91 (.ZN (n_105_91), .A (n_101_93), .B (n_95_96), .C1 (n_91_98), .C2 (n_85_101) );
AOI211_X1 g_107_90 (.ZN (n_107_90), .A (n_103_92), .B (n_97_95), .C1 (n_93_97), .C2 (n_87_100) );
AOI211_X1 g_109_89 (.ZN (n_109_89), .A (n_105_91), .B (n_99_94), .C1 (n_95_96), .C2 (n_89_99) );
AOI211_X1 g_108_91 (.ZN (n_108_91), .A (n_107_90), .B (n_101_93), .C1 (n_97_95), .C2 (n_91_98) );
AOI211_X1 g_110_90 (.ZN (n_110_90), .A (n_109_89), .B (n_103_92), .C1 (n_99_94), .C2 (n_93_97) );
AOI211_X1 g_109_92 (.ZN (n_109_92), .A (n_108_91), .B (n_105_91), .C1 (n_101_93), .C2 (n_95_96) );
AOI211_X1 g_111_91 (.ZN (n_111_91), .A (n_110_90), .B (n_107_90), .C1 (n_103_92), .C2 (n_97_95) );
AOI211_X1 g_113_90 (.ZN (n_113_90), .A (n_109_92), .B (n_109_89), .C1 (n_105_91), .C2 (n_99_94) );
AOI211_X1 g_115_89 (.ZN (n_115_89), .A (n_111_91), .B (n_108_91), .C1 (n_107_90), .C2 (n_101_93) );
AOI211_X1 g_117_88 (.ZN (n_117_88), .A (n_113_90), .B (n_110_90), .C1 (n_109_89), .C2 (n_103_92) );
AOI211_X1 g_119_87 (.ZN (n_119_87), .A (n_115_89), .B (n_109_92), .C1 (n_108_91), .C2 (n_105_91) );
AOI211_X1 g_121_86 (.ZN (n_121_86), .A (n_117_88), .B (n_111_91), .C1 (n_110_90), .C2 (n_107_90) );
AOI211_X1 g_120_88 (.ZN (n_120_88), .A (n_119_87), .B (n_113_90), .C1 (n_109_92), .C2 (n_109_89) );
AOI211_X1 g_118_87 (.ZN (n_118_87), .A (n_121_86), .B (n_115_89), .C1 (n_111_91), .C2 (n_108_91) );
AOI211_X1 g_120_86 (.ZN (n_120_86), .A (n_120_88), .B (n_117_88), .C1 (n_113_90), .C2 (n_110_90) );
AOI211_X1 g_122_85 (.ZN (n_122_85), .A (n_118_87), .B (n_119_87), .C1 (n_115_89), .C2 (n_109_92) );
AOI211_X1 g_124_86 (.ZN (n_124_86), .A (n_120_86), .B (n_121_86), .C1 (n_117_88), .C2 (n_111_91) );
AOI211_X1 g_122_87 (.ZN (n_122_87), .A (n_122_85), .B (n_120_88), .C1 (n_119_87), .C2 (n_113_90) );
AOI211_X1 g_124_88 (.ZN (n_124_88), .A (n_124_86), .B (n_118_87), .C1 (n_121_86), .C2 (n_115_89) );
AOI211_X1 g_123_86 (.ZN (n_123_86), .A (n_122_87), .B (n_120_86), .C1 (n_120_88), .C2 (n_117_88) );
AOI211_X1 g_125_85 (.ZN (n_125_85), .A (n_124_88), .B (n_122_85), .C1 (n_118_87), .C2 (n_119_87) );
AOI211_X1 g_127_84 (.ZN (n_127_84), .A (n_123_86), .B (n_124_86), .C1 (n_120_86), .C2 (n_121_86) );
AOI211_X1 g_129_83 (.ZN (n_129_83), .A (n_125_85), .B (n_122_87), .C1 (n_122_85), .C2 (n_120_88) );
AOI211_X1 g_131_82 (.ZN (n_131_82), .A (n_127_84), .B (n_124_88), .C1 (n_124_86), .C2 (n_118_87) );
AOI211_X1 g_133_81 (.ZN (n_133_81), .A (n_129_83), .B (n_123_86), .C1 (n_122_87), .C2 (n_120_86) );
AOI211_X1 g_135_80 (.ZN (n_135_80), .A (n_131_82), .B (n_125_85), .C1 (n_124_88), .C2 (n_122_85) );
AOI211_X1 g_137_79 (.ZN (n_137_79), .A (n_133_81), .B (n_127_84), .C1 (n_123_86), .C2 (n_124_86) );
AOI211_X1 g_139_78 (.ZN (n_139_78), .A (n_135_80), .B (n_129_83), .C1 (n_125_85), .C2 (n_122_87) );
AOI211_X1 g_141_77 (.ZN (n_141_77), .A (n_137_79), .B (n_131_82), .C1 (n_127_84), .C2 (n_124_88) );
AOI211_X1 g_143_76 (.ZN (n_143_76), .A (n_139_78), .B (n_133_81), .C1 (n_129_83), .C2 (n_123_86) );
AOI211_X1 g_142_78 (.ZN (n_142_78), .A (n_141_77), .B (n_135_80), .C1 (n_131_82), .C2 (n_125_85) );
AOI211_X1 g_140_79 (.ZN (n_140_79), .A (n_143_76), .B (n_137_79), .C1 (n_133_81), .C2 (n_127_84) );
AOI211_X1 g_138_80 (.ZN (n_138_80), .A (n_142_78), .B (n_139_78), .C1 (n_135_80), .C2 (n_129_83) );
AOI211_X1 g_136_81 (.ZN (n_136_81), .A (n_140_79), .B (n_141_77), .C1 (n_137_79), .C2 (n_131_82) );
AOI211_X1 g_134_82 (.ZN (n_134_82), .A (n_138_80), .B (n_143_76), .C1 (n_139_78), .C2 (n_133_81) );
AOI211_X1 g_132_83 (.ZN (n_132_83), .A (n_136_81), .B (n_142_78), .C1 (n_141_77), .C2 (n_135_80) );
AOI211_X1 g_130_84 (.ZN (n_130_84), .A (n_134_82), .B (n_140_79), .C1 (n_143_76), .C2 (n_137_79) );
AOI211_X1 g_128_85 (.ZN (n_128_85), .A (n_132_83), .B (n_138_80), .C1 (n_142_78), .C2 (n_139_78) );
AOI211_X1 g_126_86 (.ZN (n_126_86), .A (n_130_84), .B (n_136_81), .C1 (n_140_79), .C2 (n_141_77) );
AOI211_X1 g_124_85 (.ZN (n_124_85), .A (n_128_85), .B (n_134_82), .C1 (n_138_80), .C2 (n_143_76) );
AOI211_X1 g_122_86 (.ZN (n_122_86), .A (n_126_86), .B (n_132_83), .C1 (n_136_81), .C2 (n_142_78) );
AOI211_X1 g_120_87 (.ZN (n_120_87), .A (n_124_85), .B (n_130_84), .C1 (n_134_82), .C2 (n_140_79) );
AOI211_X1 g_118_88 (.ZN (n_118_88), .A (n_122_86), .B (n_128_85), .C1 (n_132_83), .C2 (n_138_80) );
AOI211_X1 g_116_89 (.ZN (n_116_89), .A (n_120_87), .B (n_126_86), .C1 (n_130_84), .C2 (n_136_81) );
AOI211_X1 g_114_90 (.ZN (n_114_90), .A (n_118_88), .B (n_124_85), .C1 (n_128_85), .C2 (n_134_82) );
AOI211_X1 g_115_88 (.ZN (n_115_88), .A (n_116_89), .B (n_122_86), .C1 (n_126_86), .C2 (n_132_83) );
AOI211_X1 g_113_89 (.ZN (n_113_89), .A (n_114_90), .B (n_120_87), .C1 (n_124_85), .C2 (n_130_84) );
AOI211_X1 g_111_90 (.ZN (n_111_90), .A (n_115_88), .B (n_118_88), .C1 (n_122_86), .C2 (n_128_85) );
AOI211_X1 g_109_91 (.ZN (n_109_91), .A (n_113_89), .B (n_116_89), .C1 (n_120_87), .C2 (n_126_86) );
AOI211_X1 g_107_92 (.ZN (n_107_92), .A (n_111_90), .B (n_114_90), .C1 (n_118_88), .C2 (n_124_85) );
AOI211_X1 g_105_93 (.ZN (n_105_93), .A (n_109_91), .B (n_115_88), .C1 (n_116_89), .C2 (n_122_86) );
AOI211_X1 g_103_94 (.ZN (n_103_94), .A (n_107_92), .B (n_113_89), .C1 (n_114_90), .C2 (n_120_87) );
AOI211_X1 g_104_92 (.ZN (n_104_92), .A (n_105_93), .B (n_111_90), .C1 (n_115_88), .C2 (n_118_88) );
AOI211_X1 g_102_93 (.ZN (n_102_93), .A (n_103_94), .B (n_109_91), .C1 (n_113_89), .C2 (n_116_89) );
AOI211_X1 g_100_94 (.ZN (n_100_94), .A (n_104_92), .B (n_107_92), .C1 (n_111_90), .C2 (n_114_90) );
AOI211_X1 g_98_95 (.ZN (n_98_95), .A (n_102_93), .B (n_105_93), .C1 (n_109_91), .C2 (n_115_88) );
AOI211_X1 g_96_96 (.ZN (n_96_96), .A (n_100_94), .B (n_103_94), .C1 (n_107_92), .C2 (n_113_89) );
AOI211_X1 g_94_97 (.ZN (n_94_97), .A (n_98_95), .B (n_104_92), .C1 (n_105_93), .C2 (n_111_90) );
AOI211_X1 g_92_98 (.ZN (n_92_98), .A (n_96_96), .B (n_102_93), .C1 (n_103_94), .C2 (n_109_91) );
AOI211_X1 g_90_99 (.ZN (n_90_99), .A (n_94_97), .B (n_100_94), .C1 (n_104_92), .C2 (n_107_92) );
AOI211_X1 g_88_100 (.ZN (n_88_100), .A (n_92_98), .B (n_98_95), .C1 (n_102_93), .C2 (n_105_93) );
AOI211_X1 g_86_101 (.ZN (n_86_101), .A (n_90_99), .B (n_96_96), .C1 (n_100_94), .C2 (n_103_94) );
AOI211_X1 g_84_102 (.ZN (n_84_102), .A (n_88_100), .B (n_94_97), .C1 (n_98_95), .C2 (n_104_92) );
AOI211_X1 g_82_103 (.ZN (n_82_103), .A (n_86_101), .B (n_92_98), .C1 (n_96_96), .C2 (n_102_93) );
AOI211_X1 g_83_101 (.ZN (n_83_101), .A (n_84_102), .B (n_90_99), .C1 (n_94_97), .C2 (n_100_94) );
AOI211_X1 g_81_102 (.ZN (n_81_102), .A (n_82_103), .B (n_88_100), .C1 (n_92_98), .C2 (n_98_95) );
AOI211_X1 g_82_100 (.ZN (n_82_100), .A (n_83_101), .B (n_86_101), .C1 (n_90_99), .C2 (n_96_96) );
AOI211_X1 g_80_101 (.ZN (n_80_101), .A (n_81_102), .B (n_84_102), .C1 (n_88_100), .C2 (n_94_97) );
AOI211_X1 g_78_102 (.ZN (n_78_102), .A (n_82_100), .B (n_82_103), .C1 (n_86_101), .C2 (n_92_98) );
AOI211_X1 g_76_103 (.ZN (n_76_103), .A (n_80_101), .B (n_83_101), .C1 (n_84_102), .C2 (n_90_99) );
AOI211_X1 g_74_104 (.ZN (n_74_104), .A (n_78_102), .B (n_81_102), .C1 (n_82_103), .C2 (n_88_100) );
AOI211_X1 g_72_105 (.ZN (n_72_105), .A (n_76_103), .B (n_82_100), .C1 (n_83_101), .C2 (n_86_101) );
AOI211_X1 g_70_106 (.ZN (n_70_106), .A (n_74_104), .B (n_80_101), .C1 (n_81_102), .C2 (n_84_102) );
AOI211_X1 g_68_107 (.ZN (n_68_107), .A (n_72_105), .B (n_78_102), .C1 (n_82_100), .C2 (n_82_103) );
AOI211_X1 g_67_109 (.ZN (n_67_109), .A (n_70_106), .B (n_76_103), .C1 (n_80_101), .C2 (n_83_101) );
AOI211_X1 g_65_108 (.ZN (n_65_108), .A (n_68_107), .B (n_74_104), .C1 (n_78_102), .C2 (n_81_102) );
AOI211_X1 g_67_107 (.ZN (n_67_107), .A (n_67_109), .B (n_72_105), .C1 (n_76_103), .C2 (n_82_100) );
AOI211_X1 g_69_106 (.ZN (n_69_106), .A (n_65_108), .B (n_70_106), .C1 (n_74_104), .C2 (n_80_101) );
AOI211_X1 g_71_105 (.ZN (n_71_105), .A (n_67_107), .B (n_68_107), .C1 (n_72_105), .C2 (n_78_102) );
AOI211_X1 g_72_107 (.ZN (n_72_107), .A (n_69_106), .B (n_67_109), .C1 (n_70_106), .C2 (n_76_103) );
AOI211_X1 g_70_108 (.ZN (n_70_108), .A (n_71_105), .B (n_65_108), .C1 (n_68_107), .C2 (n_74_104) );
AOI211_X1 g_68_109 (.ZN (n_68_109), .A (n_72_107), .B (n_67_107), .C1 (n_67_109), .C2 (n_72_105) );
AOI211_X1 g_66_110 (.ZN (n_66_110), .A (n_70_108), .B (n_69_106), .C1 (n_65_108), .C2 (n_70_106) );
AOI211_X1 g_64_111 (.ZN (n_64_111), .A (n_68_109), .B (n_71_105), .C1 (n_67_107), .C2 (n_68_107) );
AOI211_X1 g_63_109 (.ZN (n_63_109), .A (n_66_110), .B (n_72_107), .C1 (n_69_106), .C2 (n_67_109) );
AOI211_X1 g_61_110 (.ZN (n_61_110), .A (n_64_111), .B (n_70_108), .C1 (n_71_105), .C2 (n_65_108) );
AOI211_X1 g_59_111 (.ZN (n_59_111), .A (n_63_109), .B (n_68_109), .C1 (n_72_107), .C2 (n_67_107) );
AOI211_X1 g_57_112 (.ZN (n_57_112), .A (n_61_110), .B (n_66_110), .C1 (n_70_108), .C2 (n_69_106) );
AOI211_X1 g_55_113 (.ZN (n_55_113), .A (n_59_111), .B (n_64_111), .C1 (n_68_109), .C2 (n_71_105) );
AOI211_X1 g_53_114 (.ZN (n_53_114), .A (n_57_112), .B (n_63_109), .C1 (n_66_110), .C2 (n_72_107) );
AOI211_X1 g_51_115 (.ZN (n_51_115), .A (n_55_113), .B (n_61_110), .C1 (n_64_111), .C2 (n_70_108) );
AOI211_X1 g_49_116 (.ZN (n_49_116), .A (n_53_114), .B (n_59_111), .C1 (n_63_109), .C2 (n_68_109) );
AOI211_X1 g_47_117 (.ZN (n_47_117), .A (n_51_115), .B (n_57_112), .C1 (n_61_110), .C2 (n_66_110) );
AOI211_X1 g_45_118 (.ZN (n_45_118), .A (n_49_116), .B (n_55_113), .C1 (n_59_111), .C2 (n_64_111) );
AOI211_X1 g_43_119 (.ZN (n_43_119), .A (n_47_117), .B (n_53_114), .C1 (n_57_112), .C2 (n_63_109) );
AOI211_X1 g_41_120 (.ZN (n_41_120), .A (n_45_118), .B (n_51_115), .C1 (n_55_113), .C2 (n_61_110) );
AOI211_X1 g_39_121 (.ZN (n_39_121), .A (n_43_119), .B (n_49_116), .C1 (n_53_114), .C2 (n_59_111) );
AOI211_X1 g_37_122 (.ZN (n_37_122), .A (n_41_120), .B (n_47_117), .C1 (n_51_115), .C2 (n_57_112) );
AOI211_X1 g_35_123 (.ZN (n_35_123), .A (n_39_121), .B (n_45_118), .C1 (n_49_116), .C2 (n_55_113) );
AOI211_X1 g_33_124 (.ZN (n_33_124), .A (n_37_122), .B (n_43_119), .C1 (n_47_117), .C2 (n_53_114) );
AOI211_X1 g_31_125 (.ZN (n_31_125), .A (n_35_123), .B (n_41_120), .C1 (n_45_118), .C2 (n_51_115) );
AOI211_X1 g_29_126 (.ZN (n_29_126), .A (n_33_124), .B (n_39_121), .C1 (n_43_119), .C2 (n_49_116) );
AOI211_X1 g_27_127 (.ZN (n_27_127), .A (n_31_125), .B (n_37_122), .C1 (n_41_120), .C2 (n_47_117) );
AOI211_X1 g_25_128 (.ZN (n_25_128), .A (n_29_126), .B (n_35_123), .C1 (n_39_121), .C2 (n_45_118) );
AOI211_X1 g_23_129 (.ZN (n_23_129), .A (n_27_127), .B (n_33_124), .C1 (n_37_122), .C2 (n_43_119) );
AOI211_X1 g_21_130 (.ZN (n_21_130), .A (n_25_128), .B (n_31_125), .C1 (n_35_123), .C2 (n_41_120) );
AOI211_X1 g_19_131 (.ZN (n_19_131), .A (n_23_129), .B (n_29_126), .C1 (n_33_124), .C2 (n_39_121) );
AOI211_X1 g_17_132 (.ZN (n_17_132), .A (n_21_130), .B (n_27_127), .C1 (n_31_125), .C2 (n_37_122) );
AOI211_X1 g_19_133 (.ZN (n_19_133), .A (n_19_131), .B (n_25_128), .C1 (n_29_126), .C2 (n_35_123) );
AOI211_X1 g_21_132 (.ZN (n_21_132), .A (n_17_132), .B (n_23_129), .C1 (n_27_127), .C2 (n_33_124) );
AOI211_X1 g_23_131 (.ZN (n_23_131), .A (n_19_133), .B (n_21_130), .C1 (n_25_128), .C2 (n_31_125) );
AOI211_X1 g_25_130 (.ZN (n_25_130), .A (n_21_132), .B (n_19_131), .C1 (n_23_129), .C2 (n_29_126) );
AOI211_X1 g_27_129 (.ZN (n_27_129), .A (n_23_131), .B (n_17_132), .C1 (n_21_130), .C2 (n_27_127) );
AOI211_X1 g_29_128 (.ZN (n_29_128), .A (n_25_130), .B (n_19_133), .C1 (n_19_131), .C2 (n_25_128) );
AOI211_X1 g_31_127 (.ZN (n_31_127), .A (n_27_129), .B (n_21_132), .C1 (n_17_132), .C2 (n_23_129) );
AOI211_X1 g_33_126 (.ZN (n_33_126), .A (n_29_128), .B (n_23_131), .C1 (n_19_133), .C2 (n_21_130) );
AOI211_X1 g_35_125 (.ZN (n_35_125), .A (n_31_127), .B (n_25_130), .C1 (n_21_132), .C2 (n_19_131) );
AOI211_X1 g_37_124 (.ZN (n_37_124), .A (n_33_126), .B (n_27_129), .C1 (n_23_131), .C2 (n_17_132) );
AOI211_X1 g_39_123 (.ZN (n_39_123), .A (n_35_125), .B (n_29_128), .C1 (n_25_130), .C2 (n_19_133) );
AOI211_X1 g_41_122 (.ZN (n_41_122), .A (n_37_124), .B (n_31_127), .C1 (n_27_129), .C2 (n_21_132) );
AOI211_X1 g_43_121 (.ZN (n_43_121), .A (n_39_123), .B (n_33_126), .C1 (n_29_128), .C2 (n_23_131) );
AOI211_X1 g_45_120 (.ZN (n_45_120), .A (n_41_122), .B (n_35_125), .C1 (n_31_127), .C2 (n_25_130) );
AOI211_X1 g_47_119 (.ZN (n_47_119), .A (n_43_121), .B (n_37_124), .C1 (n_33_126), .C2 (n_27_129) );
AOI211_X1 g_49_118 (.ZN (n_49_118), .A (n_45_120), .B (n_39_123), .C1 (n_35_125), .C2 (n_29_128) );
AOI211_X1 g_51_117 (.ZN (n_51_117), .A (n_47_119), .B (n_41_122), .C1 (n_37_124), .C2 (n_31_127) );
AOI211_X1 g_53_116 (.ZN (n_53_116), .A (n_49_118), .B (n_43_121), .C1 (n_39_123), .C2 (n_33_126) );
AOI211_X1 g_55_115 (.ZN (n_55_115), .A (n_51_117), .B (n_45_120), .C1 (n_41_122), .C2 (n_35_125) );
AOI211_X1 g_57_114 (.ZN (n_57_114), .A (n_53_116), .B (n_47_119), .C1 (n_43_121), .C2 (n_37_124) );
AOI211_X1 g_59_113 (.ZN (n_59_113), .A (n_55_115), .B (n_49_118), .C1 (n_45_120), .C2 (n_39_123) );
AOI211_X1 g_61_112 (.ZN (n_61_112), .A (n_57_114), .B (n_51_117), .C1 (n_47_119), .C2 (n_41_122) );
AOI211_X1 g_63_111 (.ZN (n_63_111), .A (n_59_113), .B (n_53_116), .C1 (n_49_118), .C2 (n_43_121) );
AOI211_X1 g_65_110 (.ZN (n_65_110), .A (n_61_112), .B (n_55_115), .C1 (n_51_117), .C2 (n_45_120) );
AOI211_X1 g_64_112 (.ZN (n_64_112), .A (n_63_111), .B (n_57_114), .C1 (n_53_116), .C2 (n_47_119) );
AOI211_X1 g_62_111 (.ZN (n_62_111), .A (n_65_110), .B (n_59_113), .C1 (n_55_115), .C2 (n_49_118) );
AOI211_X1 g_64_110 (.ZN (n_64_110), .A (n_64_112), .B (n_61_112), .C1 (n_57_114), .C2 (n_51_117) );
AOI211_X1 g_66_109 (.ZN (n_66_109), .A (n_62_111), .B (n_63_111), .C1 (n_59_113), .C2 (n_53_116) );
AOI211_X1 g_68_108 (.ZN (n_68_108), .A (n_64_110), .B (n_65_110), .C1 (n_61_112), .C2 (n_55_115) );
AOI211_X1 g_70_107 (.ZN (n_70_107), .A (n_66_109), .B (n_64_112), .C1 (n_63_111), .C2 (n_57_114) );
AOI211_X1 g_72_106 (.ZN (n_72_106), .A (n_68_108), .B (n_62_111), .C1 (n_65_110), .C2 (n_59_113) );
AOI211_X1 g_74_105 (.ZN (n_74_105), .A (n_70_107), .B (n_64_110), .C1 (n_64_112), .C2 (n_61_112) );
AOI211_X1 g_76_104 (.ZN (n_76_104), .A (n_72_106), .B (n_66_109), .C1 (n_62_111), .C2 (n_63_111) );
AOI211_X1 g_78_103 (.ZN (n_78_103), .A (n_74_105), .B (n_68_108), .C1 (n_64_110), .C2 (n_65_110) );
AOI211_X1 g_80_102 (.ZN (n_80_102), .A (n_76_104), .B (n_70_107), .C1 (n_66_109), .C2 (n_64_112) );
AOI211_X1 g_79_104 (.ZN (n_79_104), .A (n_78_103), .B (n_72_106), .C1 (n_68_108), .C2 (n_62_111) );
AOI211_X1 g_81_103 (.ZN (n_81_103), .A (n_80_102), .B (n_74_105), .C1 (n_70_107), .C2 (n_64_110) );
AOI211_X1 g_83_102 (.ZN (n_83_102), .A (n_79_104), .B (n_76_104), .C1 (n_72_106), .C2 (n_66_109) );
AOI211_X1 g_82_104 (.ZN (n_82_104), .A (n_81_103), .B (n_78_103), .C1 (n_74_105), .C2 (n_68_108) );
AOI211_X1 g_80_103 (.ZN (n_80_103), .A (n_83_102), .B (n_80_102), .C1 (n_76_104), .C2 (n_70_107) );
AOI211_X1 g_82_102 (.ZN (n_82_102), .A (n_82_104), .B (n_79_104), .C1 (n_78_103), .C2 (n_72_106) );
AOI211_X1 g_84_101 (.ZN (n_84_101), .A (n_80_103), .B (n_81_103), .C1 (n_80_102), .C2 (n_74_105) );
AOI211_X1 g_86_100 (.ZN (n_86_100), .A (n_82_102), .B (n_83_102), .C1 (n_79_104), .C2 (n_76_104) );
AOI211_X1 g_88_99 (.ZN (n_88_99), .A (n_84_101), .B (n_82_104), .C1 (n_81_103), .C2 (n_78_103) );
AOI211_X1 g_87_101 (.ZN (n_87_101), .A (n_86_100), .B (n_80_103), .C1 (n_83_102), .C2 (n_80_102) );
AOI211_X1 g_85_102 (.ZN (n_85_102), .A (n_88_99), .B (n_82_102), .C1 (n_82_104), .C2 (n_79_104) );
AOI211_X1 g_83_103 (.ZN (n_83_103), .A (n_87_101), .B (n_84_101), .C1 (n_80_103), .C2 (n_81_103) );
AOI211_X1 g_81_104 (.ZN (n_81_104), .A (n_85_102), .B (n_86_100), .C1 (n_82_102), .C2 (n_83_102) );
AOI211_X1 g_79_103 (.ZN (n_79_103), .A (n_83_103), .B (n_88_99), .C1 (n_84_101), .C2 (n_82_104) );
AOI211_X1 g_77_104 (.ZN (n_77_104), .A (n_81_104), .B (n_87_101), .C1 (n_86_100), .C2 (n_80_103) );
AOI211_X1 g_75_105 (.ZN (n_75_105), .A (n_79_103), .B (n_85_102), .C1 (n_88_99), .C2 (n_82_102) );
AOI211_X1 g_73_106 (.ZN (n_73_106), .A (n_77_104), .B (n_83_103), .C1 (n_87_101), .C2 (n_84_101) );
AOI211_X1 g_71_107 (.ZN (n_71_107), .A (n_75_105), .B (n_81_104), .C1 (n_85_102), .C2 (n_86_100) );
AOI211_X1 g_69_108 (.ZN (n_69_108), .A (n_73_106), .B (n_79_103), .C1 (n_83_103), .C2 (n_88_99) );
AOI211_X1 g_68_110 (.ZN (n_68_110), .A (n_71_107), .B (n_77_104), .C1 (n_81_104), .C2 (n_87_101) );
AOI211_X1 g_66_111 (.ZN (n_66_111), .A (n_69_108), .B (n_75_105), .C1 (n_79_103), .C2 (n_85_102) );
AOI211_X1 g_65_113 (.ZN (n_65_113), .A (n_68_110), .B (n_73_106), .C1 (n_77_104), .C2 (n_83_103) );
AOI211_X1 g_63_112 (.ZN (n_63_112), .A (n_66_111), .B (n_71_107), .C1 (n_75_105), .C2 (n_81_104) );
AOI211_X1 g_65_111 (.ZN (n_65_111), .A (n_65_113), .B (n_69_108), .C1 (n_73_106), .C2 (n_79_103) );
AOI211_X1 g_67_110 (.ZN (n_67_110), .A (n_63_112), .B (n_68_110), .C1 (n_71_107), .C2 (n_77_104) );
AOI211_X1 g_69_109 (.ZN (n_69_109), .A (n_65_111), .B (n_66_111), .C1 (n_69_108), .C2 (n_75_105) );
AOI211_X1 g_71_108 (.ZN (n_71_108), .A (n_67_110), .B (n_65_113), .C1 (n_68_110), .C2 (n_73_106) );
AOI211_X1 g_73_107 (.ZN (n_73_107), .A (n_69_109), .B (n_63_112), .C1 (n_66_111), .C2 (n_71_107) );
AOI211_X1 g_75_106 (.ZN (n_75_106), .A (n_71_108), .B (n_65_111), .C1 (n_65_113), .C2 (n_69_108) );
AOI211_X1 g_77_105 (.ZN (n_77_105), .A (n_73_107), .B (n_67_110), .C1 (n_63_112), .C2 (n_68_110) );
AOI211_X1 g_76_107 (.ZN (n_76_107), .A (n_75_106), .B (n_69_109), .C1 (n_65_111), .C2 (n_66_111) );
AOI211_X1 g_74_108 (.ZN (n_74_108), .A (n_77_105), .B (n_71_108), .C1 (n_67_110), .C2 (n_65_113) );
AOI211_X1 g_72_109 (.ZN (n_72_109), .A (n_76_107), .B (n_73_107), .C1 (n_69_109), .C2 (n_63_112) );
AOI211_X1 g_70_110 (.ZN (n_70_110), .A (n_74_108), .B (n_75_106), .C1 (n_71_108), .C2 (n_65_111) );
AOI211_X1 g_68_111 (.ZN (n_68_111), .A (n_72_109), .B (n_77_105), .C1 (n_73_107), .C2 (n_67_110) );
AOI211_X1 g_66_112 (.ZN (n_66_112), .A (n_70_110), .B (n_76_107), .C1 (n_75_106), .C2 (n_69_109) );
AOI211_X1 g_64_113 (.ZN (n_64_113), .A (n_68_111), .B (n_74_108), .C1 (n_77_105), .C2 (n_71_108) );
AOI211_X1 g_62_112 (.ZN (n_62_112), .A (n_66_112), .B (n_72_109), .C1 (n_76_107), .C2 (n_73_107) );
AOI211_X1 g_60_113 (.ZN (n_60_113), .A (n_64_113), .B (n_70_110), .C1 (n_74_108), .C2 (n_75_106) );
AOI211_X1 g_58_114 (.ZN (n_58_114), .A (n_62_112), .B (n_68_111), .C1 (n_72_109), .C2 (n_77_105) );
AOI211_X1 g_56_115 (.ZN (n_56_115), .A (n_60_113), .B (n_66_112), .C1 (n_70_110), .C2 (n_76_107) );
AOI211_X1 g_54_116 (.ZN (n_54_116), .A (n_58_114), .B (n_64_113), .C1 (n_68_111), .C2 (n_74_108) );
AOI211_X1 g_52_117 (.ZN (n_52_117), .A (n_56_115), .B (n_62_112), .C1 (n_66_112), .C2 (n_72_109) );
AOI211_X1 g_50_118 (.ZN (n_50_118), .A (n_54_116), .B (n_60_113), .C1 (n_64_113), .C2 (n_70_110) );
AOI211_X1 g_48_119 (.ZN (n_48_119), .A (n_52_117), .B (n_58_114), .C1 (n_62_112), .C2 (n_68_111) );
AOI211_X1 g_46_120 (.ZN (n_46_120), .A (n_50_118), .B (n_56_115), .C1 (n_60_113), .C2 (n_66_112) );
AOI211_X1 g_44_121 (.ZN (n_44_121), .A (n_48_119), .B (n_54_116), .C1 (n_58_114), .C2 (n_64_113) );
AOI211_X1 g_42_122 (.ZN (n_42_122), .A (n_46_120), .B (n_52_117), .C1 (n_56_115), .C2 (n_62_112) );
AOI211_X1 g_40_123 (.ZN (n_40_123), .A (n_44_121), .B (n_50_118), .C1 (n_54_116), .C2 (n_60_113) );
AOI211_X1 g_38_124 (.ZN (n_38_124), .A (n_42_122), .B (n_48_119), .C1 (n_52_117), .C2 (n_58_114) );
AOI211_X1 g_36_125 (.ZN (n_36_125), .A (n_40_123), .B (n_46_120), .C1 (n_50_118), .C2 (n_56_115) );
AOI211_X1 g_34_126 (.ZN (n_34_126), .A (n_38_124), .B (n_44_121), .C1 (n_48_119), .C2 (n_54_116) );
AOI211_X1 g_32_127 (.ZN (n_32_127), .A (n_36_125), .B (n_42_122), .C1 (n_46_120), .C2 (n_52_117) );
AOI211_X1 g_33_125 (.ZN (n_33_125), .A (n_34_126), .B (n_40_123), .C1 (n_44_121), .C2 (n_50_118) );
AOI211_X1 g_31_126 (.ZN (n_31_126), .A (n_32_127), .B (n_38_124), .C1 (n_42_122), .C2 (n_48_119) );
AOI211_X1 g_29_127 (.ZN (n_29_127), .A (n_33_125), .B (n_36_125), .C1 (n_40_123), .C2 (n_46_120) );
AOI211_X1 g_27_128 (.ZN (n_27_128), .A (n_31_126), .B (n_34_126), .C1 (n_38_124), .C2 (n_44_121) );
AOI211_X1 g_25_129 (.ZN (n_25_129), .A (n_29_127), .B (n_32_127), .C1 (n_36_125), .C2 (n_42_122) );
AOI211_X1 g_23_130 (.ZN (n_23_130), .A (n_27_128), .B (n_33_125), .C1 (n_34_126), .C2 (n_40_123) );
AOI211_X1 g_21_131 (.ZN (n_21_131), .A (n_25_129), .B (n_31_126), .C1 (n_32_127), .C2 (n_38_124) );
AOI211_X1 g_19_132 (.ZN (n_19_132), .A (n_23_130), .B (n_29_127), .C1 (n_33_125), .C2 (n_36_125) );
AOI211_X1 g_17_133 (.ZN (n_17_133), .A (n_21_131), .B (n_27_128), .C1 (n_31_126), .C2 (n_34_126) );
AOI211_X1 g_15_134 (.ZN (n_15_134), .A (n_19_132), .B (n_25_129), .C1 (n_29_127), .C2 (n_32_127) );
AOI211_X1 g_13_135 (.ZN (n_13_135), .A (n_17_133), .B (n_23_130), .C1 (n_27_128), .C2 (n_33_125) );
AOI211_X1 g_11_136 (.ZN (n_11_136), .A (n_15_134), .B (n_21_131), .C1 (n_25_129), .C2 (n_31_126) );
AOI211_X1 g_9_137 (.ZN (n_9_137), .A (n_13_135), .B (n_19_132), .C1 (n_23_130), .C2 (n_29_127) );
AOI211_X1 g_7_138 (.ZN (n_7_138), .A (n_11_136), .B (n_17_133), .C1 (n_21_131), .C2 (n_27_128) );
AOI211_X1 g_6_140 (.ZN (n_6_140), .A (n_9_137), .B (n_15_134), .C1 (n_19_132), .C2 (n_25_129) );
AOI211_X1 g_8_139 (.ZN (n_8_139), .A (n_7_138), .B (n_13_135), .C1 (n_17_133), .C2 (n_23_130) );
AOI211_X1 g_10_138 (.ZN (n_10_138), .A (n_6_140), .B (n_11_136), .C1 (n_15_134), .C2 (n_21_131) );
AOI211_X1 g_12_137 (.ZN (n_12_137), .A (n_8_139), .B (n_9_137), .C1 (n_13_135), .C2 (n_19_132) );
AOI211_X1 g_14_136 (.ZN (n_14_136), .A (n_10_138), .B (n_7_138), .C1 (n_11_136), .C2 (n_17_133) );
AOI211_X1 g_16_135 (.ZN (n_16_135), .A (n_12_137), .B (n_6_140), .C1 (n_9_137), .C2 (n_15_134) );
AOI211_X1 g_18_134 (.ZN (n_18_134), .A (n_14_136), .B (n_8_139), .C1 (n_7_138), .C2 (n_13_135) );
AOI211_X1 g_20_133 (.ZN (n_20_133), .A (n_16_135), .B (n_10_138), .C1 (n_6_140), .C2 (n_11_136) );
AOI211_X1 g_22_132 (.ZN (n_22_132), .A (n_18_134), .B (n_12_137), .C1 (n_8_139), .C2 (n_9_137) );
AOI211_X1 g_24_131 (.ZN (n_24_131), .A (n_20_133), .B (n_14_136), .C1 (n_10_138), .C2 (n_7_138) );
AOI211_X1 g_26_130 (.ZN (n_26_130), .A (n_22_132), .B (n_16_135), .C1 (n_12_137), .C2 (n_6_140) );
AOI211_X1 g_28_129 (.ZN (n_28_129), .A (n_24_131), .B (n_18_134), .C1 (n_14_136), .C2 (n_8_139) );
AOI211_X1 g_30_128 (.ZN (n_30_128), .A (n_26_130), .B (n_20_133), .C1 (n_16_135), .C2 (n_10_138) );
AOI211_X1 g_29_130 (.ZN (n_29_130), .A (n_28_129), .B (n_22_132), .C1 (n_18_134), .C2 (n_12_137) );
AOI211_X1 g_28_128 (.ZN (n_28_128), .A (n_30_128), .B (n_24_131), .C1 (n_20_133), .C2 (n_14_136) );
AOI211_X1 g_30_127 (.ZN (n_30_127), .A (n_29_130), .B (n_26_130), .C1 (n_22_132), .C2 (n_16_135) );
AOI211_X1 g_32_126 (.ZN (n_32_126), .A (n_28_128), .B (n_28_129), .C1 (n_24_131), .C2 (n_18_134) );
AOI211_X1 g_34_125 (.ZN (n_34_125), .A (n_30_127), .B (n_30_128), .C1 (n_26_130), .C2 (n_20_133) );
AOI211_X1 g_36_124 (.ZN (n_36_124), .A (n_32_126), .B (n_29_130), .C1 (n_28_129), .C2 (n_22_132) );
AOI211_X1 g_38_123 (.ZN (n_38_123), .A (n_34_125), .B (n_28_128), .C1 (n_30_128), .C2 (n_24_131) );
AOI211_X1 g_40_122 (.ZN (n_40_122), .A (n_36_124), .B (n_30_127), .C1 (n_29_130), .C2 (n_26_130) );
AOI211_X1 g_42_121 (.ZN (n_42_121), .A (n_38_123), .B (n_32_126), .C1 (n_28_128), .C2 (n_28_129) );
AOI211_X1 g_44_120 (.ZN (n_44_120), .A (n_40_122), .B (n_34_125), .C1 (n_30_127), .C2 (n_30_128) );
AOI211_X1 g_46_119 (.ZN (n_46_119), .A (n_42_121), .B (n_36_124), .C1 (n_32_126), .C2 (n_29_130) );
AOI211_X1 g_48_118 (.ZN (n_48_118), .A (n_44_120), .B (n_38_123), .C1 (n_34_125), .C2 (n_28_128) );
AOI211_X1 g_50_117 (.ZN (n_50_117), .A (n_46_119), .B (n_40_122), .C1 (n_36_124), .C2 (n_30_127) );
AOI211_X1 g_52_116 (.ZN (n_52_116), .A (n_48_118), .B (n_42_121), .C1 (n_38_123), .C2 (n_32_126) );
AOI211_X1 g_54_115 (.ZN (n_54_115), .A (n_50_117), .B (n_44_120), .C1 (n_40_122), .C2 (n_34_125) );
AOI211_X1 g_56_114 (.ZN (n_56_114), .A (n_52_116), .B (n_46_119), .C1 (n_42_121), .C2 (n_36_124) );
AOI211_X1 g_58_113 (.ZN (n_58_113), .A (n_54_115), .B (n_48_118), .C1 (n_44_120), .C2 (n_38_123) );
AOI211_X1 g_60_112 (.ZN (n_60_112), .A (n_56_114), .B (n_50_117), .C1 (n_46_119), .C2 (n_40_122) );
AOI211_X1 g_62_113 (.ZN (n_62_113), .A (n_58_113), .B (n_52_116), .C1 (n_48_118), .C2 (n_42_121) );
AOI211_X1 g_60_114 (.ZN (n_60_114), .A (n_60_112), .B (n_54_115), .C1 (n_50_117), .C2 (n_44_120) );
AOI211_X1 g_58_115 (.ZN (n_58_115), .A (n_62_113), .B (n_56_114), .C1 (n_52_116), .C2 (n_46_119) );
AOI211_X1 g_56_116 (.ZN (n_56_116), .A (n_60_114), .B (n_58_113), .C1 (n_54_115), .C2 (n_48_118) );
AOI211_X1 g_54_117 (.ZN (n_54_117), .A (n_58_115), .B (n_60_112), .C1 (n_56_114), .C2 (n_50_117) );
AOI211_X1 g_52_118 (.ZN (n_52_118), .A (n_56_116), .B (n_62_113), .C1 (n_58_113), .C2 (n_52_116) );
AOI211_X1 g_50_119 (.ZN (n_50_119), .A (n_54_117), .B (n_60_114), .C1 (n_60_112), .C2 (n_54_115) );
AOI211_X1 g_48_120 (.ZN (n_48_120), .A (n_52_118), .B (n_58_115), .C1 (n_62_113), .C2 (n_56_114) );
AOI211_X1 g_46_121 (.ZN (n_46_121), .A (n_50_119), .B (n_56_116), .C1 (n_60_114), .C2 (n_58_113) );
AOI211_X1 g_44_122 (.ZN (n_44_122), .A (n_48_120), .B (n_54_117), .C1 (n_58_115), .C2 (n_60_112) );
AOI211_X1 g_42_123 (.ZN (n_42_123), .A (n_46_121), .B (n_52_118), .C1 (n_56_116), .C2 (n_62_113) );
AOI211_X1 g_40_124 (.ZN (n_40_124), .A (n_44_122), .B (n_50_119), .C1 (n_54_117), .C2 (n_60_114) );
AOI211_X1 g_38_125 (.ZN (n_38_125), .A (n_42_123), .B (n_48_120), .C1 (n_52_118), .C2 (n_58_115) );
AOI211_X1 g_36_126 (.ZN (n_36_126), .A (n_40_124), .B (n_46_121), .C1 (n_50_119), .C2 (n_56_116) );
AOI211_X1 g_34_127 (.ZN (n_34_127), .A (n_38_125), .B (n_44_122), .C1 (n_48_120), .C2 (n_54_117) );
AOI211_X1 g_32_128 (.ZN (n_32_128), .A (n_36_126), .B (n_42_123), .C1 (n_46_121), .C2 (n_52_118) );
AOI211_X1 g_30_129 (.ZN (n_30_129), .A (n_34_127), .B (n_40_124), .C1 (n_44_122), .C2 (n_50_119) );
AOI211_X1 g_28_130 (.ZN (n_28_130), .A (n_32_128), .B (n_38_125), .C1 (n_42_123), .C2 (n_48_120) );
AOI211_X1 g_26_129 (.ZN (n_26_129), .A (n_30_129), .B (n_36_126), .C1 (n_40_124), .C2 (n_46_121) );
AOI211_X1 g_24_130 (.ZN (n_24_130), .A (n_28_130), .B (n_34_127), .C1 (n_38_125), .C2 (n_44_122) );
AOI211_X1 g_22_131 (.ZN (n_22_131), .A (n_26_129), .B (n_32_128), .C1 (n_36_126), .C2 (n_42_123) );
AOI211_X1 g_20_132 (.ZN (n_20_132), .A (n_24_130), .B (n_30_129), .C1 (n_34_127), .C2 (n_40_124) );
AOI211_X1 g_18_133 (.ZN (n_18_133), .A (n_22_131), .B (n_28_130), .C1 (n_32_128), .C2 (n_38_125) );
AOI211_X1 g_16_134 (.ZN (n_16_134), .A (n_20_132), .B (n_26_129), .C1 (n_30_129), .C2 (n_36_126) );
AOI211_X1 g_14_135 (.ZN (n_14_135), .A (n_18_133), .B (n_24_130), .C1 (n_28_130), .C2 (n_34_127) );
AOI211_X1 g_13_137 (.ZN (n_13_137), .A (n_16_134), .B (n_22_131), .C1 (n_26_129), .C2 (n_32_128) );
AOI211_X1 g_15_136 (.ZN (n_15_136), .A (n_14_135), .B (n_20_132), .C1 (n_24_130), .C2 (n_30_129) );
AOI211_X1 g_17_135 (.ZN (n_17_135), .A (n_13_137), .B (n_18_133), .C1 (n_22_131), .C2 (n_28_130) );
AOI211_X1 g_19_134 (.ZN (n_19_134), .A (n_15_136), .B (n_16_134), .C1 (n_20_132), .C2 (n_26_129) );
AOI211_X1 g_21_133 (.ZN (n_21_133), .A (n_17_135), .B (n_14_135), .C1 (n_18_133), .C2 (n_24_130) );
AOI211_X1 g_23_132 (.ZN (n_23_132), .A (n_19_134), .B (n_13_137), .C1 (n_16_134), .C2 (n_22_131) );
AOI211_X1 g_25_131 (.ZN (n_25_131), .A (n_21_133), .B (n_15_136), .C1 (n_14_135), .C2 (n_20_132) );
AOI211_X1 g_27_130 (.ZN (n_27_130), .A (n_23_132), .B (n_17_135), .C1 (n_13_137), .C2 (n_18_133) );
AOI211_X1 g_29_129 (.ZN (n_29_129), .A (n_25_131), .B (n_19_134), .C1 (n_15_136), .C2 (n_16_134) );
AOI211_X1 g_31_128 (.ZN (n_31_128), .A (n_27_130), .B (n_21_133), .C1 (n_17_135), .C2 (n_14_135) );
AOI211_X1 g_33_127 (.ZN (n_33_127), .A (n_29_129), .B (n_23_132), .C1 (n_19_134), .C2 (n_13_137) );
AOI211_X1 g_35_126 (.ZN (n_35_126), .A (n_31_128), .B (n_25_131), .C1 (n_21_133), .C2 (n_15_136) );
AOI211_X1 g_37_125 (.ZN (n_37_125), .A (n_33_127), .B (n_27_130), .C1 (n_23_132), .C2 (n_17_135) );
AOI211_X1 g_39_124 (.ZN (n_39_124), .A (n_35_126), .B (n_29_129), .C1 (n_25_131), .C2 (n_19_134) );
AOI211_X1 g_41_123 (.ZN (n_41_123), .A (n_37_125), .B (n_31_128), .C1 (n_27_130), .C2 (n_21_133) );
AOI211_X1 g_43_122 (.ZN (n_43_122), .A (n_39_124), .B (n_33_127), .C1 (n_29_129), .C2 (n_23_132) );
AOI211_X1 g_45_121 (.ZN (n_45_121), .A (n_41_123), .B (n_35_126), .C1 (n_31_128), .C2 (n_25_131) );
AOI211_X1 g_47_120 (.ZN (n_47_120), .A (n_43_122), .B (n_37_125), .C1 (n_33_127), .C2 (n_27_130) );
AOI211_X1 g_49_119 (.ZN (n_49_119), .A (n_45_121), .B (n_39_124), .C1 (n_35_126), .C2 (n_29_129) );
AOI211_X1 g_51_118 (.ZN (n_51_118), .A (n_47_120), .B (n_41_123), .C1 (n_37_125), .C2 (n_31_128) );
AOI211_X1 g_53_117 (.ZN (n_53_117), .A (n_49_119), .B (n_43_122), .C1 (n_39_124), .C2 (n_33_127) );
AOI211_X1 g_55_116 (.ZN (n_55_116), .A (n_51_118), .B (n_45_121), .C1 (n_41_123), .C2 (n_35_126) );
AOI211_X1 g_57_115 (.ZN (n_57_115), .A (n_53_117), .B (n_47_120), .C1 (n_43_122), .C2 (n_37_125) );
AOI211_X1 g_59_114 (.ZN (n_59_114), .A (n_55_116), .B (n_49_119), .C1 (n_45_121), .C2 (n_39_124) );
AOI211_X1 g_61_113 (.ZN (n_61_113), .A (n_57_115), .B (n_51_118), .C1 (n_47_120), .C2 (n_41_123) );
AOI211_X1 g_63_114 (.ZN (n_63_114), .A (n_59_114), .B (n_53_117), .C1 (n_49_119), .C2 (n_43_122) );
AOI211_X1 g_61_115 (.ZN (n_61_115), .A (n_61_113), .B (n_55_116), .C1 (n_51_118), .C2 (n_45_121) );
AOI211_X1 g_59_116 (.ZN (n_59_116), .A (n_63_114), .B (n_57_115), .C1 (n_53_117), .C2 (n_47_120) );
AOI211_X1 g_57_117 (.ZN (n_57_117), .A (n_61_115), .B (n_59_114), .C1 (n_55_116), .C2 (n_49_119) );
AOI211_X1 g_55_118 (.ZN (n_55_118), .A (n_59_116), .B (n_61_113), .C1 (n_57_115), .C2 (n_51_118) );
AOI211_X1 g_53_119 (.ZN (n_53_119), .A (n_57_117), .B (n_63_114), .C1 (n_59_114), .C2 (n_53_117) );
AOI211_X1 g_51_120 (.ZN (n_51_120), .A (n_55_118), .B (n_61_115), .C1 (n_61_113), .C2 (n_55_116) );
AOI211_X1 g_49_121 (.ZN (n_49_121), .A (n_53_119), .B (n_59_116), .C1 (n_63_114), .C2 (n_57_115) );
AOI211_X1 g_47_122 (.ZN (n_47_122), .A (n_51_120), .B (n_57_117), .C1 (n_61_115), .C2 (n_59_114) );
AOI211_X1 g_45_123 (.ZN (n_45_123), .A (n_49_121), .B (n_55_118), .C1 (n_59_116), .C2 (n_61_113) );
AOI211_X1 g_43_124 (.ZN (n_43_124), .A (n_47_122), .B (n_53_119), .C1 (n_57_117), .C2 (n_63_114) );
AOI211_X1 g_41_125 (.ZN (n_41_125), .A (n_45_123), .B (n_51_120), .C1 (n_55_118), .C2 (n_61_115) );
AOI211_X1 g_39_126 (.ZN (n_39_126), .A (n_43_124), .B (n_49_121), .C1 (n_53_119), .C2 (n_59_116) );
AOI211_X1 g_37_127 (.ZN (n_37_127), .A (n_41_125), .B (n_47_122), .C1 (n_51_120), .C2 (n_57_117) );
AOI211_X1 g_35_128 (.ZN (n_35_128), .A (n_39_126), .B (n_45_123), .C1 (n_49_121), .C2 (n_55_118) );
AOI211_X1 g_33_129 (.ZN (n_33_129), .A (n_37_127), .B (n_43_124), .C1 (n_47_122), .C2 (n_53_119) );
AOI211_X1 g_31_130 (.ZN (n_31_130), .A (n_35_128), .B (n_41_125), .C1 (n_45_123), .C2 (n_51_120) );
AOI211_X1 g_29_131 (.ZN (n_29_131), .A (n_33_129), .B (n_39_126), .C1 (n_43_124), .C2 (n_49_121) );
AOI211_X1 g_27_132 (.ZN (n_27_132), .A (n_31_130), .B (n_37_127), .C1 (n_41_125), .C2 (n_47_122) );
AOI211_X1 g_25_133 (.ZN (n_25_133), .A (n_29_131), .B (n_35_128), .C1 (n_39_126), .C2 (n_45_123) );
AOI211_X1 g_26_131 (.ZN (n_26_131), .A (n_27_132), .B (n_33_129), .C1 (n_37_127), .C2 (n_43_124) );
AOI211_X1 g_24_132 (.ZN (n_24_132), .A (n_25_133), .B (n_31_130), .C1 (n_35_128), .C2 (n_41_125) );
AOI211_X1 g_22_133 (.ZN (n_22_133), .A (n_26_131), .B (n_29_131), .C1 (n_33_129), .C2 (n_39_126) );
AOI211_X1 g_20_134 (.ZN (n_20_134), .A (n_24_132), .B (n_27_132), .C1 (n_31_130), .C2 (n_37_127) );
AOI211_X1 g_18_135 (.ZN (n_18_135), .A (n_22_133), .B (n_25_133), .C1 (n_29_131), .C2 (n_35_128) );
AOI211_X1 g_16_136 (.ZN (n_16_136), .A (n_20_134), .B (n_26_131), .C1 (n_27_132), .C2 (n_33_129) );
AOI211_X1 g_14_137 (.ZN (n_14_137), .A (n_18_135), .B (n_24_132), .C1 (n_25_133), .C2 (n_31_130) );
AOI211_X1 g_12_138 (.ZN (n_12_138), .A (n_16_136), .B (n_22_133), .C1 (n_26_131), .C2 (n_29_131) );
AOI211_X1 g_10_139 (.ZN (n_10_139), .A (n_14_137), .B (n_20_134), .C1 (n_24_132), .C2 (n_27_132) );
AOI211_X1 g_8_140 (.ZN (n_8_140), .A (n_12_138), .B (n_18_135), .C1 (n_22_133), .C2 (n_25_133) );
AOI211_X1 g_6_139 (.ZN (n_6_139), .A (n_10_139), .B (n_16_136), .C1 (n_20_134), .C2 (n_26_131) );
AOI211_X1 g_5_141 (.ZN (n_5_141), .A (n_8_140), .B (n_14_137), .C1 (n_18_135), .C2 (n_24_132) );
AOI211_X1 g_4_143 (.ZN (n_4_143), .A (n_6_139), .B (n_12_138), .C1 (n_16_136), .C2 (n_22_133) );
AOI211_X1 g_5_145 (.ZN (n_5_145), .A (n_5_141), .B (n_10_139), .C1 (n_14_137), .C2 (n_20_134) );
AOI211_X1 g_7_144 (.ZN (n_7_144), .A (n_4_143), .B (n_8_140), .C1 (n_12_138), .C2 (n_18_135) );
AOI211_X1 g_6_142 (.ZN (n_6_142), .A (n_5_145), .B (n_6_139), .C1 (n_10_139), .C2 (n_16_136) );
AOI211_X1 g_7_140 (.ZN (n_7_140), .A (n_7_144), .B (n_5_141), .C1 (n_8_140), .C2 (n_14_137) );
AOI211_X1 g_9_139 (.ZN (n_9_139), .A (n_6_142), .B (n_4_143), .C1 (n_6_139), .C2 (n_12_138) );
AOI211_X1 g_11_138 (.ZN (n_11_138), .A (n_7_140), .B (n_5_145), .C1 (n_5_141), .C2 (n_10_139) );
AOI211_X1 g_10_140 (.ZN (n_10_140), .A (n_9_139), .B (n_7_144), .C1 (n_4_143), .C2 (n_8_140) );
AOI211_X1 g_8_141 (.ZN (n_8_141), .A (n_11_138), .B (n_6_142), .C1 (n_5_145), .C2 (n_6_139) );
AOI211_X1 g_9_143 (.ZN (n_9_143), .A (n_10_140), .B (n_7_140), .C1 (n_7_144), .C2 (n_5_141) );
AOI211_X1 g_7_142 (.ZN (n_7_142), .A (n_8_141), .B (n_9_139), .C1 (n_6_142), .C2 (n_4_143) );
AOI211_X1 g_6_144 (.ZN (n_6_144), .A (n_9_143), .B (n_11_138), .C1 (n_7_140), .C2 (n_5_145) );
AOI211_X1 g_7_146 (.ZN (n_7_146), .A (n_7_142), .B (n_10_140), .C1 (n_9_139), .C2 (n_7_144) );
AOI211_X1 g_9_147 (.ZN (n_9_147), .A (n_6_144), .B (n_8_141), .C1 (n_11_138), .C2 (n_6_142) );
AOI211_X1 g_8_145 (.ZN (n_8_145), .A (n_7_146), .B (n_9_143), .C1 (n_10_140), .C2 (n_7_140) );
AOI211_X1 g_10_146 (.ZN (n_10_146), .A (n_9_147), .B (n_7_142), .C1 (n_8_141), .C2 (n_9_139) );
AOI211_X1 g_11_148 (.ZN (n_11_148), .A (n_8_145), .B (n_6_144), .C1 (n_9_143), .C2 (n_11_138) );
AOI211_X1 g_12_146 (.ZN (n_12_146), .A (n_10_146), .B (n_7_146), .C1 (n_7_142), .C2 (n_10_140) );
AOI211_X1 g_10_145 (.ZN (n_10_145), .A (n_11_148), .B (n_9_147), .C1 (n_6_144), .C2 (n_8_141) );
AOI211_X1 g_8_144 (.ZN (n_8_144), .A (n_12_146), .B (n_8_145), .C1 (n_7_146), .C2 (n_9_143) );
AOI211_X1 g_6_143 (.ZN (n_6_143), .A (n_10_145), .B (n_10_146), .C1 (n_9_147), .C2 (n_7_142) );
AOI211_X1 g_7_141 (.ZN (n_7_141), .A (n_8_144), .B (n_11_148), .C1 (n_8_145), .C2 (n_6_144) );
AOI211_X1 g_9_142 (.ZN (n_9_142), .A (n_6_143), .B (n_12_146), .C1 (n_10_146), .C2 (n_7_146) );
AOI211_X1 g_11_141 (.ZN (n_11_141), .A (n_7_141), .B (n_10_145), .C1 (n_11_148), .C2 (n_9_147) );
AOI211_X1 g_12_139 (.ZN (n_12_139), .A (n_9_142), .B (n_8_144), .C1 (n_12_146), .C2 (n_8_145) );
AOI211_X1 g_14_138 (.ZN (n_14_138), .A (n_11_141), .B (n_6_143), .C1 (n_10_145), .C2 (n_10_146) );
AOI211_X1 g_16_137 (.ZN (n_16_137), .A (n_12_139), .B (n_7_141), .C1 (n_8_144), .C2 (n_11_148) );
AOI211_X1 g_18_136 (.ZN (n_18_136), .A (n_14_138), .B (n_9_142), .C1 (n_6_143), .C2 (n_12_146) );
AOI211_X1 g_20_135 (.ZN (n_20_135), .A (n_16_137), .B (n_11_141), .C1 (n_7_141), .C2 (n_10_145) );
AOI211_X1 g_22_134 (.ZN (n_22_134), .A (n_18_136), .B (n_12_139), .C1 (n_9_142), .C2 (n_8_144) );
AOI211_X1 g_24_133 (.ZN (n_24_133), .A (n_20_135), .B (n_14_138), .C1 (n_11_141), .C2 (n_6_143) );
AOI211_X1 g_26_132 (.ZN (n_26_132), .A (n_22_134), .B (n_16_137), .C1 (n_12_139), .C2 (n_7_141) );
AOI211_X1 g_28_131 (.ZN (n_28_131), .A (n_24_133), .B (n_18_136), .C1 (n_14_138), .C2 (n_9_142) );
AOI211_X1 g_30_130 (.ZN (n_30_130), .A (n_26_132), .B (n_20_135), .C1 (n_16_137), .C2 (n_11_141) );
AOI211_X1 g_32_129 (.ZN (n_32_129), .A (n_28_131), .B (n_22_134), .C1 (n_18_136), .C2 (n_12_139) );
AOI211_X1 g_34_128 (.ZN (n_34_128), .A (n_30_130), .B (n_24_133), .C1 (n_20_135), .C2 (n_14_138) );
AOI211_X1 g_36_127 (.ZN (n_36_127), .A (n_32_129), .B (n_26_132), .C1 (n_22_134), .C2 (n_16_137) );
AOI211_X1 g_38_126 (.ZN (n_38_126), .A (n_34_128), .B (n_28_131), .C1 (n_24_133), .C2 (n_18_136) );
AOI211_X1 g_40_125 (.ZN (n_40_125), .A (n_36_127), .B (n_30_130), .C1 (n_26_132), .C2 (n_20_135) );
AOI211_X1 g_42_124 (.ZN (n_42_124), .A (n_38_126), .B (n_32_129), .C1 (n_28_131), .C2 (n_22_134) );
AOI211_X1 g_44_123 (.ZN (n_44_123), .A (n_40_125), .B (n_34_128), .C1 (n_30_130), .C2 (n_24_133) );
AOI211_X1 g_46_122 (.ZN (n_46_122), .A (n_42_124), .B (n_36_127), .C1 (n_32_129), .C2 (n_26_132) );
AOI211_X1 g_48_121 (.ZN (n_48_121), .A (n_44_123), .B (n_38_126), .C1 (n_34_128), .C2 (n_28_131) );
AOI211_X1 g_50_120 (.ZN (n_50_120), .A (n_46_122), .B (n_40_125), .C1 (n_36_127), .C2 (n_30_130) );
AOI211_X1 g_52_119 (.ZN (n_52_119), .A (n_48_121), .B (n_42_124), .C1 (n_38_126), .C2 (n_32_129) );
AOI211_X1 g_54_118 (.ZN (n_54_118), .A (n_50_120), .B (n_44_123), .C1 (n_40_125), .C2 (n_34_128) );
AOI211_X1 g_56_117 (.ZN (n_56_117), .A (n_52_119), .B (n_46_122), .C1 (n_42_124), .C2 (n_36_127) );
AOI211_X1 g_58_116 (.ZN (n_58_116), .A (n_54_118), .B (n_48_121), .C1 (n_44_123), .C2 (n_38_126) );
AOI211_X1 g_60_115 (.ZN (n_60_115), .A (n_56_117), .B (n_50_120), .C1 (n_46_122), .C2 (n_40_125) );
AOI211_X1 g_62_114 (.ZN (n_62_114), .A (n_58_116), .B (n_52_119), .C1 (n_48_121), .C2 (n_42_124) );
AOI211_X1 g_61_116 (.ZN (n_61_116), .A (n_60_115), .B (n_54_118), .C1 (n_50_120), .C2 (n_44_123) );
AOI211_X1 g_59_115 (.ZN (n_59_115), .A (n_62_114), .B (n_56_117), .C1 (n_52_119), .C2 (n_46_122) );
AOI211_X1 g_61_114 (.ZN (n_61_114), .A (n_61_116), .B (n_58_116), .C1 (n_54_118), .C2 (n_48_121) );
AOI211_X1 g_63_113 (.ZN (n_63_113), .A (n_59_115), .B (n_60_115), .C1 (n_56_117), .C2 (n_50_120) );
AOI211_X1 g_65_112 (.ZN (n_65_112), .A (n_61_114), .B (n_62_114), .C1 (n_58_116), .C2 (n_52_119) );
AOI211_X1 g_67_111 (.ZN (n_67_111), .A (n_63_113), .B (n_61_116), .C1 (n_60_115), .C2 (n_54_118) );
AOI211_X1 g_69_110 (.ZN (n_69_110), .A (n_65_112), .B (n_59_115), .C1 (n_62_114), .C2 (n_56_117) );
AOI211_X1 g_71_109 (.ZN (n_71_109), .A (n_67_111), .B (n_61_114), .C1 (n_61_116), .C2 (n_58_116) );
AOI211_X1 g_73_108 (.ZN (n_73_108), .A (n_69_110), .B (n_63_113), .C1 (n_59_115), .C2 (n_60_115) );
AOI211_X1 g_75_107 (.ZN (n_75_107), .A (n_71_109), .B (n_65_112), .C1 (n_61_114), .C2 (n_62_114) );
AOI211_X1 g_76_105 (.ZN (n_76_105), .A (n_73_108), .B (n_67_111), .C1 (n_63_113), .C2 (n_61_116) );
AOI211_X1 g_78_104 (.ZN (n_78_104), .A (n_75_107), .B (n_69_110), .C1 (n_65_112), .C2 (n_59_115) );
AOI211_X1 g_77_106 (.ZN (n_77_106), .A (n_76_105), .B (n_71_109), .C1 (n_67_111), .C2 (n_61_114) );
AOI211_X1 g_79_105 (.ZN (n_79_105), .A (n_78_104), .B (n_73_108), .C1 (n_69_110), .C2 (n_63_113) );
AOI211_X1 g_78_107 (.ZN (n_78_107), .A (n_77_106), .B (n_75_107), .C1 (n_71_109), .C2 (n_65_112) );
AOI211_X1 g_76_106 (.ZN (n_76_106), .A (n_79_105), .B (n_76_105), .C1 (n_73_108), .C2 (n_67_111) );
AOI211_X1 g_78_105 (.ZN (n_78_105), .A (n_78_107), .B (n_78_104), .C1 (n_75_107), .C2 (n_69_110) );
AOI211_X1 g_80_104 (.ZN (n_80_104), .A (n_76_106), .B (n_77_106), .C1 (n_76_105), .C2 (n_71_109) );
AOI211_X1 g_79_106 (.ZN (n_79_106), .A (n_78_105), .B (n_79_105), .C1 (n_78_104), .C2 (n_73_108) );
AOI211_X1 g_81_105 (.ZN (n_81_105), .A (n_80_104), .B (n_78_107), .C1 (n_77_106), .C2 (n_75_107) );
AOI211_X1 g_83_104 (.ZN (n_83_104), .A (n_79_106), .B (n_76_106), .C1 (n_79_105), .C2 (n_76_105) );
AOI211_X1 g_85_103 (.ZN (n_85_103), .A (n_81_105), .B (n_78_105), .C1 (n_78_107), .C2 (n_78_104) );
AOI211_X1 g_87_102 (.ZN (n_87_102), .A (n_83_104), .B (n_80_104), .C1 (n_76_106), .C2 (n_77_106) );
AOI211_X1 g_89_101 (.ZN (n_89_101), .A (n_85_103), .B (n_79_106), .C1 (n_78_105), .C2 (n_79_105) );
AOI211_X1 g_91_100 (.ZN (n_91_100), .A (n_87_102), .B (n_81_105), .C1 (n_80_104), .C2 (n_78_107) );
AOI211_X1 g_93_99 (.ZN (n_93_99), .A (n_89_101), .B (n_83_104), .C1 (n_79_106), .C2 (n_76_106) );
AOI211_X1 g_95_98 (.ZN (n_95_98), .A (n_91_100), .B (n_85_103), .C1 (n_81_105), .C2 (n_78_105) );
AOI211_X1 g_97_97 (.ZN (n_97_97), .A (n_93_99), .B (n_87_102), .C1 (n_83_104), .C2 (n_80_104) );
AOI211_X1 g_99_96 (.ZN (n_99_96), .A (n_95_98), .B (n_89_101), .C1 (n_85_103), .C2 (n_79_106) );
AOI211_X1 g_101_95 (.ZN (n_101_95), .A (n_97_97), .B (n_91_100), .C1 (n_87_102), .C2 (n_81_105) );
AOI211_X1 g_100_97 (.ZN (n_100_97), .A (n_99_96), .B (n_93_99), .C1 (n_89_101), .C2 (n_83_104) );
AOI211_X1 g_98_96 (.ZN (n_98_96), .A (n_101_95), .B (n_95_98), .C1 (n_91_100), .C2 (n_85_103) );
AOI211_X1 g_100_95 (.ZN (n_100_95), .A (n_100_97), .B (n_97_97), .C1 (n_93_99), .C2 (n_87_102) );
AOI211_X1 g_102_94 (.ZN (n_102_94), .A (n_98_96), .B (n_99_96), .C1 (n_95_98), .C2 (n_89_101) );
AOI211_X1 g_104_93 (.ZN (n_104_93), .A (n_100_95), .B (n_101_95), .C1 (n_97_97), .C2 (n_91_100) );
AOI211_X1 g_106_92 (.ZN (n_106_92), .A (n_102_94), .B (n_100_97), .C1 (n_99_96), .C2 (n_93_99) );
AOI211_X1 g_105_94 (.ZN (n_105_94), .A (n_104_93), .B (n_98_96), .C1 (n_101_95), .C2 (n_95_98) );
AOI211_X1 g_107_93 (.ZN (n_107_93), .A (n_106_92), .B (n_100_95), .C1 (n_100_97), .C2 (n_97_97) );
AOI211_X1 g_106_95 (.ZN (n_106_95), .A (n_105_94), .B (n_102_94), .C1 (n_98_96), .C2 (n_99_96) );
AOI211_X1 g_104_94 (.ZN (n_104_94), .A (n_107_93), .B (n_104_93), .C1 (n_100_95), .C2 (n_101_95) );
AOI211_X1 g_106_93 (.ZN (n_106_93), .A (n_106_95), .B (n_106_92), .C1 (n_102_94), .C2 (n_100_97) );
AOI211_X1 g_108_92 (.ZN (n_108_92), .A (n_104_94), .B (n_105_94), .C1 (n_104_93), .C2 (n_98_96) );
AOI211_X1 g_110_91 (.ZN (n_110_91), .A (n_106_93), .B (n_107_93), .C1 (n_106_92), .C2 (n_100_95) );
AOI211_X1 g_112_90 (.ZN (n_112_90), .A (n_108_92), .B (n_106_95), .C1 (n_105_94), .C2 (n_102_94) );
AOI211_X1 g_114_89 (.ZN (n_114_89), .A (n_110_91), .B (n_104_94), .C1 (n_107_93), .C2 (n_104_93) );
AOI211_X1 g_116_88 (.ZN (n_116_88), .A (n_112_90), .B (n_106_93), .C1 (n_106_95), .C2 (n_106_92) );
AOI211_X1 g_118_89 (.ZN (n_118_89), .A (n_114_89), .B (n_108_92), .C1 (n_104_94), .C2 (n_105_94) );
AOI211_X1 g_116_90 (.ZN (n_116_90), .A (n_116_88), .B (n_110_91), .C1 (n_106_93), .C2 (n_107_93) );
AOI211_X1 g_114_91 (.ZN (n_114_91), .A (n_118_89), .B (n_112_90), .C1 (n_108_92), .C2 (n_106_95) );
AOI211_X1 g_112_92 (.ZN (n_112_92), .A (n_116_90), .B (n_114_89), .C1 (n_110_91), .C2 (n_104_94) );
AOI211_X1 g_110_93 (.ZN (n_110_93), .A (n_114_91), .B (n_116_88), .C1 (n_112_90), .C2 (n_106_93) );
AOI211_X1 g_108_94 (.ZN (n_108_94), .A (n_112_92), .B (n_118_89), .C1 (n_114_89), .C2 (n_108_92) );
AOI211_X1 g_107_96 (.ZN (n_107_96), .A (n_110_93), .B (n_116_90), .C1 (n_116_88), .C2 (n_110_91) );
AOI211_X1 g_106_94 (.ZN (n_106_94), .A (n_108_94), .B (n_114_91), .C1 (n_118_89), .C2 (n_112_90) );
AOI211_X1 g_108_93 (.ZN (n_108_93), .A (n_107_96), .B (n_112_92), .C1 (n_116_90), .C2 (n_114_89) );
AOI211_X1 g_110_92 (.ZN (n_110_92), .A (n_106_94), .B (n_110_93), .C1 (n_114_91), .C2 (n_116_88) );
AOI211_X1 g_112_91 (.ZN (n_112_91), .A (n_108_93), .B (n_108_94), .C1 (n_112_92), .C2 (n_118_89) );
AOI211_X1 g_111_93 (.ZN (n_111_93), .A (n_110_92), .B (n_107_96), .C1 (n_110_93), .C2 (n_116_90) );
AOI211_X1 g_113_92 (.ZN (n_113_92), .A (n_112_91), .B (n_106_94), .C1 (n_108_94), .C2 (n_114_91) );
AOI211_X1 g_115_91 (.ZN (n_115_91), .A (n_111_93), .B (n_108_93), .C1 (n_107_96), .C2 (n_112_92) );
AOI211_X1 g_117_90 (.ZN (n_117_90), .A (n_113_92), .B (n_110_92), .C1 (n_106_94), .C2 (n_110_93) );
AOI211_X1 g_119_89 (.ZN (n_119_89), .A (n_115_91), .B (n_112_91), .C1 (n_108_93), .C2 (n_108_94) );
AOI211_X1 g_121_88 (.ZN (n_121_88), .A (n_117_90), .B (n_111_93), .C1 (n_110_92), .C2 (n_107_96) );
AOI211_X1 g_123_87 (.ZN (n_123_87), .A (n_119_89), .B (n_113_92), .C1 (n_112_91), .C2 (n_106_94) );
AOI211_X1 g_122_89 (.ZN (n_122_89), .A (n_121_88), .B (n_115_91), .C1 (n_111_93), .C2 (n_108_93) );
AOI211_X1 g_121_87 (.ZN (n_121_87), .A (n_123_87), .B (n_117_90), .C1 (n_113_92), .C2 (n_110_92) );
AOI211_X1 g_119_88 (.ZN (n_119_88), .A (n_122_89), .B (n_119_89), .C1 (n_115_91), .C2 (n_112_91) );
AOI211_X1 g_117_89 (.ZN (n_117_89), .A (n_121_87), .B (n_121_88), .C1 (n_117_90), .C2 (n_111_93) );
AOI211_X1 g_115_90 (.ZN (n_115_90), .A (n_119_88), .B (n_123_87), .C1 (n_119_89), .C2 (n_113_92) );
AOI211_X1 g_113_91 (.ZN (n_113_91), .A (n_117_89), .B (n_122_89), .C1 (n_121_88), .C2 (n_115_91) );
AOI211_X1 g_111_92 (.ZN (n_111_92), .A (n_115_90), .B (n_121_87), .C1 (n_123_87), .C2 (n_117_90) );
AOI211_X1 g_109_93 (.ZN (n_109_93), .A (n_113_91), .B (n_119_88), .C1 (n_122_89), .C2 (n_119_89) );
AOI211_X1 g_107_94 (.ZN (n_107_94), .A (n_111_92), .B (n_117_89), .C1 (n_121_87), .C2 (n_121_88) );
AOI211_X1 g_105_95 (.ZN (n_105_95), .A (n_109_93), .B (n_115_90), .C1 (n_119_88), .C2 (n_123_87) );
AOI211_X1 g_103_96 (.ZN (n_103_96), .A (n_107_94), .B (n_113_91), .C1 (n_117_89), .C2 (n_122_89) );
AOI211_X1 g_101_97 (.ZN (n_101_97), .A (n_105_95), .B (n_111_92), .C1 (n_115_90), .C2 (n_121_87) );
AOI211_X1 g_102_95 (.ZN (n_102_95), .A (n_103_96), .B (n_109_93), .C1 (n_113_91), .C2 (n_119_88) );
AOI211_X1 g_100_96 (.ZN (n_100_96), .A (n_101_97), .B (n_107_94), .C1 (n_111_92), .C2 (n_117_89) );
AOI211_X1 g_98_97 (.ZN (n_98_97), .A (n_102_95), .B (n_105_95), .C1 (n_109_93), .C2 (n_115_90) );
AOI211_X1 g_96_98 (.ZN (n_96_98), .A (n_100_96), .B (n_103_96), .C1 (n_107_94), .C2 (n_113_91) );
AOI211_X1 g_94_99 (.ZN (n_94_99), .A (n_98_97), .B (n_101_97), .C1 (n_105_95), .C2 (n_111_92) );
AOI211_X1 g_92_100 (.ZN (n_92_100), .A (n_96_98), .B (n_102_95), .C1 (n_103_96), .C2 (n_109_93) );
AOI211_X1 g_90_101 (.ZN (n_90_101), .A (n_94_99), .B (n_100_96), .C1 (n_101_97), .C2 (n_107_94) );
AOI211_X1 g_88_102 (.ZN (n_88_102), .A (n_92_100), .B (n_98_97), .C1 (n_102_95), .C2 (n_105_95) );
AOI211_X1 g_86_103 (.ZN (n_86_103), .A (n_90_101), .B (n_96_98), .C1 (n_100_96), .C2 (n_103_96) );
AOI211_X1 g_84_104 (.ZN (n_84_104), .A (n_88_102), .B (n_94_99), .C1 (n_98_97), .C2 (n_101_97) );
AOI211_X1 g_82_105 (.ZN (n_82_105), .A (n_86_103), .B (n_92_100), .C1 (n_96_98), .C2 (n_102_95) );
AOI211_X1 g_80_106 (.ZN (n_80_106), .A (n_84_104), .B (n_90_101), .C1 (n_94_99), .C2 (n_100_96) );
AOI211_X1 g_82_107 (.ZN (n_82_107), .A (n_82_105), .B (n_88_102), .C1 (n_92_100), .C2 (n_98_97) );
AOI211_X1 g_84_106 (.ZN (n_84_106), .A (n_80_106), .B (n_86_103), .C1 (n_90_101), .C2 (n_96_98) );
AOI211_X1 g_86_105 (.ZN (n_86_105), .A (n_82_107), .B (n_84_104), .C1 (n_88_102), .C2 (n_94_99) );
AOI211_X1 g_88_104 (.ZN (n_88_104), .A (n_84_106), .B (n_82_105), .C1 (n_86_103), .C2 (n_92_100) );
AOI211_X1 g_90_103 (.ZN (n_90_103), .A (n_86_105), .B (n_80_106), .C1 (n_84_104), .C2 (n_90_101) );
AOI211_X1 g_92_102 (.ZN (n_92_102), .A (n_88_104), .B (n_82_107), .C1 (n_82_105), .C2 (n_88_102) );
AOI211_X1 g_94_101 (.ZN (n_94_101), .A (n_90_103), .B (n_84_106), .C1 (n_80_106), .C2 (n_86_103) );
AOI211_X1 g_96_100 (.ZN (n_96_100), .A (n_92_102), .B (n_86_105), .C1 (n_82_107), .C2 (n_84_104) );
AOI211_X1 g_97_98 (.ZN (n_97_98), .A (n_94_101), .B (n_88_104), .C1 (n_84_106), .C2 (n_82_105) );
AOI211_X1 g_99_97 (.ZN (n_99_97), .A (n_96_100), .B (n_90_103), .C1 (n_86_105), .C2 (n_80_106) );
AOI211_X1 g_101_96 (.ZN (n_101_96), .A (n_97_98), .B (n_92_102), .C1 (n_88_104), .C2 (n_82_107) );
AOI211_X1 g_103_95 (.ZN (n_103_95), .A (n_99_97), .B (n_94_101), .C1 (n_90_103), .C2 (n_84_106) );
AOI211_X1 g_102_97 (.ZN (n_102_97), .A (n_101_96), .B (n_96_100), .C1 (n_92_102), .C2 (n_86_105) );
AOI211_X1 g_104_96 (.ZN (n_104_96), .A (n_103_95), .B (n_97_98), .C1 (n_94_101), .C2 (n_88_104) );
AOI211_X1 g_103_98 (.ZN (n_103_98), .A (n_102_97), .B (n_99_97), .C1 (n_96_100), .C2 (n_90_103) );
AOI211_X1 g_102_96 (.ZN (n_102_96), .A (n_104_96), .B (n_101_96), .C1 (n_97_98), .C2 (n_92_102) );
AOI211_X1 g_104_95 (.ZN (n_104_95), .A (n_103_98), .B (n_103_95), .C1 (n_99_97), .C2 (n_94_101) );
AOI211_X1 g_105_97 (.ZN (n_105_97), .A (n_102_96), .B (n_102_97), .C1 (n_101_96), .C2 (n_96_100) );
AOI211_X1 g_104_99 (.ZN (n_104_99), .A (n_104_95), .B (n_104_96), .C1 (n_103_95), .C2 (n_97_98) );
AOI211_X1 g_103_97 (.ZN (n_103_97), .A (n_105_97), .B (n_103_98), .C1 (n_102_97), .C2 (n_99_97) );
AOI211_X1 g_105_96 (.ZN (n_105_96), .A (n_104_99), .B (n_102_96), .C1 (n_104_96), .C2 (n_101_96) );
AOI211_X1 g_107_95 (.ZN (n_107_95), .A (n_103_97), .B (n_104_95), .C1 (n_103_98), .C2 (n_103_95) );
AOI211_X1 g_109_94 (.ZN (n_109_94), .A (n_105_96), .B (n_105_97), .C1 (n_102_96), .C2 (n_102_97) );
AOI211_X1 g_108_96 (.ZN (n_108_96), .A (n_107_95), .B (n_104_99), .C1 (n_104_95), .C2 (n_104_96) );
AOI211_X1 g_110_95 (.ZN (n_110_95), .A (n_109_94), .B (n_103_97), .C1 (n_105_97), .C2 (n_103_98) );
AOI211_X1 g_112_94 (.ZN (n_112_94), .A (n_108_96), .B (n_105_96), .C1 (n_104_99), .C2 (n_102_96) );
AOI211_X1 g_114_93 (.ZN (n_114_93), .A (n_110_95), .B (n_107_95), .C1 (n_103_97), .C2 (n_104_95) );
AOI211_X1 g_116_92 (.ZN (n_116_92), .A (n_112_94), .B (n_109_94), .C1 (n_105_96), .C2 (n_105_97) );
AOI211_X1 g_118_91 (.ZN (n_118_91), .A (n_114_93), .B (n_108_96), .C1 (n_107_95), .C2 (n_104_99) );
AOI211_X1 g_120_90 (.ZN (n_120_90), .A (n_116_92), .B (n_110_95), .C1 (n_109_94), .C2 (n_103_97) );
AOI211_X1 g_119_92 (.ZN (n_119_92), .A (n_118_91), .B (n_112_94), .C1 (n_108_96), .C2 (n_105_96) );
AOI211_X1 g_118_90 (.ZN (n_118_90), .A (n_120_90), .B (n_114_93), .C1 (n_110_95), .C2 (n_107_95) );
AOI211_X1 g_120_89 (.ZN (n_120_89), .A (n_119_92), .B (n_116_92), .C1 (n_112_94), .C2 (n_109_94) );
AOI211_X1 g_122_88 (.ZN (n_122_88), .A (n_118_90), .B (n_118_91), .C1 (n_114_93), .C2 (n_108_96) );
AOI211_X1 g_124_87 (.ZN (n_124_87), .A (n_120_89), .B (n_120_90), .C1 (n_116_92), .C2 (n_110_95) );
AOI211_X1 g_123_89 (.ZN (n_123_89), .A (n_122_88), .B (n_119_92), .C1 (n_118_91), .C2 (n_112_94) );
AOI211_X1 g_125_88 (.ZN (n_125_88), .A (n_124_87), .B (n_118_90), .C1 (n_120_90), .C2 (n_114_93) );
AOI211_X1 g_127_87 (.ZN (n_127_87), .A (n_123_89), .B (n_120_89), .C1 (n_119_92), .C2 (n_116_92) );
AOI211_X1 g_129_86 (.ZN (n_129_86), .A (n_125_88), .B (n_122_88), .C1 (n_118_90), .C2 (n_118_91) );
AOI211_X1 g_128_84 (.ZN (n_128_84), .A (n_127_87), .B (n_124_87), .C1 (n_120_89), .C2 (n_120_90) );
AOI211_X1 g_130_83 (.ZN (n_130_83), .A (n_129_86), .B (n_123_89), .C1 (n_122_88), .C2 (n_119_92) );
AOI211_X1 g_132_82 (.ZN (n_132_82), .A (n_128_84), .B (n_125_88), .C1 (n_124_87), .C2 (n_118_90) );
AOI211_X1 g_134_81 (.ZN (n_134_81), .A (n_130_83), .B (n_127_87), .C1 (n_123_89), .C2 (n_120_89) );
AOI211_X1 g_136_80 (.ZN (n_136_80), .A (n_132_82), .B (n_129_86), .C1 (n_125_88), .C2 (n_122_88) );
AOI211_X1 g_135_82 (.ZN (n_135_82), .A (n_134_81), .B (n_128_84), .C1 (n_127_87), .C2 (n_124_87) );
AOI211_X1 g_137_81 (.ZN (n_137_81), .A (n_136_80), .B (n_130_83), .C1 (n_129_86), .C2 (n_123_89) );
AOI211_X1 g_139_80 (.ZN (n_139_80), .A (n_135_82), .B (n_132_82), .C1 (n_128_84), .C2 (n_125_88) );
AOI211_X1 g_141_79 (.ZN (n_141_79), .A (n_137_81), .B (n_134_81), .C1 (n_130_83), .C2 (n_127_87) );
AOI211_X1 g_143_78 (.ZN (n_143_78), .A (n_139_80), .B (n_136_80), .C1 (n_132_82), .C2 (n_129_86) );
AOI211_X1 g_142_80 (.ZN (n_142_80), .A (n_141_79), .B (n_135_82), .C1 (n_134_81), .C2 (n_128_84) );
AOI211_X1 g_141_78 (.ZN (n_141_78), .A (n_143_78), .B (n_137_81), .C1 (n_136_80), .C2 (n_130_83) );
AOI211_X1 g_143_77 (.ZN (n_143_77), .A (n_142_80), .B (n_139_80), .C1 (n_135_82), .C2 (n_132_82) );
AOI211_X1 g_145_76 (.ZN (n_145_76), .A (n_141_78), .B (n_141_79), .C1 (n_137_81), .C2 (n_134_81) );
AOI211_X1 g_146_78 (.ZN (n_146_78), .A (n_143_77), .B (n_143_78), .C1 (n_139_80), .C2 (n_136_80) );
AOI211_X1 g_144_79 (.ZN (n_144_79), .A (n_145_76), .B (n_142_80), .C1 (n_141_79), .C2 (n_135_82) );
AOI211_X1 g_146_80 (.ZN (n_146_80), .A (n_146_78), .B (n_141_78), .C1 (n_143_78), .C2 (n_137_81) );
AOI211_X1 g_148_79 (.ZN (n_148_79), .A (n_144_79), .B (n_143_77), .C1 (n_142_80), .C2 (n_139_80) );
AOI211_X1 g_147_77 (.ZN (n_147_77), .A (n_146_80), .B (n_145_76), .C1 (n_141_78), .C2 (n_141_79) );
AOI211_X1 g_145_78 (.ZN (n_145_78), .A (n_148_79), .B (n_146_78), .C1 (n_143_77), .C2 (n_143_78) );
AOI211_X1 g_143_79 (.ZN (n_143_79), .A (n_147_77), .B (n_144_79), .C1 (n_145_76), .C2 (n_142_80) );
AOI211_X1 g_144_81 (.ZN (n_144_81), .A (n_145_78), .B (n_146_80), .C1 (n_146_78), .C2 (n_141_78) );
AOI211_X1 g_146_82 (.ZN (n_146_82), .A (n_143_79), .B (n_148_79), .C1 (n_144_79), .C2 (n_143_77) );
AOI211_X1 g_148_83 (.ZN (n_148_83), .A (n_144_81), .B (n_147_77), .C1 (n_146_80), .C2 (n_145_76) );
AOI211_X1 g_147_81 (.ZN (n_147_81), .A (n_146_82), .B (n_145_78), .C1 (n_148_79), .C2 (n_146_78) );
AOI211_X1 g_146_79 (.ZN (n_146_79), .A (n_148_83), .B (n_143_79), .C1 (n_147_77), .C2 (n_144_79) );
AOI211_X1 g_144_78 (.ZN (n_144_78), .A (n_147_81), .B (n_144_81), .C1 (n_145_78), .C2 (n_146_80) );
AOI211_X1 g_145_80 (.ZN (n_145_80), .A (n_146_79), .B (n_146_82), .C1 (n_143_79), .C2 (n_148_79) );
AOI211_X1 g_143_81 (.ZN (n_143_81), .A (n_144_78), .B (n_148_83), .C1 (n_144_81), .C2 (n_147_77) );
AOI211_X1 g_142_79 (.ZN (n_142_79), .A (n_145_80), .B (n_147_81), .C1 (n_146_82), .C2 (n_145_78) );
AOI211_X1 g_144_80 (.ZN (n_144_80), .A (n_143_81), .B (n_146_79), .C1 (n_148_83), .C2 (n_143_79) );
AOI211_X1 g_145_82 (.ZN (n_145_82), .A (n_142_79), .B (n_144_78), .C1 (n_147_81), .C2 (n_144_81) );
AOI211_X1 g_146_84 (.ZN (n_146_84), .A (n_144_80), .B (n_145_80), .C1 (n_146_79), .C2 (n_146_82) );
AOI211_X1 g_144_83 (.ZN (n_144_83), .A (n_145_82), .B (n_143_81), .C1 (n_144_78), .C2 (n_148_83) );
AOI211_X1 g_145_81 (.ZN (n_145_81), .A (n_146_84), .B (n_142_79), .C1 (n_145_80), .C2 (n_147_81) );
AOI211_X1 g_143_80 (.ZN (n_143_80), .A (n_144_83), .B (n_144_80), .C1 (n_143_81), .C2 (n_146_79) );
AOI211_X1 g_141_81 (.ZN (n_141_81), .A (n_145_81), .B (n_145_82), .C1 (n_142_79), .C2 (n_144_78) );
AOI211_X1 g_143_82 (.ZN (n_143_82), .A (n_143_80), .B (n_146_84), .C1 (n_144_80), .C2 (n_145_80) );
AOI211_X1 g_144_84 (.ZN (n_144_84), .A (n_141_81), .B (n_144_83), .C1 (n_145_82), .C2 (n_143_81) );
AOI211_X1 g_146_83 (.ZN (n_146_83), .A (n_143_82), .B (n_145_81), .C1 (n_146_84), .C2 (n_142_79) );
AOI211_X1 g_144_82 (.ZN (n_144_82), .A (n_144_84), .B (n_143_80), .C1 (n_144_83), .C2 (n_144_80) );
AOI211_X1 g_142_81 (.ZN (n_142_81), .A (n_146_83), .B (n_141_81), .C1 (n_145_81), .C2 (n_145_82) );
AOI211_X1 g_140_80 (.ZN (n_140_80), .A (n_144_82), .B (n_143_82), .C1 (n_143_80), .C2 (n_146_84) );
AOI211_X1 g_139_82 (.ZN (n_139_82), .A (n_142_81), .B (n_144_84), .C1 (n_141_81), .C2 (n_144_83) );
AOI211_X1 g_137_83 (.ZN (n_137_83), .A (n_140_80), .B (n_146_83), .C1 (n_143_82), .C2 (n_145_81) );
AOI211_X1 g_138_81 (.ZN (n_138_81), .A (n_139_82), .B (n_144_82), .C1 (n_144_84), .C2 (n_143_80) );
AOI211_X1 g_139_79 (.ZN (n_139_79), .A (n_137_83), .B (n_142_81), .C1 (n_146_83), .C2 (n_141_81) );
AOI211_X1 g_137_80 (.ZN (n_137_80), .A (n_138_81), .B (n_140_80), .C1 (n_144_82), .C2 (n_143_82) );
AOI211_X1 g_136_82 (.ZN (n_136_82), .A (n_139_79), .B (n_139_82), .C1 (n_142_81), .C2 (n_144_84) );
AOI211_X1 g_134_83 (.ZN (n_134_83), .A (n_137_80), .B (n_137_83), .C1 (n_140_80), .C2 (n_146_83) );
AOI211_X1 g_132_84 (.ZN (n_132_84), .A (n_136_82), .B (n_138_81), .C1 (n_139_82), .C2 (n_144_82) );
AOI211_X1 g_130_85 (.ZN (n_130_85), .A (n_134_83), .B (n_139_79), .C1 (n_137_83), .C2 (n_142_81) );
AOI211_X1 g_128_86 (.ZN (n_128_86), .A (n_132_84), .B (n_137_80), .C1 (n_138_81), .C2 (n_140_80) );
AOI211_X1 g_126_87 (.ZN (n_126_87), .A (n_130_85), .B (n_136_82), .C1 (n_139_79), .C2 (n_139_82) );
AOI211_X1 g_125_89 (.ZN (n_125_89), .A (n_128_86), .B (n_134_83), .C1 (n_137_80), .C2 (n_137_83) );
AOI211_X1 g_123_88 (.ZN (n_123_88), .A (n_126_87), .B (n_132_84), .C1 (n_136_82), .C2 (n_138_81) );
AOI211_X1 g_125_87 (.ZN (n_125_87), .A (n_125_89), .B (n_130_85), .C1 (n_134_83), .C2 (n_139_79) );
AOI211_X1 g_127_86 (.ZN (n_127_86), .A (n_123_88), .B (n_128_86), .C1 (n_132_84), .C2 (n_137_80) );
AOI211_X1 g_129_85 (.ZN (n_129_85), .A (n_125_87), .B (n_126_87), .C1 (n_130_85), .C2 (n_136_82) );
AOI211_X1 g_131_84 (.ZN (n_131_84), .A (n_127_86), .B (n_125_89), .C1 (n_128_86), .C2 (n_134_83) );
AOI211_X1 g_133_83 (.ZN (n_133_83), .A (n_129_85), .B (n_123_88), .C1 (n_126_87), .C2 (n_132_84) );
AOI211_X1 g_135_84 (.ZN (n_135_84), .A (n_131_84), .B (n_125_87), .C1 (n_125_89), .C2 (n_130_85) );
AOI211_X1 g_133_85 (.ZN (n_133_85), .A (n_133_83), .B (n_127_86), .C1 (n_123_88), .C2 (n_128_86) );
AOI211_X1 g_131_86 (.ZN (n_131_86), .A (n_135_84), .B (n_129_85), .C1 (n_125_87), .C2 (n_126_87) );
AOI211_X1 g_129_87 (.ZN (n_129_87), .A (n_133_85), .B (n_131_84), .C1 (n_127_86), .C2 (n_125_89) );
AOI211_X1 g_127_88 (.ZN (n_127_88), .A (n_131_86), .B (n_133_83), .C1 (n_129_85), .C2 (n_123_88) );
AOI211_X1 g_126_90 (.ZN (n_126_90), .A (n_129_87), .B (n_135_84), .C1 (n_131_84), .C2 (n_125_87) );
AOI211_X1 g_124_89 (.ZN (n_124_89), .A (n_127_88), .B (n_133_85), .C1 (n_133_83), .C2 (n_127_86) );
AOI211_X1 g_126_88 (.ZN (n_126_88), .A (n_126_90), .B (n_131_86), .C1 (n_135_84), .C2 (n_129_85) );
AOI211_X1 g_128_87 (.ZN (n_128_87), .A (n_124_89), .B (n_129_87), .C1 (n_133_85), .C2 (n_131_84) );
AOI211_X1 g_130_86 (.ZN (n_130_86), .A (n_126_88), .B (n_127_88), .C1 (n_131_86), .C2 (n_133_83) );
AOI211_X1 g_132_85 (.ZN (n_132_85), .A (n_128_87), .B (n_126_90), .C1 (n_129_87), .C2 (n_135_84) );
AOI211_X1 g_134_84 (.ZN (n_134_84), .A (n_130_86), .B (n_124_89), .C1 (n_127_88), .C2 (n_133_85) );
AOI211_X1 g_136_83 (.ZN (n_136_83), .A (n_132_85), .B (n_126_88), .C1 (n_126_90), .C2 (n_131_86) );
AOI211_X1 g_138_82 (.ZN (n_138_82), .A (n_134_84), .B (n_128_87), .C1 (n_124_89), .C2 (n_129_87) );
AOI211_X1 g_140_81 (.ZN (n_140_81), .A (n_136_83), .B (n_130_86), .C1 (n_126_88), .C2 (n_127_88) );
AOI211_X1 g_141_83 (.ZN (n_141_83), .A (n_138_82), .B (n_132_85), .C1 (n_128_87), .C2 (n_126_90) );
AOI211_X1 g_139_84 (.ZN (n_139_84), .A (n_140_81), .B (n_134_84), .C1 (n_130_86), .C2 (n_124_89) );
AOI211_X1 g_140_82 (.ZN (n_140_82), .A (n_141_83), .B (n_136_83), .C1 (n_132_85), .C2 (n_126_88) );
AOI211_X1 g_141_80 (.ZN (n_141_80), .A (n_139_84), .B (n_138_82), .C1 (n_134_84), .C2 (n_128_87) );
AOI211_X1 g_142_82 (.ZN (n_142_82), .A (n_140_82), .B (n_140_81), .C1 (n_136_83), .C2 (n_130_86) );
AOI211_X1 g_143_84 (.ZN (n_143_84), .A (n_141_80), .B (n_141_83), .C1 (n_138_82), .C2 (n_132_85) );
AOI211_X1 g_145_85 (.ZN (n_145_85), .A (n_142_82), .B (n_139_84), .C1 (n_140_81), .C2 (n_134_84) );
AOI211_X1 g_143_86 (.ZN (n_143_86), .A (n_143_84), .B (n_140_82), .C1 (n_141_83), .C2 (n_136_83) );
AOI211_X1 g_142_84 (.ZN (n_142_84), .A (n_145_85), .B (n_141_80), .C1 (n_139_84), .C2 (n_138_82) );
AOI211_X1 g_141_82 (.ZN (n_141_82), .A (n_143_86), .B (n_142_82), .C1 (n_140_82), .C2 (n_140_81) );
AOI211_X1 g_139_81 (.ZN (n_139_81), .A (n_142_84), .B (n_143_84), .C1 (n_141_80), .C2 (n_141_83) );
AOI211_X1 g_140_83 (.ZN (n_140_83), .A (n_141_82), .B (n_145_85), .C1 (n_142_82), .C2 (n_139_84) );
AOI211_X1 g_141_85 (.ZN (n_141_85), .A (n_139_81), .B (n_143_86), .C1 (n_143_84), .C2 (n_140_82) );
AOI211_X1 g_142_83 (.ZN (n_142_83), .A (n_140_83), .B (n_142_84), .C1 (n_145_85), .C2 (n_141_80) );
AOI211_X1 g_140_84 (.ZN (n_140_84), .A (n_141_85), .B (n_141_82), .C1 (n_143_86), .C2 (n_142_82) );
AOI211_X1 g_138_83 (.ZN (n_138_83), .A (n_142_83), .B (n_139_81), .C1 (n_142_84), .C2 (n_143_84) );
AOI211_X1 g_137_85 (.ZN (n_137_85), .A (n_140_84), .B (n_140_83), .C1 (n_141_82), .C2 (n_145_85) );
AOI211_X1 g_135_86 (.ZN (n_135_86), .A (n_138_83), .B (n_141_85), .C1 (n_139_81), .C2 (n_143_86) );
AOI211_X1 g_136_84 (.ZN (n_136_84), .A (n_137_85), .B (n_142_83), .C1 (n_140_83), .C2 (n_142_84) );
AOI211_X1 g_137_82 (.ZN (n_137_82), .A (n_135_86), .B (n_140_84), .C1 (n_141_85), .C2 (n_141_82) );
AOI211_X1 g_135_83 (.ZN (n_135_83), .A (n_136_84), .B (n_138_83), .C1 (n_142_83), .C2 (n_139_81) );
AOI211_X1 g_133_84 (.ZN (n_133_84), .A (n_137_82), .B (n_137_85), .C1 (n_140_84), .C2 (n_140_83) );
AOI211_X1 g_131_85 (.ZN (n_131_85), .A (n_135_83), .B (n_135_86), .C1 (n_138_83), .C2 (n_141_85) );
AOI211_X1 g_130_87 (.ZN (n_130_87), .A (n_133_84), .B (n_136_84), .C1 (n_137_85), .C2 (n_142_83) );
AOI211_X1 g_132_86 (.ZN (n_132_86), .A (n_131_85), .B (n_137_82), .C1 (n_135_86), .C2 (n_140_84) );
AOI211_X1 g_134_85 (.ZN (n_134_85), .A (n_130_87), .B (n_135_83), .C1 (n_136_84), .C2 (n_138_83) );
AOI211_X1 g_133_87 (.ZN (n_133_87), .A (n_132_86), .B (n_133_84), .C1 (n_137_82), .C2 (n_137_85) );
AOI211_X1 g_131_88 (.ZN (n_131_88), .A (n_134_85), .B (n_131_85), .C1 (n_135_83), .C2 (n_135_86) );
AOI211_X1 g_129_89 (.ZN (n_129_89), .A (n_133_87), .B (n_130_87), .C1 (n_133_84), .C2 (n_136_84) );
AOI211_X1 g_127_90 (.ZN (n_127_90), .A (n_131_88), .B (n_132_86), .C1 (n_131_85), .C2 (n_137_82) );
AOI211_X1 g_128_88 (.ZN (n_128_88), .A (n_129_89), .B (n_134_85), .C1 (n_130_87), .C2 (n_135_83) );
AOI211_X1 g_126_89 (.ZN (n_126_89), .A (n_127_90), .B (n_133_87), .C1 (n_132_86), .C2 (n_133_84) );
AOI211_X1 g_124_90 (.ZN (n_124_90), .A (n_128_88), .B (n_131_88), .C1 (n_134_85), .C2 (n_131_85) );
AOI211_X1 g_122_91 (.ZN (n_122_91), .A (n_126_89), .B (n_129_89), .C1 (n_133_87), .C2 (n_130_87) );
AOI211_X1 g_121_89 (.ZN (n_121_89), .A (n_124_90), .B (n_127_90), .C1 (n_131_88), .C2 (n_132_86) );
AOI211_X1 g_119_90 (.ZN (n_119_90), .A (n_122_91), .B (n_128_88), .C1 (n_129_89), .C2 (n_134_85) );
AOI211_X1 g_117_91 (.ZN (n_117_91), .A (n_121_89), .B (n_126_89), .C1 (n_127_90), .C2 (n_133_87) );
AOI211_X1 g_115_92 (.ZN (n_115_92), .A (n_119_90), .B (n_124_90), .C1 (n_128_88), .C2 (n_131_88) );
AOI211_X1 g_113_93 (.ZN (n_113_93), .A (n_117_91), .B (n_122_91), .C1 (n_126_89), .C2 (n_129_89) );
AOI211_X1 g_111_94 (.ZN (n_111_94), .A (n_115_92), .B (n_121_89), .C1 (n_124_90), .C2 (n_127_90) );
AOI211_X1 g_109_95 (.ZN (n_109_95), .A (n_113_93), .B (n_119_90), .C1 (n_122_91), .C2 (n_128_88) );
AOI211_X1 g_108_97 (.ZN (n_108_97), .A (n_111_94), .B (n_117_91), .C1 (n_121_89), .C2 (n_126_89) );
AOI211_X1 g_106_96 (.ZN (n_106_96), .A (n_109_95), .B (n_115_92), .C1 (n_119_90), .C2 (n_124_90) );
AOI211_X1 g_108_95 (.ZN (n_108_95), .A (n_108_97), .B (n_113_93), .C1 (n_117_91), .C2 (n_122_91) );
AOI211_X1 g_110_94 (.ZN (n_110_94), .A (n_106_96), .B (n_111_94), .C1 (n_115_92), .C2 (n_121_89) );
AOI211_X1 g_112_93 (.ZN (n_112_93), .A (n_108_95), .B (n_109_95), .C1 (n_113_93), .C2 (n_119_90) );
AOI211_X1 g_114_92 (.ZN (n_114_92), .A (n_110_94), .B (n_108_97), .C1 (n_111_94), .C2 (n_117_91) );
AOI211_X1 g_116_91 (.ZN (n_116_91), .A (n_112_93), .B (n_106_96), .C1 (n_109_95), .C2 (n_115_92) );
AOI211_X1 g_117_93 (.ZN (n_117_93), .A (n_114_92), .B (n_108_95), .C1 (n_108_97), .C2 (n_113_93) );
AOI211_X1 g_115_94 (.ZN (n_115_94), .A (n_116_91), .B (n_110_94), .C1 (n_106_96), .C2 (n_111_94) );
AOI211_X1 g_113_95 (.ZN (n_113_95), .A (n_117_93), .B (n_112_93), .C1 (n_108_95), .C2 (n_109_95) );
AOI211_X1 g_111_96 (.ZN (n_111_96), .A (n_115_94), .B (n_114_92), .C1 (n_110_94), .C2 (n_108_97) );
AOI211_X1 g_109_97 (.ZN (n_109_97), .A (n_113_95), .B (n_116_91), .C1 (n_112_93), .C2 (n_106_96) );
AOI211_X1 g_107_98 (.ZN (n_107_98), .A (n_111_96), .B (n_117_93), .C1 (n_114_92), .C2 (n_108_95) );
AOI211_X1 g_105_99 (.ZN (n_105_99), .A (n_109_97), .B (n_115_94), .C1 (n_116_91), .C2 (n_110_94) );
AOI211_X1 g_106_97 (.ZN (n_106_97), .A (n_107_98), .B (n_113_95), .C1 (n_117_93), .C2 (n_112_93) );
AOI211_X1 g_104_98 (.ZN (n_104_98), .A (n_105_99), .B (n_111_96), .C1 (n_115_94), .C2 (n_114_92) );
AOI211_X1 g_102_99 (.ZN (n_102_99), .A (n_106_97), .B (n_109_97), .C1 (n_113_95), .C2 (n_116_91) );
AOI211_X1 g_100_98 (.ZN (n_100_98), .A (n_104_98), .B (n_107_98), .C1 (n_111_96), .C2 (n_117_93) );
AOI211_X1 g_98_99 (.ZN (n_98_99), .A (n_102_99), .B (n_105_99), .C1 (n_109_97), .C2 (n_115_94) );
AOI211_X1 g_100_100 (.ZN (n_100_100), .A (n_100_98), .B (n_106_97), .C1 (n_107_98), .C2 (n_113_95) );
AOI211_X1 g_101_98 (.ZN (n_101_98), .A (n_98_99), .B (n_104_98), .C1 (n_105_99), .C2 (n_111_96) );
AOI211_X1 g_99_99 (.ZN (n_99_99), .A (n_100_100), .B (n_102_99), .C1 (n_106_97), .C2 (n_109_97) );
AOI211_X1 g_98_101 (.ZN (n_98_101), .A (n_101_98), .B (n_100_98), .C1 (n_104_98), .C2 (n_107_98) );
AOI211_X1 g_97_99 (.ZN (n_97_99), .A (n_99_99), .B (n_98_99), .C1 (n_102_99), .C2 (n_105_99) );
AOI211_X1 g_99_98 (.ZN (n_99_98), .A (n_98_101), .B (n_100_100), .C1 (n_100_98), .C2 (n_106_97) );
AOI211_X1 g_101_99 (.ZN (n_101_99), .A (n_97_99), .B (n_101_98), .C1 (n_98_99), .C2 (n_104_98) );
AOI211_X1 g_99_100 (.ZN (n_99_100), .A (n_99_98), .B (n_99_99), .C1 (n_100_100), .C2 (n_102_99) );
AOI211_X1 g_98_98 (.ZN (n_98_98), .A (n_101_99), .B (n_98_101), .C1 (n_101_98), .C2 (n_100_98) );
AOI211_X1 g_96_97 (.ZN (n_96_97), .A (n_99_100), .B (n_97_99), .C1 (n_99_99), .C2 (n_98_99) );
AOI211_X1 g_95_99 (.ZN (n_95_99), .A (n_98_98), .B (n_99_98), .C1 (n_98_101), .C2 (n_100_100) );
AOI211_X1 g_93_100 (.ZN (n_93_100), .A (n_96_97), .B (n_101_99), .C1 (n_97_99), .C2 (n_101_98) );
AOI211_X1 g_94_98 (.ZN (n_94_98), .A (n_95_99), .B (n_99_100), .C1 (n_99_98), .C2 (n_99_99) );
AOI211_X1 g_92_99 (.ZN (n_92_99), .A (n_93_100), .B (n_98_98), .C1 (n_101_99), .C2 (n_98_101) );
AOI211_X1 g_91_101 (.ZN (n_91_101), .A (n_94_98), .B (n_96_97), .C1 (n_99_100), .C2 (n_97_99) );
AOI211_X1 g_89_102 (.ZN (n_89_102), .A (n_92_99), .B (n_95_99), .C1 (n_98_98), .C2 (n_99_98) );
AOI211_X1 g_90_100 (.ZN (n_90_100), .A (n_91_101), .B (n_93_100), .C1 (n_96_97), .C2 (n_101_99) );
AOI211_X1 g_88_101 (.ZN (n_88_101), .A (n_89_102), .B (n_94_98), .C1 (n_95_99), .C2 (n_99_100) );
AOI211_X1 g_87_103 (.ZN (n_87_103), .A (n_90_100), .B (n_92_99), .C1 (n_93_100), .C2 (n_98_98) );
AOI211_X1 g_85_104 (.ZN (n_85_104), .A (n_88_101), .B (n_91_101), .C1 (n_94_98), .C2 (n_96_97) );
AOI211_X1 g_86_102 (.ZN (n_86_102), .A (n_87_103), .B (n_89_102), .C1 (n_92_99), .C2 (n_95_99) );
AOI211_X1 g_84_103 (.ZN (n_84_103), .A (n_85_104), .B (n_90_100), .C1 (n_91_101), .C2 (n_93_100) );
AOI211_X1 g_83_105 (.ZN (n_83_105), .A (n_86_102), .B (n_88_101), .C1 (n_89_102), .C2 (n_94_98) );
AOI211_X1 g_81_106 (.ZN (n_81_106), .A (n_84_103), .B (n_87_103), .C1 (n_90_100), .C2 (n_92_99) );
AOI211_X1 g_80_108 (.ZN (n_80_108), .A (n_83_105), .B (n_85_104), .C1 (n_88_101), .C2 (n_91_101) );
AOI211_X1 g_78_109 (.ZN (n_78_109), .A (n_81_106), .B (n_86_102), .C1 (n_87_103), .C2 (n_89_102) );
AOI211_X1 g_77_107 (.ZN (n_77_107), .A (n_80_108), .B (n_84_103), .C1 (n_85_104), .C2 (n_90_100) );
AOI211_X1 g_75_108 (.ZN (n_75_108), .A (n_78_109), .B (n_83_105), .C1 (n_86_102), .C2 (n_88_101) );
AOI211_X1 g_73_109 (.ZN (n_73_109), .A (n_77_107), .B (n_81_106), .C1 (n_84_103), .C2 (n_87_103) );
AOI211_X1 g_74_107 (.ZN (n_74_107), .A (n_75_108), .B (n_80_108), .C1 (n_83_105), .C2 (n_85_104) );
AOI211_X1 g_76_108 (.ZN (n_76_108), .A (n_73_109), .B (n_78_109), .C1 (n_81_106), .C2 (n_86_102) );
AOI211_X1 g_74_109 (.ZN (n_74_109), .A (n_74_107), .B (n_77_107), .C1 (n_80_108), .C2 (n_84_103) );
AOI211_X1 g_72_108 (.ZN (n_72_108), .A (n_76_108), .B (n_75_108), .C1 (n_78_109), .C2 (n_83_105) );
AOI211_X1 g_70_109 (.ZN (n_70_109), .A (n_74_109), .B (n_73_109), .C1 (n_77_107), .C2 (n_81_106) );
AOI211_X1 g_72_110 (.ZN (n_72_110), .A (n_72_108), .B (n_74_107), .C1 (n_75_108), .C2 (n_80_108) );
AOI211_X1 g_70_111 (.ZN (n_70_111), .A (n_70_109), .B (n_76_108), .C1 (n_73_109), .C2 (n_78_109) );
AOI211_X1 g_68_112 (.ZN (n_68_112), .A (n_72_110), .B (n_74_109), .C1 (n_74_107), .C2 (n_77_107) );
AOI211_X1 g_66_113 (.ZN (n_66_113), .A (n_70_111), .B (n_72_108), .C1 (n_76_108), .C2 (n_75_108) );
AOI211_X1 g_64_114 (.ZN (n_64_114), .A (n_68_112), .B (n_70_109), .C1 (n_74_109), .C2 (n_73_109) );
AOI211_X1 g_62_115 (.ZN (n_62_115), .A (n_66_113), .B (n_72_110), .C1 (n_72_108), .C2 (n_74_107) );
AOI211_X1 g_60_116 (.ZN (n_60_116), .A (n_64_114), .B (n_70_111), .C1 (n_70_109), .C2 (n_76_108) );
AOI211_X1 g_58_117 (.ZN (n_58_117), .A (n_62_115), .B (n_68_112), .C1 (n_72_110), .C2 (n_74_109) );
AOI211_X1 g_56_118 (.ZN (n_56_118), .A (n_60_116), .B (n_66_113), .C1 (n_70_111), .C2 (n_72_108) );
AOI211_X1 g_57_116 (.ZN (n_57_116), .A (n_58_117), .B (n_64_114), .C1 (n_68_112), .C2 (n_70_109) );
AOI211_X1 g_55_117 (.ZN (n_55_117), .A (n_56_118), .B (n_62_115), .C1 (n_66_113), .C2 (n_72_110) );
AOI211_X1 g_53_118 (.ZN (n_53_118), .A (n_57_116), .B (n_60_116), .C1 (n_64_114), .C2 (n_70_111) );
AOI211_X1 g_51_119 (.ZN (n_51_119), .A (n_55_117), .B (n_58_117), .C1 (n_62_115), .C2 (n_68_112) );
AOI211_X1 g_49_120 (.ZN (n_49_120), .A (n_53_118), .B (n_56_118), .C1 (n_60_116), .C2 (n_66_113) );
AOI211_X1 g_47_121 (.ZN (n_47_121), .A (n_51_119), .B (n_57_116), .C1 (n_58_117), .C2 (n_64_114) );
AOI211_X1 g_45_122 (.ZN (n_45_122), .A (n_49_120), .B (n_55_117), .C1 (n_56_118), .C2 (n_62_115) );
AOI211_X1 g_43_123 (.ZN (n_43_123), .A (n_47_121), .B (n_53_118), .C1 (n_57_116), .C2 (n_60_116) );
AOI211_X1 g_41_124 (.ZN (n_41_124), .A (n_45_122), .B (n_51_119), .C1 (n_55_117), .C2 (n_58_117) );
AOI211_X1 g_39_125 (.ZN (n_39_125), .A (n_43_123), .B (n_49_120), .C1 (n_53_118), .C2 (n_56_118) );
AOI211_X1 g_37_126 (.ZN (n_37_126), .A (n_41_124), .B (n_47_121), .C1 (n_51_119), .C2 (n_57_116) );
AOI211_X1 g_35_127 (.ZN (n_35_127), .A (n_39_125), .B (n_45_122), .C1 (n_49_120), .C2 (n_55_117) );
AOI211_X1 g_33_128 (.ZN (n_33_128), .A (n_37_126), .B (n_43_123), .C1 (n_47_121), .C2 (n_53_118) );
AOI211_X1 g_31_129 (.ZN (n_31_129), .A (n_35_127), .B (n_41_124), .C1 (n_45_122), .C2 (n_51_119) );
AOI211_X1 g_30_131 (.ZN (n_30_131), .A (n_33_128), .B (n_39_125), .C1 (n_43_123), .C2 (n_49_120) );
AOI211_X1 g_32_130 (.ZN (n_32_130), .A (n_31_129), .B (n_37_126), .C1 (n_41_124), .C2 (n_47_121) );
AOI211_X1 g_34_129 (.ZN (n_34_129), .A (n_30_131), .B (n_35_127), .C1 (n_39_125), .C2 (n_45_122) );
AOI211_X1 g_36_128 (.ZN (n_36_128), .A (n_32_130), .B (n_33_128), .C1 (n_37_126), .C2 (n_43_123) );
AOI211_X1 g_38_127 (.ZN (n_38_127), .A (n_34_129), .B (n_31_129), .C1 (n_35_127), .C2 (n_41_124) );
AOI211_X1 g_40_126 (.ZN (n_40_126), .A (n_36_128), .B (n_30_131), .C1 (n_33_128), .C2 (n_39_125) );
AOI211_X1 g_42_125 (.ZN (n_42_125), .A (n_38_127), .B (n_32_130), .C1 (n_31_129), .C2 (n_37_126) );
AOI211_X1 g_44_124 (.ZN (n_44_124), .A (n_40_126), .B (n_34_129), .C1 (n_30_131), .C2 (n_35_127) );
AOI211_X1 g_46_123 (.ZN (n_46_123), .A (n_42_125), .B (n_36_128), .C1 (n_32_130), .C2 (n_33_128) );
AOI211_X1 g_48_122 (.ZN (n_48_122), .A (n_44_124), .B (n_38_127), .C1 (n_34_129), .C2 (n_31_129) );
AOI211_X1 g_50_121 (.ZN (n_50_121), .A (n_46_123), .B (n_40_126), .C1 (n_36_128), .C2 (n_30_131) );
AOI211_X1 g_52_120 (.ZN (n_52_120), .A (n_48_122), .B (n_42_125), .C1 (n_38_127), .C2 (n_32_130) );
AOI211_X1 g_54_119 (.ZN (n_54_119), .A (n_50_121), .B (n_44_124), .C1 (n_40_126), .C2 (n_34_129) );
AOI211_X1 g_53_121 (.ZN (n_53_121), .A (n_52_120), .B (n_46_123), .C1 (n_42_125), .C2 (n_36_128) );
AOI211_X1 g_55_120 (.ZN (n_55_120), .A (n_54_119), .B (n_48_122), .C1 (n_44_124), .C2 (n_38_127) );
AOI211_X1 g_57_119 (.ZN (n_57_119), .A (n_53_121), .B (n_50_121), .C1 (n_46_123), .C2 (n_40_126) );
AOI211_X1 g_59_118 (.ZN (n_59_118), .A (n_55_120), .B (n_52_120), .C1 (n_48_122), .C2 (n_42_125) );
AOI211_X1 g_61_117 (.ZN (n_61_117), .A (n_57_119), .B (n_54_119), .C1 (n_50_121), .C2 (n_44_124) );
AOI211_X1 g_63_116 (.ZN (n_63_116), .A (n_59_118), .B (n_53_121), .C1 (n_52_120), .C2 (n_46_123) );
AOI211_X1 g_65_115 (.ZN (n_65_115), .A (n_61_117), .B (n_55_120), .C1 (n_54_119), .C2 (n_48_122) );
AOI211_X1 g_67_114 (.ZN (n_67_114), .A (n_63_116), .B (n_57_119), .C1 (n_53_121), .C2 (n_50_121) );
AOI211_X1 g_69_113 (.ZN (n_69_113), .A (n_65_115), .B (n_59_118), .C1 (n_55_120), .C2 (n_52_120) );
AOI211_X1 g_67_112 (.ZN (n_67_112), .A (n_67_114), .B (n_61_117), .C1 (n_57_119), .C2 (n_54_119) );
AOI211_X1 g_69_111 (.ZN (n_69_111), .A (n_69_113), .B (n_63_116), .C1 (n_59_118), .C2 (n_53_121) );
AOI211_X1 g_71_110 (.ZN (n_71_110), .A (n_67_112), .B (n_65_115), .C1 (n_61_117), .C2 (n_55_120) );
AOI211_X1 g_70_112 (.ZN (n_70_112), .A (n_69_111), .B (n_67_114), .C1 (n_63_116), .C2 (n_57_119) );
AOI211_X1 g_72_111 (.ZN (n_72_111), .A (n_71_110), .B (n_69_113), .C1 (n_65_115), .C2 (n_59_118) );
AOI211_X1 g_74_110 (.ZN (n_74_110), .A (n_70_112), .B (n_67_112), .C1 (n_67_114), .C2 (n_61_117) );
AOI211_X1 g_76_109 (.ZN (n_76_109), .A (n_72_111), .B (n_69_111), .C1 (n_69_113), .C2 (n_63_116) );
AOI211_X1 g_78_108 (.ZN (n_78_108), .A (n_74_110), .B (n_71_110), .C1 (n_67_112), .C2 (n_65_115) );
AOI211_X1 g_80_107 (.ZN (n_80_107), .A (n_76_109), .B (n_70_112), .C1 (n_69_111), .C2 (n_67_114) );
AOI211_X1 g_78_106 (.ZN (n_78_106), .A (n_78_108), .B (n_72_111), .C1 (n_71_110), .C2 (n_69_113) );
AOI211_X1 g_80_105 (.ZN (n_80_105), .A (n_80_107), .B (n_74_110), .C1 (n_70_112), .C2 (n_67_112) );
AOI211_X1 g_79_107 (.ZN (n_79_107), .A (n_78_106), .B (n_76_109), .C1 (n_72_111), .C2 (n_69_111) );
AOI211_X1 g_77_108 (.ZN (n_77_108), .A (n_80_105), .B (n_78_108), .C1 (n_74_110), .C2 (n_71_110) );
AOI211_X1 g_75_109 (.ZN (n_75_109), .A (n_79_107), .B (n_80_107), .C1 (n_76_109), .C2 (n_70_112) );
AOI211_X1 g_73_110 (.ZN (n_73_110), .A (n_77_108), .B (n_78_106), .C1 (n_78_108), .C2 (n_72_111) );
AOI211_X1 g_71_111 (.ZN (n_71_111), .A (n_75_109), .B (n_80_105), .C1 (n_80_107), .C2 (n_74_110) );
AOI211_X1 g_69_112 (.ZN (n_69_112), .A (n_73_110), .B (n_79_107), .C1 (n_78_106), .C2 (n_76_109) );
AOI211_X1 g_67_113 (.ZN (n_67_113), .A (n_71_111), .B (n_77_108), .C1 (n_80_105), .C2 (n_78_108) );
AOI211_X1 g_65_114 (.ZN (n_65_114), .A (n_69_112), .B (n_75_109), .C1 (n_79_107), .C2 (n_80_107) );
AOI211_X1 g_63_115 (.ZN (n_63_115), .A (n_67_113), .B (n_73_110), .C1 (n_77_108), .C2 (n_78_106) );
AOI211_X1 g_62_117 (.ZN (n_62_117), .A (n_65_114), .B (n_71_111), .C1 (n_75_109), .C2 (n_80_105) );
AOI211_X1 g_64_116 (.ZN (n_64_116), .A (n_63_115), .B (n_69_112), .C1 (n_73_110), .C2 (n_79_107) );
AOI211_X1 g_66_115 (.ZN (n_66_115), .A (n_62_117), .B (n_67_113), .C1 (n_71_111), .C2 (n_77_108) );
AOI211_X1 g_68_114 (.ZN (n_68_114), .A (n_64_116), .B (n_65_114), .C1 (n_69_112), .C2 (n_75_109) );
AOI211_X1 g_70_113 (.ZN (n_70_113), .A (n_66_115), .B (n_63_115), .C1 (n_67_113), .C2 (n_73_110) );
AOI211_X1 g_72_112 (.ZN (n_72_112), .A (n_68_114), .B (n_62_117), .C1 (n_65_114), .C2 (n_71_111) );
AOI211_X1 g_74_111 (.ZN (n_74_111), .A (n_70_113), .B (n_64_116), .C1 (n_63_115), .C2 (n_69_112) );
AOI211_X1 g_76_110 (.ZN (n_76_110), .A (n_72_112), .B (n_66_115), .C1 (n_62_117), .C2 (n_67_113) );
AOI211_X1 g_75_112 (.ZN (n_75_112), .A (n_74_111), .B (n_68_114), .C1 (n_64_116), .C2 (n_65_114) );
AOI211_X1 g_73_111 (.ZN (n_73_111), .A (n_76_110), .B (n_70_113), .C1 (n_66_115), .C2 (n_63_115) );
AOI211_X1 g_71_112 (.ZN (n_71_112), .A (n_75_112), .B (n_72_112), .C1 (n_68_114), .C2 (n_62_117) );
AOI211_X1 g_73_113 (.ZN (n_73_113), .A (n_73_111), .B (n_74_111), .C1 (n_70_113), .C2 (n_64_116) );
AOI211_X1 g_71_114 (.ZN (n_71_114), .A (n_71_112), .B (n_76_110), .C1 (n_72_112), .C2 (n_66_115) );
AOI211_X1 g_69_115 (.ZN (n_69_115), .A (n_73_113), .B (n_75_112), .C1 (n_74_111), .C2 (n_68_114) );
AOI211_X1 g_68_113 (.ZN (n_68_113), .A (n_71_114), .B (n_73_111), .C1 (n_76_110), .C2 (n_70_113) );
AOI211_X1 g_66_114 (.ZN (n_66_114), .A (n_69_115), .B (n_71_112), .C1 (n_75_112), .C2 (n_72_112) );
AOI211_X1 g_64_115 (.ZN (n_64_115), .A (n_68_113), .B (n_73_113), .C1 (n_73_111), .C2 (n_74_111) );
AOI211_X1 g_62_116 (.ZN (n_62_116), .A (n_66_114), .B (n_71_114), .C1 (n_71_112), .C2 (n_76_110) );
AOI211_X1 g_60_117 (.ZN (n_60_117), .A (n_64_115), .B (n_69_115), .C1 (n_73_113), .C2 (n_75_112) );
AOI211_X1 g_58_118 (.ZN (n_58_118), .A (n_62_116), .B (n_68_113), .C1 (n_71_114), .C2 (n_73_111) );
AOI211_X1 g_56_119 (.ZN (n_56_119), .A (n_60_117), .B (n_66_114), .C1 (n_69_115), .C2 (n_71_112) );
AOI211_X1 g_54_120 (.ZN (n_54_120), .A (n_58_118), .B (n_64_115), .C1 (n_68_113), .C2 (n_73_113) );
AOI211_X1 g_52_121 (.ZN (n_52_121), .A (n_56_119), .B (n_62_116), .C1 (n_66_114), .C2 (n_71_114) );
AOI211_X1 g_50_122 (.ZN (n_50_122), .A (n_54_120), .B (n_60_117), .C1 (n_64_115), .C2 (n_69_115) );
AOI211_X1 g_48_123 (.ZN (n_48_123), .A (n_52_121), .B (n_58_118), .C1 (n_62_116), .C2 (n_68_113) );
AOI211_X1 g_46_124 (.ZN (n_46_124), .A (n_50_122), .B (n_56_119), .C1 (n_60_117), .C2 (n_66_114) );
AOI211_X1 g_44_125 (.ZN (n_44_125), .A (n_48_123), .B (n_54_120), .C1 (n_58_118), .C2 (n_64_115) );
AOI211_X1 g_42_126 (.ZN (n_42_126), .A (n_46_124), .B (n_52_121), .C1 (n_56_119), .C2 (n_62_116) );
AOI211_X1 g_40_127 (.ZN (n_40_127), .A (n_44_125), .B (n_50_122), .C1 (n_54_120), .C2 (n_60_117) );
AOI211_X1 g_38_128 (.ZN (n_38_128), .A (n_42_126), .B (n_48_123), .C1 (n_52_121), .C2 (n_58_118) );
AOI211_X1 g_36_129 (.ZN (n_36_129), .A (n_40_127), .B (n_46_124), .C1 (n_50_122), .C2 (n_56_119) );
AOI211_X1 g_34_130 (.ZN (n_34_130), .A (n_38_128), .B (n_44_125), .C1 (n_48_123), .C2 (n_54_120) );
AOI211_X1 g_32_131 (.ZN (n_32_131), .A (n_36_129), .B (n_42_126), .C1 (n_46_124), .C2 (n_52_121) );
AOI211_X1 g_30_132 (.ZN (n_30_132), .A (n_34_130), .B (n_40_127), .C1 (n_44_125), .C2 (n_50_122) );
AOI211_X1 g_28_133 (.ZN (n_28_133), .A (n_32_131), .B (n_38_128), .C1 (n_42_126), .C2 (n_48_123) );
AOI211_X1 g_27_131 (.ZN (n_27_131), .A (n_30_132), .B (n_36_129), .C1 (n_40_127), .C2 (n_46_124) );
AOI211_X1 g_25_132 (.ZN (n_25_132), .A (n_28_133), .B (n_34_130), .C1 (n_38_128), .C2 (n_44_125) );
AOI211_X1 g_23_133 (.ZN (n_23_133), .A (n_27_131), .B (n_32_131), .C1 (n_36_129), .C2 (n_42_126) );
AOI211_X1 g_21_134 (.ZN (n_21_134), .A (n_25_132), .B (n_30_132), .C1 (n_34_130), .C2 (n_40_127) );
AOI211_X1 g_19_135 (.ZN (n_19_135), .A (n_23_133), .B (n_28_133), .C1 (n_32_131), .C2 (n_38_128) );
AOI211_X1 g_17_136 (.ZN (n_17_136), .A (n_21_134), .B (n_27_131), .C1 (n_30_132), .C2 (n_36_129) );
AOI211_X1 g_15_137 (.ZN (n_15_137), .A (n_19_135), .B (n_25_132), .C1 (n_28_133), .C2 (n_34_130) );
AOI211_X1 g_13_138 (.ZN (n_13_138), .A (n_17_136), .B (n_23_133), .C1 (n_27_131), .C2 (n_32_131) );
AOI211_X1 g_11_139 (.ZN (n_11_139), .A (n_15_137), .B (n_21_134), .C1 (n_25_132), .C2 (n_30_132) );
AOI211_X1 g_9_140 (.ZN (n_9_140), .A (n_13_138), .B (n_19_135), .C1 (n_23_133), .C2 (n_28_133) );
AOI211_X1 g_8_142 (.ZN (n_8_142), .A (n_11_139), .B (n_17_136), .C1 (n_21_134), .C2 (n_27_131) );
AOI211_X1 g_10_141 (.ZN (n_10_141), .A (n_9_140), .B (n_15_137), .C1 (n_19_135), .C2 (n_25_132) );
AOI211_X1 g_12_140 (.ZN (n_12_140), .A (n_8_142), .B (n_13_138), .C1 (n_17_136), .C2 (n_23_133) );
AOI211_X1 g_14_139 (.ZN (n_14_139), .A (n_10_141), .B (n_11_139), .C1 (n_15_137), .C2 (n_21_134) );
AOI211_X1 g_16_138 (.ZN (n_16_138), .A (n_12_140), .B (n_9_140), .C1 (n_13_138), .C2 (n_19_135) );
AOI211_X1 g_18_137 (.ZN (n_18_137), .A (n_14_139), .B (n_8_142), .C1 (n_11_139), .C2 (n_17_136) );
AOI211_X1 g_20_136 (.ZN (n_20_136), .A (n_16_138), .B (n_10_141), .C1 (n_9_140), .C2 (n_15_137) );
AOI211_X1 g_22_135 (.ZN (n_22_135), .A (n_18_137), .B (n_12_140), .C1 (n_8_142), .C2 (n_13_138) );
AOI211_X1 g_24_134 (.ZN (n_24_134), .A (n_20_136), .B (n_14_139), .C1 (n_10_141), .C2 (n_11_139) );
AOI211_X1 g_26_133 (.ZN (n_26_133), .A (n_22_135), .B (n_16_138), .C1 (n_12_140), .C2 (n_9_140) );
AOI211_X1 g_28_132 (.ZN (n_28_132), .A (n_24_134), .B (n_18_137), .C1 (n_14_139), .C2 (n_8_142) );
AOI211_X1 g_27_134 (.ZN (n_27_134), .A (n_26_133), .B (n_20_136), .C1 (n_16_138), .C2 (n_10_141) );
AOI211_X1 g_29_133 (.ZN (n_29_133), .A (n_28_132), .B (n_22_135), .C1 (n_18_137), .C2 (n_12_140) );
AOI211_X1 g_31_132 (.ZN (n_31_132), .A (n_27_134), .B (n_24_134), .C1 (n_20_136), .C2 (n_14_139) );
AOI211_X1 g_33_131 (.ZN (n_33_131), .A (n_29_133), .B (n_26_133), .C1 (n_22_135), .C2 (n_16_138) );
AOI211_X1 g_35_130 (.ZN (n_35_130), .A (n_31_132), .B (n_28_132), .C1 (n_24_134), .C2 (n_18_137) );
AOI211_X1 g_37_129 (.ZN (n_37_129), .A (n_33_131), .B (n_27_134), .C1 (n_26_133), .C2 (n_20_136) );
AOI211_X1 g_39_128 (.ZN (n_39_128), .A (n_35_130), .B (n_29_133), .C1 (n_28_132), .C2 (n_22_135) );
AOI211_X1 g_41_127 (.ZN (n_41_127), .A (n_37_129), .B (n_31_132), .C1 (n_27_134), .C2 (n_24_134) );
AOI211_X1 g_43_126 (.ZN (n_43_126), .A (n_39_128), .B (n_33_131), .C1 (n_29_133), .C2 (n_26_133) );
AOI211_X1 g_45_125 (.ZN (n_45_125), .A (n_41_127), .B (n_35_130), .C1 (n_31_132), .C2 (n_28_132) );
AOI211_X1 g_47_124 (.ZN (n_47_124), .A (n_43_126), .B (n_37_129), .C1 (n_33_131), .C2 (n_27_134) );
AOI211_X1 g_49_123 (.ZN (n_49_123), .A (n_45_125), .B (n_39_128), .C1 (n_35_130), .C2 (n_29_133) );
AOI211_X1 g_51_122 (.ZN (n_51_122), .A (n_47_124), .B (n_41_127), .C1 (n_37_129), .C2 (n_31_132) );
AOI211_X1 g_50_124 (.ZN (n_50_124), .A (n_49_123), .B (n_43_126), .C1 (n_39_128), .C2 (n_33_131) );
AOI211_X1 g_49_122 (.ZN (n_49_122), .A (n_51_122), .B (n_45_125), .C1 (n_41_127), .C2 (n_35_130) );
AOI211_X1 g_51_121 (.ZN (n_51_121), .A (n_50_124), .B (n_47_124), .C1 (n_43_126), .C2 (n_37_129) );
AOI211_X1 g_53_120 (.ZN (n_53_120), .A (n_49_122), .B (n_49_123), .C1 (n_45_125), .C2 (n_39_128) );
AOI211_X1 g_55_119 (.ZN (n_55_119), .A (n_51_121), .B (n_51_122), .C1 (n_47_124), .C2 (n_41_127) );
AOI211_X1 g_57_118 (.ZN (n_57_118), .A (n_53_120), .B (n_50_124), .C1 (n_49_123), .C2 (n_43_126) );
AOI211_X1 g_59_117 (.ZN (n_59_117), .A (n_55_119), .B (n_49_122), .C1 (n_51_122), .C2 (n_45_125) );
AOI211_X1 g_58_119 (.ZN (n_58_119), .A (n_57_118), .B (n_51_121), .C1 (n_50_124), .C2 (n_47_124) );
AOI211_X1 g_60_118 (.ZN (n_60_118), .A (n_59_117), .B (n_53_120), .C1 (n_49_122), .C2 (n_49_123) );
AOI211_X1 g_59_120 (.ZN (n_59_120), .A (n_58_119), .B (n_55_119), .C1 (n_51_121), .C2 (n_51_122) );
AOI211_X1 g_61_119 (.ZN (n_61_119), .A (n_60_118), .B (n_57_118), .C1 (n_53_120), .C2 (n_50_124) );
AOI211_X1 g_63_118 (.ZN (n_63_118), .A (n_59_120), .B (n_59_117), .C1 (n_55_119), .C2 (n_49_122) );
AOI211_X1 g_65_117 (.ZN (n_65_117), .A (n_61_119), .B (n_58_119), .C1 (n_57_118), .C2 (n_51_121) );
AOI211_X1 g_67_116 (.ZN (n_67_116), .A (n_63_118), .B (n_60_118), .C1 (n_59_117), .C2 (n_53_120) );
AOI211_X1 g_66_118 (.ZN (n_66_118), .A (n_65_117), .B (n_59_120), .C1 (n_58_119), .C2 (n_55_119) );
AOI211_X1 g_65_116 (.ZN (n_65_116), .A (n_67_116), .B (n_61_119), .C1 (n_60_118), .C2 (n_57_118) );
AOI211_X1 g_67_115 (.ZN (n_67_115), .A (n_66_118), .B (n_63_118), .C1 (n_59_120), .C2 (n_59_117) );
AOI211_X1 g_69_114 (.ZN (n_69_114), .A (n_65_116), .B (n_65_117), .C1 (n_61_119), .C2 (n_58_119) );
AOI211_X1 g_71_113 (.ZN (n_71_113), .A (n_67_115), .B (n_67_116), .C1 (n_63_118), .C2 (n_60_118) );
AOI211_X1 g_73_112 (.ZN (n_73_112), .A (n_69_114), .B (n_66_118), .C1 (n_65_117), .C2 (n_59_120) );
AOI211_X1 g_75_111 (.ZN (n_75_111), .A (n_71_113), .B (n_65_116), .C1 (n_67_116), .C2 (n_61_119) );
AOI211_X1 g_77_110 (.ZN (n_77_110), .A (n_73_112), .B (n_67_115), .C1 (n_66_118), .C2 (n_63_118) );
AOI211_X1 g_79_109 (.ZN (n_79_109), .A (n_75_111), .B (n_69_114), .C1 (n_65_116), .C2 (n_65_117) );
AOI211_X1 g_81_108 (.ZN (n_81_108), .A (n_77_110), .B (n_71_113), .C1 (n_67_115), .C2 (n_67_116) );
AOI211_X1 g_82_106 (.ZN (n_82_106), .A (n_79_109), .B (n_73_112), .C1 (n_69_114), .C2 (n_66_118) );
AOI211_X1 g_84_105 (.ZN (n_84_105), .A (n_81_108), .B (n_75_111), .C1 (n_71_113), .C2 (n_65_116) );
AOI211_X1 g_86_104 (.ZN (n_86_104), .A (n_82_106), .B (n_77_110), .C1 (n_73_112), .C2 (n_67_115) );
AOI211_X1 g_88_103 (.ZN (n_88_103), .A (n_84_105), .B (n_79_109), .C1 (n_75_111), .C2 (n_69_114) );
AOI211_X1 g_90_102 (.ZN (n_90_102), .A (n_86_104), .B (n_81_108), .C1 (n_77_110), .C2 (n_71_113) );
AOI211_X1 g_92_101 (.ZN (n_92_101), .A (n_88_103), .B (n_82_106), .C1 (n_79_109), .C2 (n_73_112) );
AOI211_X1 g_94_100 (.ZN (n_94_100), .A (n_90_102), .B (n_84_105), .C1 (n_81_108), .C2 (n_75_111) );
AOI211_X1 g_96_99 (.ZN (n_96_99), .A (n_92_101), .B (n_86_104), .C1 (n_82_106), .C2 (n_77_110) );
AOI211_X1 g_95_101 (.ZN (n_95_101), .A (n_94_100), .B (n_88_103), .C1 (n_84_105), .C2 (n_79_109) );
AOI211_X1 g_97_100 (.ZN (n_97_100), .A (n_96_99), .B (n_90_102), .C1 (n_86_104), .C2 (n_81_108) );
AOI211_X1 g_96_102 (.ZN (n_96_102), .A (n_95_101), .B (n_92_101), .C1 (n_88_103), .C2 (n_82_106) );
AOI211_X1 g_95_100 (.ZN (n_95_100), .A (n_97_100), .B (n_94_100), .C1 (n_90_102), .C2 (n_84_105) );
AOI211_X1 g_93_101 (.ZN (n_93_101), .A (n_96_102), .B (n_96_99), .C1 (n_92_101), .C2 (n_86_104) );
AOI211_X1 g_91_102 (.ZN (n_91_102), .A (n_95_100), .B (n_95_101), .C1 (n_94_100), .C2 (n_88_103) );
AOI211_X1 g_89_103 (.ZN (n_89_103), .A (n_93_101), .B (n_97_100), .C1 (n_96_99), .C2 (n_90_102) );
AOI211_X1 g_87_104 (.ZN (n_87_104), .A (n_91_102), .B (n_96_102), .C1 (n_95_101), .C2 (n_92_101) );
AOI211_X1 g_85_105 (.ZN (n_85_105), .A (n_89_103), .B (n_95_100), .C1 (n_97_100), .C2 (n_94_100) );
AOI211_X1 g_83_106 (.ZN (n_83_106), .A (n_87_104), .B (n_93_101), .C1 (n_96_102), .C2 (n_96_99) );
AOI211_X1 g_81_107 (.ZN (n_81_107), .A (n_85_105), .B (n_91_102), .C1 (n_95_100), .C2 (n_95_101) );
AOI211_X1 g_79_108 (.ZN (n_79_108), .A (n_83_106), .B (n_89_103), .C1 (n_93_101), .C2 (n_97_100) );
AOI211_X1 g_77_109 (.ZN (n_77_109), .A (n_81_107), .B (n_87_104), .C1 (n_91_102), .C2 (n_96_102) );
AOI211_X1 g_75_110 (.ZN (n_75_110), .A (n_79_108), .B (n_85_105), .C1 (n_89_103), .C2 (n_95_100) );
AOI211_X1 g_77_111 (.ZN (n_77_111), .A (n_77_109), .B (n_83_106), .C1 (n_87_104), .C2 (n_93_101) );
AOI211_X1 g_79_110 (.ZN (n_79_110), .A (n_75_110), .B (n_81_107), .C1 (n_85_105), .C2 (n_91_102) );
AOI211_X1 g_81_109 (.ZN (n_81_109), .A (n_77_111), .B (n_79_108), .C1 (n_83_106), .C2 (n_89_103) );
AOI211_X1 g_83_108 (.ZN (n_83_108), .A (n_79_110), .B (n_77_109), .C1 (n_81_107), .C2 (n_87_104) );
AOI211_X1 g_85_107 (.ZN (n_85_107), .A (n_81_109), .B (n_75_110), .C1 (n_79_108), .C2 (n_85_105) );
AOI211_X1 g_87_106 (.ZN (n_87_106), .A (n_83_108), .B (n_77_111), .C1 (n_77_109), .C2 (n_83_106) );
AOI211_X1 g_89_105 (.ZN (n_89_105), .A (n_85_107), .B (n_79_110), .C1 (n_75_110), .C2 (n_81_107) );
AOI211_X1 g_91_104 (.ZN (n_91_104), .A (n_87_106), .B (n_81_109), .C1 (n_77_111), .C2 (n_79_108) );
AOI211_X1 g_93_103 (.ZN (n_93_103), .A (n_89_105), .B (n_83_108), .C1 (n_79_110), .C2 (n_77_109) );
AOI211_X1 g_95_102 (.ZN (n_95_102), .A (n_91_104), .B (n_85_107), .C1 (n_81_109), .C2 (n_75_110) );
AOI211_X1 g_97_101 (.ZN (n_97_101), .A (n_93_103), .B (n_87_106), .C1 (n_83_108), .C2 (n_77_111) );
AOI211_X1 g_96_103 (.ZN (n_96_103), .A (n_95_102), .B (n_89_105), .C1 (n_85_107), .C2 (n_79_110) );
AOI211_X1 g_94_102 (.ZN (n_94_102), .A (n_97_101), .B (n_91_104), .C1 (n_87_106), .C2 (n_81_109) );
AOI211_X1 g_96_101 (.ZN (n_96_101), .A (n_96_103), .B (n_93_103), .C1 (n_89_105), .C2 (n_83_108) );
AOI211_X1 g_98_100 (.ZN (n_98_100), .A (n_94_102), .B (n_95_102), .C1 (n_91_104), .C2 (n_85_107) );
AOI211_X1 g_100_99 (.ZN (n_100_99), .A (n_96_101), .B (n_97_101), .C1 (n_93_103), .C2 (n_87_106) );
AOI211_X1 g_102_98 (.ZN (n_102_98), .A (n_98_100), .B (n_96_103), .C1 (n_95_102), .C2 (n_89_105) );
AOI211_X1 g_104_97 (.ZN (n_104_97), .A (n_100_99), .B (n_94_102), .C1 (n_97_101), .C2 (n_91_104) );
AOI211_X1 g_106_98 (.ZN (n_106_98), .A (n_102_98), .B (n_96_101), .C1 (n_96_103), .C2 (n_93_103) );
AOI211_X1 g_105_100 (.ZN (n_105_100), .A (n_104_97), .B (n_98_100), .C1 (n_94_102), .C2 (n_95_102) );
AOI211_X1 g_103_99 (.ZN (n_103_99), .A (n_106_98), .B (n_100_99), .C1 (n_96_101), .C2 (n_97_101) );
AOI211_X1 g_105_98 (.ZN (n_105_98), .A (n_105_100), .B (n_102_98), .C1 (n_98_100), .C2 (n_96_103) );
AOI211_X1 g_107_97 (.ZN (n_107_97), .A (n_103_99), .B (n_104_97), .C1 (n_100_99), .C2 (n_94_102) );
AOI211_X1 g_109_96 (.ZN (n_109_96), .A (n_105_98), .B (n_106_98), .C1 (n_102_98), .C2 (n_96_101) );
AOI211_X1 g_111_95 (.ZN (n_111_95), .A (n_107_97), .B (n_105_100), .C1 (n_104_97), .C2 (n_98_100) );
AOI211_X1 g_113_94 (.ZN (n_113_94), .A (n_109_96), .B (n_103_99), .C1 (n_106_98), .C2 (n_100_99) );
AOI211_X1 g_115_93 (.ZN (n_115_93), .A (n_111_95), .B (n_105_98), .C1 (n_105_100), .C2 (n_102_98) );
AOI211_X1 g_117_92 (.ZN (n_117_92), .A (n_113_94), .B (n_107_97), .C1 (n_103_99), .C2 (n_104_97) );
AOI211_X1 g_119_91 (.ZN (n_119_91), .A (n_115_93), .B (n_109_96), .C1 (n_105_98), .C2 (n_106_98) );
AOI211_X1 g_121_90 (.ZN (n_121_90), .A (n_117_92), .B (n_111_95), .C1 (n_107_97), .C2 (n_105_100) );
AOI211_X1 g_120_92 (.ZN (n_120_92), .A (n_119_91), .B (n_113_94), .C1 (n_109_96), .C2 (n_103_99) );
AOI211_X1 g_118_93 (.ZN (n_118_93), .A (n_121_90), .B (n_115_93), .C1 (n_111_95), .C2 (n_105_98) );
AOI211_X1 g_116_94 (.ZN (n_116_94), .A (n_120_92), .B (n_117_92), .C1 (n_113_94), .C2 (n_107_97) );
AOI211_X1 g_114_95 (.ZN (n_114_95), .A (n_118_93), .B (n_119_91), .C1 (n_115_93), .C2 (n_109_96) );
AOI211_X1 g_112_96 (.ZN (n_112_96), .A (n_116_94), .B (n_121_90), .C1 (n_117_92), .C2 (n_111_95) );
AOI211_X1 g_110_97 (.ZN (n_110_97), .A (n_114_95), .B (n_120_92), .C1 (n_119_91), .C2 (n_113_94) );
AOI211_X1 g_108_98 (.ZN (n_108_98), .A (n_112_96), .B (n_118_93), .C1 (n_121_90), .C2 (n_115_93) );
AOI211_X1 g_106_99 (.ZN (n_106_99), .A (n_110_97), .B (n_116_94), .C1 (n_120_92), .C2 (n_117_92) );
AOI211_X1 g_104_100 (.ZN (n_104_100), .A (n_108_98), .B (n_114_95), .C1 (n_118_93), .C2 (n_119_91) );
AOI211_X1 g_102_101 (.ZN (n_102_101), .A (n_106_99), .B (n_112_96), .C1 (n_116_94), .C2 (n_121_90) );
AOI211_X1 g_100_102 (.ZN (n_100_102), .A (n_104_100), .B (n_110_97), .C1 (n_114_95), .C2 (n_120_92) );
AOI211_X1 g_101_100 (.ZN (n_101_100), .A (n_102_101), .B (n_108_98), .C1 (n_112_96), .C2 (n_118_93) );
AOI211_X1 g_99_101 (.ZN (n_99_101), .A (n_100_102), .B (n_106_99), .C1 (n_110_97), .C2 (n_116_94) );
AOI211_X1 g_97_102 (.ZN (n_97_102), .A (n_101_100), .B (n_104_100), .C1 (n_108_98), .C2 (n_114_95) );
AOI211_X1 g_95_103 (.ZN (n_95_103), .A (n_99_101), .B (n_102_101), .C1 (n_106_99), .C2 (n_112_96) );
AOI211_X1 g_93_102 (.ZN (n_93_102), .A (n_97_102), .B (n_100_102), .C1 (n_104_100), .C2 (n_110_97) );
AOI211_X1 g_91_103 (.ZN (n_91_103), .A (n_95_103), .B (n_101_100), .C1 (n_102_101), .C2 (n_108_98) );
AOI211_X1 g_89_104 (.ZN (n_89_104), .A (n_93_102), .B (n_99_101), .C1 (n_100_102), .C2 (n_106_99) );
AOI211_X1 g_87_105 (.ZN (n_87_105), .A (n_91_103), .B (n_97_102), .C1 (n_101_100), .C2 (n_104_100) );
AOI211_X1 g_85_106 (.ZN (n_85_106), .A (n_89_104), .B (n_95_103), .C1 (n_99_101), .C2 (n_102_101) );
AOI211_X1 g_83_107 (.ZN (n_83_107), .A (n_87_105), .B (n_93_102), .C1 (n_97_102), .C2 (n_100_102) );
AOI211_X1 g_82_109 (.ZN (n_82_109), .A (n_85_106), .B (n_91_103), .C1 (n_95_103), .C2 (n_101_100) );
AOI211_X1 g_84_108 (.ZN (n_84_108), .A (n_83_107), .B (n_89_104), .C1 (n_93_102), .C2 (n_99_101) );
AOI211_X1 g_86_107 (.ZN (n_86_107), .A (n_82_109), .B (n_87_105), .C1 (n_91_103), .C2 (n_97_102) );
AOI211_X1 g_88_106 (.ZN (n_88_106), .A (n_84_108), .B (n_85_106), .C1 (n_89_104), .C2 (n_95_103) );
AOI211_X1 g_90_105 (.ZN (n_90_105), .A (n_86_107), .B (n_83_107), .C1 (n_87_105), .C2 (n_93_102) );
AOI211_X1 g_92_104 (.ZN (n_92_104), .A (n_88_106), .B (n_82_109), .C1 (n_85_106), .C2 (n_91_103) );
AOI211_X1 g_94_103 (.ZN (n_94_103), .A (n_90_105), .B (n_84_108), .C1 (n_83_107), .C2 (n_89_104) );
AOI211_X1 g_96_104 (.ZN (n_96_104), .A (n_92_104), .B (n_86_107), .C1 (n_82_109), .C2 (n_87_105) );
AOI211_X1 g_98_103 (.ZN (n_98_103), .A (n_94_103), .B (n_88_106), .C1 (n_84_108), .C2 (n_85_106) );
AOI211_X1 g_97_105 (.ZN (n_97_105), .A (n_96_104), .B (n_90_105), .C1 (n_86_107), .C2 (n_83_107) );
AOI211_X1 g_95_104 (.ZN (n_95_104), .A (n_98_103), .B (n_92_104), .C1 (n_88_106), .C2 (n_82_109) );
AOI211_X1 g_97_103 (.ZN (n_97_103), .A (n_97_105), .B (n_94_103), .C1 (n_90_105), .C2 (n_84_108) );
AOI211_X1 g_99_102 (.ZN (n_99_102), .A (n_95_104), .B (n_96_104), .C1 (n_92_104), .C2 (n_86_107) );
AOI211_X1 g_101_101 (.ZN (n_101_101), .A (n_97_103), .B (n_98_103), .C1 (n_94_103), .C2 (n_88_106) );
AOI211_X1 g_103_100 (.ZN (n_103_100), .A (n_99_102), .B (n_97_105), .C1 (n_96_104), .C2 (n_90_105) );
AOI211_X1 g_104_102 (.ZN (n_104_102), .A (n_101_101), .B (n_95_104), .C1 (n_98_103), .C2 (n_92_104) );
AOI211_X1 g_106_101 (.ZN (n_106_101), .A (n_103_100), .B (n_97_103), .C1 (n_97_105), .C2 (n_94_103) );
AOI211_X1 g_107_99 (.ZN (n_107_99), .A (n_104_102), .B (n_99_102), .C1 (n_95_104), .C2 (n_96_104) );
AOI211_X1 g_109_98 (.ZN (n_109_98), .A (n_106_101), .B (n_101_101), .C1 (n_97_103), .C2 (n_98_103) );
AOI211_X1 g_110_96 (.ZN (n_110_96), .A (n_107_99), .B (n_103_100), .C1 (n_99_102), .C2 (n_97_105) );
AOI211_X1 g_112_95 (.ZN (n_112_95), .A (n_109_98), .B (n_104_102), .C1 (n_101_101), .C2 (n_95_104) );
AOI211_X1 g_114_94 (.ZN (n_114_94), .A (n_110_96), .B (n_106_101), .C1 (n_103_100), .C2 (n_97_103) );
AOI211_X1 g_116_93 (.ZN (n_116_93), .A (n_112_95), .B (n_107_99), .C1 (n_104_102), .C2 (n_99_102) );
AOI211_X1 g_118_92 (.ZN (n_118_92), .A (n_114_94), .B (n_109_98), .C1 (n_106_101), .C2 (n_101_101) );
AOI211_X1 g_120_91 (.ZN (n_120_91), .A (n_116_93), .B (n_110_96), .C1 (n_107_99), .C2 (n_103_100) );
AOI211_X1 g_122_90 (.ZN (n_122_90), .A (n_118_92), .B (n_112_95), .C1 (n_109_98), .C2 (n_104_102) );
AOI211_X1 g_124_91 (.ZN (n_124_91), .A (n_120_91), .B (n_114_94), .C1 (n_110_96), .C2 (n_106_101) );
AOI211_X1 g_122_92 (.ZN (n_122_92), .A (n_122_90), .B (n_116_93), .C1 (n_112_95), .C2 (n_107_99) );
AOI211_X1 g_123_90 (.ZN (n_123_90), .A (n_124_91), .B (n_118_92), .C1 (n_114_94), .C2 (n_109_98) );
AOI211_X1 g_121_91 (.ZN (n_121_91), .A (n_122_92), .B (n_120_91), .C1 (n_116_93), .C2 (n_110_96) );
AOI211_X1 g_120_93 (.ZN (n_120_93), .A (n_123_90), .B (n_122_90), .C1 (n_118_92), .C2 (n_112_95) );
AOI211_X1 g_118_94 (.ZN (n_118_94), .A (n_121_91), .B (n_124_91), .C1 (n_120_91), .C2 (n_114_94) );
AOI211_X1 g_116_95 (.ZN (n_116_95), .A (n_120_93), .B (n_122_92), .C1 (n_122_90), .C2 (n_116_93) );
AOI211_X1 g_114_96 (.ZN (n_114_96), .A (n_118_94), .B (n_123_90), .C1 (n_124_91), .C2 (n_118_92) );
AOI211_X1 g_112_97 (.ZN (n_112_97), .A (n_116_95), .B (n_121_91), .C1 (n_122_92), .C2 (n_120_91) );
AOI211_X1 g_110_98 (.ZN (n_110_98), .A (n_114_96), .B (n_120_93), .C1 (n_123_90), .C2 (n_122_90) );
AOI211_X1 g_108_99 (.ZN (n_108_99), .A (n_112_97), .B (n_118_94), .C1 (n_121_91), .C2 (n_124_91) );
AOI211_X1 g_106_100 (.ZN (n_106_100), .A (n_110_98), .B (n_116_95), .C1 (n_120_93), .C2 (n_122_92) );
AOI211_X1 g_104_101 (.ZN (n_104_101), .A (n_108_99), .B (n_114_96), .C1 (n_118_94), .C2 (n_123_90) );
AOI211_X1 g_102_100 (.ZN (n_102_100), .A (n_106_100), .B (n_112_97), .C1 (n_116_95), .C2 (n_121_91) );
AOI211_X1 g_100_101 (.ZN (n_100_101), .A (n_104_101), .B (n_110_98), .C1 (n_114_96), .C2 (n_120_93) );
AOI211_X1 g_98_102 (.ZN (n_98_102), .A (n_102_100), .B (n_108_99), .C1 (n_112_97), .C2 (n_118_94) );
AOI211_X1 g_99_104 (.ZN (n_99_104), .A (n_100_101), .B (n_106_100), .C1 (n_110_98), .C2 (n_116_95) );
AOI211_X1 g_101_103 (.ZN (n_101_103), .A (n_98_102), .B (n_104_101), .C1 (n_108_99), .C2 (n_114_96) );
AOI211_X1 g_103_102 (.ZN (n_103_102), .A (n_99_104), .B (n_102_100), .C1 (n_106_100), .C2 (n_112_97) );
AOI211_X1 g_105_101 (.ZN (n_105_101), .A (n_101_103), .B (n_100_101), .C1 (n_104_101), .C2 (n_110_98) );
AOI211_X1 g_107_100 (.ZN (n_107_100), .A (n_103_102), .B (n_98_102), .C1 (n_102_100), .C2 (n_108_99) );
AOI211_X1 g_109_99 (.ZN (n_109_99), .A (n_105_101), .B (n_99_104), .C1 (n_100_101), .C2 (n_106_100) );
AOI211_X1 g_111_98 (.ZN (n_111_98), .A (n_107_100), .B (n_101_103), .C1 (n_98_102), .C2 (n_104_101) );
AOI211_X1 g_113_97 (.ZN (n_113_97), .A (n_109_99), .B (n_103_102), .C1 (n_99_104), .C2 (n_102_100) );
AOI211_X1 g_115_96 (.ZN (n_115_96), .A (n_111_98), .B (n_105_101), .C1 (n_101_103), .C2 (n_100_101) );
AOI211_X1 g_117_95 (.ZN (n_117_95), .A (n_113_97), .B (n_107_100), .C1 (n_103_102), .C2 (n_98_102) );
AOI211_X1 g_119_94 (.ZN (n_119_94), .A (n_115_96), .B (n_109_99), .C1 (n_105_101), .C2 (n_99_104) );
AOI211_X1 g_121_93 (.ZN (n_121_93), .A (n_117_95), .B (n_111_98), .C1 (n_107_100), .C2 (n_101_103) );
AOI211_X1 g_123_92 (.ZN (n_123_92), .A (n_119_94), .B (n_113_97), .C1 (n_109_99), .C2 (n_103_102) );
AOI211_X1 g_125_91 (.ZN (n_125_91), .A (n_121_93), .B (n_115_96), .C1 (n_111_98), .C2 (n_105_101) );
AOI211_X1 g_124_93 (.ZN (n_124_93), .A (n_123_92), .B (n_117_95), .C1 (n_113_97), .C2 (n_107_100) );
AOI211_X1 g_123_91 (.ZN (n_123_91), .A (n_125_91), .B (n_119_94), .C1 (n_115_96), .C2 (n_109_99) );
AOI211_X1 g_125_90 (.ZN (n_125_90), .A (n_124_93), .B (n_121_93), .C1 (n_117_95), .C2 (n_111_98) );
AOI211_X1 g_127_89 (.ZN (n_127_89), .A (n_123_91), .B (n_123_92), .C1 (n_119_94), .C2 (n_113_97) );
AOI211_X1 g_129_88 (.ZN (n_129_88), .A (n_125_90), .B (n_125_91), .C1 (n_121_93), .C2 (n_115_96) );
AOI211_X1 g_131_87 (.ZN (n_131_87), .A (n_127_89), .B (n_124_93), .C1 (n_123_92), .C2 (n_117_95) );
AOI211_X1 g_133_86 (.ZN (n_133_86), .A (n_129_88), .B (n_123_91), .C1 (n_125_91), .C2 (n_119_94) );
AOI211_X1 g_135_85 (.ZN (n_135_85), .A (n_131_87), .B (n_125_90), .C1 (n_124_93), .C2 (n_121_93) );
AOI211_X1 g_137_84 (.ZN (n_137_84), .A (n_133_86), .B (n_127_89), .C1 (n_123_91), .C2 (n_123_92) );
AOI211_X1 g_139_83 (.ZN (n_139_83), .A (n_135_85), .B (n_129_88), .C1 (n_125_90), .C2 (n_125_91) );
AOI211_X1 g_138_85 (.ZN (n_138_85), .A (n_137_84), .B (n_131_87), .C1 (n_127_89), .C2 (n_124_93) );
AOI211_X1 g_136_86 (.ZN (n_136_86), .A (n_139_83), .B (n_133_86), .C1 (n_129_88), .C2 (n_123_91) );
AOI211_X1 g_134_87 (.ZN (n_134_87), .A (n_138_85), .B (n_135_85), .C1 (n_131_87), .C2 (n_125_90) );
AOI211_X1 g_132_88 (.ZN (n_132_88), .A (n_136_86), .B (n_137_84), .C1 (n_133_86), .C2 (n_127_89) );
AOI211_X1 g_130_89 (.ZN (n_130_89), .A (n_134_87), .B (n_139_83), .C1 (n_135_85), .C2 (n_129_88) );
AOI211_X1 g_128_90 (.ZN (n_128_90), .A (n_132_88), .B (n_138_85), .C1 (n_137_84), .C2 (n_131_87) );
AOI211_X1 g_126_91 (.ZN (n_126_91), .A (n_130_89), .B (n_136_86), .C1 (n_139_83), .C2 (n_133_86) );
AOI211_X1 g_124_92 (.ZN (n_124_92), .A (n_128_90), .B (n_134_87), .C1 (n_138_85), .C2 (n_135_85) );
AOI211_X1 g_122_93 (.ZN (n_122_93), .A (n_126_91), .B (n_132_88), .C1 (n_136_86), .C2 (n_137_84) );
AOI211_X1 g_120_94 (.ZN (n_120_94), .A (n_124_92), .B (n_130_89), .C1 (n_134_87), .C2 (n_139_83) );
AOI211_X1 g_121_92 (.ZN (n_121_92), .A (n_122_93), .B (n_128_90), .C1 (n_132_88), .C2 (n_138_85) );
AOI211_X1 g_119_93 (.ZN (n_119_93), .A (n_120_94), .B (n_126_91), .C1 (n_130_89), .C2 (n_136_86) );
AOI211_X1 g_117_94 (.ZN (n_117_94), .A (n_121_92), .B (n_124_92), .C1 (n_128_90), .C2 (n_134_87) );
AOI211_X1 g_115_95 (.ZN (n_115_95), .A (n_119_93), .B (n_122_93), .C1 (n_126_91), .C2 (n_132_88) );
AOI211_X1 g_113_96 (.ZN (n_113_96), .A (n_117_94), .B (n_120_94), .C1 (n_124_92), .C2 (n_130_89) );
AOI211_X1 g_111_97 (.ZN (n_111_97), .A (n_115_95), .B (n_121_92), .C1 (n_122_93), .C2 (n_128_90) );
AOI211_X1 g_110_99 (.ZN (n_110_99), .A (n_113_96), .B (n_119_93), .C1 (n_120_94), .C2 (n_126_91) );
AOI211_X1 g_108_100 (.ZN (n_108_100), .A (n_111_97), .B (n_117_94), .C1 (n_121_92), .C2 (n_124_92) );
AOI211_X1 g_107_102 (.ZN (n_107_102), .A (n_110_99), .B (n_115_95), .C1 (n_119_93), .C2 (n_122_93) );
AOI211_X1 g_109_101 (.ZN (n_109_101), .A (n_108_100), .B (n_113_96), .C1 (n_117_94), .C2 (n_120_94) );
AOI211_X1 g_111_100 (.ZN (n_111_100), .A (n_107_102), .B (n_111_97), .C1 (n_115_95), .C2 (n_121_92) );
AOI211_X1 g_112_98 (.ZN (n_112_98), .A (n_109_101), .B (n_110_99), .C1 (n_113_96), .C2 (n_119_93) );
AOI211_X1 g_114_97 (.ZN (n_114_97), .A (n_111_100), .B (n_108_100), .C1 (n_111_97), .C2 (n_117_94) );
AOI211_X1 g_116_96 (.ZN (n_116_96), .A (n_112_98), .B (n_107_102), .C1 (n_110_99), .C2 (n_115_95) );
AOI211_X1 g_118_95 (.ZN (n_118_95), .A (n_114_97), .B (n_109_101), .C1 (n_108_100), .C2 (n_113_96) );
AOI211_X1 g_117_97 (.ZN (n_117_97), .A (n_116_96), .B (n_111_100), .C1 (n_107_102), .C2 (n_111_97) );
AOI211_X1 g_119_96 (.ZN (n_119_96), .A (n_118_95), .B (n_112_98), .C1 (n_109_101), .C2 (n_110_99) );
AOI211_X1 g_121_95 (.ZN (n_121_95), .A (n_117_97), .B (n_114_97), .C1 (n_111_100), .C2 (n_108_100) );
AOI211_X1 g_123_94 (.ZN (n_123_94), .A (n_119_96), .B (n_116_96), .C1 (n_112_98), .C2 (n_107_102) );
AOI211_X1 g_125_93 (.ZN (n_125_93), .A (n_121_95), .B (n_118_95), .C1 (n_114_97), .C2 (n_109_101) );
AOI211_X1 g_127_92 (.ZN (n_127_92), .A (n_123_94), .B (n_117_97), .C1 (n_116_96), .C2 (n_111_100) );
AOI211_X1 g_129_91 (.ZN (n_129_91), .A (n_125_93), .B (n_119_96), .C1 (n_118_95), .C2 (n_112_98) );
AOI211_X1 g_128_89 (.ZN (n_128_89), .A (n_127_92), .B (n_121_95), .C1 (n_117_97), .C2 (n_114_97) );
AOI211_X1 g_130_88 (.ZN (n_130_88), .A (n_129_91), .B (n_123_94), .C1 (n_119_96), .C2 (n_116_96) );
AOI211_X1 g_132_87 (.ZN (n_132_87), .A (n_128_89), .B (n_125_93), .C1 (n_121_95), .C2 (n_118_95) );
AOI211_X1 g_134_86 (.ZN (n_134_86), .A (n_130_88), .B (n_127_92), .C1 (n_123_94), .C2 (n_117_97) );
AOI211_X1 g_136_85 (.ZN (n_136_85), .A (n_132_87), .B (n_129_91), .C1 (n_125_93), .C2 (n_119_96) );
AOI211_X1 g_138_84 (.ZN (n_138_84), .A (n_134_86), .B (n_128_89), .C1 (n_127_92), .C2 (n_121_95) );
AOI211_X1 g_139_86 (.ZN (n_139_86), .A (n_136_85), .B (n_130_88), .C1 (n_129_91), .C2 (n_123_94) );
AOI211_X1 g_137_87 (.ZN (n_137_87), .A (n_138_84), .B (n_132_87), .C1 (n_128_89), .C2 (n_125_93) );
AOI211_X1 g_135_88 (.ZN (n_135_88), .A (n_139_86), .B (n_134_86), .C1 (n_130_88), .C2 (n_127_92) );
AOI211_X1 g_133_89 (.ZN (n_133_89), .A (n_137_87), .B (n_136_85), .C1 (n_132_87), .C2 (n_129_91) );
AOI211_X1 g_131_90 (.ZN (n_131_90), .A (n_135_88), .B (n_138_84), .C1 (n_134_86), .C2 (n_128_89) );
AOI211_X1 g_130_92 (.ZN (n_130_92), .A (n_133_89), .B (n_139_86), .C1 (n_136_85), .C2 (n_130_88) );
AOI211_X1 g_129_90 (.ZN (n_129_90), .A (n_131_90), .B (n_137_87), .C1 (n_138_84), .C2 (n_132_87) );
AOI211_X1 g_131_89 (.ZN (n_131_89), .A (n_130_92), .B (n_135_88), .C1 (n_139_86), .C2 (n_134_86) );
AOI211_X1 g_133_88 (.ZN (n_133_88), .A (n_129_90), .B (n_133_89), .C1 (n_137_87), .C2 (n_136_85) );
AOI211_X1 g_135_87 (.ZN (n_135_87), .A (n_131_89), .B (n_131_90), .C1 (n_135_88), .C2 (n_138_84) );
AOI211_X1 g_137_86 (.ZN (n_137_86), .A (n_133_88), .B (n_130_92), .C1 (n_133_89), .C2 (n_139_86) );
AOI211_X1 g_139_85 (.ZN (n_139_85), .A (n_135_87), .B (n_129_90), .C1 (n_131_90), .C2 (n_137_87) );
AOI211_X1 g_141_84 (.ZN (n_141_84), .A (n_137_86), .B (n_131_89), .C1 (n_130_92), .C2 (n_135_88) );
AOI211_X1 g_143_83 (.ZN (n_143_83), .A (n_139_85), .B (n_133_88), .C1 (n_129_90), .C2 (n_133_89) );
AOI211_X1 g_144_85 (.ZN (n_144_85), .A (n_141_84), .B (n_135_87), .C1 (n_131_89), .C2 (n_131_90) );
AOI211_X1 g_146_86 (.ZN (n_146_86), .A (n_143_83), .B (n_137_86), .C1 (n_133_88), .C2 (n_130_92) );
AOI211_X1 g_145_84 (.ZN (n_145_84), .A (n_144_85), .B (n_139_85), .C1 (n_135_87), .C2 (n_129_90) );
AOI211_X1 g_147_85 (.ZN (n_147_85), .A (n_146_86), .B (n_141_84), .C1 (n_137_86), .C2 (n_131_89) );
AOI211_X1 g_148_87 (.ZN (n_148_87), .A (n_145_84), .B (n_143_83), .C1 (n_139_85), .C2 (n_133_88) );
AOI211_X1 g_146_88 (.ZN (n_146_88), .A (n_147_85), .B (n_144_85), .C1 (n_141_84), .C2 (n_135_87) );
AOI211_X1 g_145_86 (.ZN (n_145_86), .A (n_148_87), .B (n_146_86), .C1 (n_143_83), .C2 (n_137_86) );
AOI211_X1 g_143_85 (.ZN (n_143_85), .A (n_146_88), .B (n_145_84), .C1 (n_144_85), .C2 (n_139_85) );
AOI211_X1 g_141_86 (.ZN (n_141_86), .A (n_145_86), .B (n_147_85), .C1 (n_146_86), .C2 (n_141_84) );
AOI211_X1 g_139_87 (.ZN (n_139_87), .A (n_143_85), .B (n_148_87), .C1 (n_145_84), .C2 (n_143_83) );
AOI211_X1 g_140_85 (.ZN (n_140_85), .A (n_141_86), .B (n_146_88), .C1 (n_147_85), .C2 (n_144_85) );
AOI211_X1 g_138_86 (.ZN (n_138_86), .A (n_139_87), .B (n_145_86), .C1 (n_148_87), .C2 (n_146_86) );
AOI211_X1 g_136_87 (.ZN (n_136_87), .A (n_140_85), .B (n_143_85), .C1 (n_146_88), .C2 (n_145_84) );
AOI211_X1 g_134_88 (.ZN (n_134_88), .A (n_138_86), .B (n_141_86), .C1 (n_145_86), .C2 (n_147_85) );
AOI211_X1 g_132_89 (.ZN (n_132_89), .A (n_136_87), .B (n_139_87), .C1 (n_143_85), .C2 (n_148_87) );
AOI211_X1 g_130_90 (.ZN (n_130_90), .A (n_134_88), .B (n_140_85), .C1 (n_141_86), .C2 (n_146_88) );
AOI211_X1 g_128_91 (.ZN (n_128_91), .A (n_132_89), .B (n_138_86), .C1 (n_139_87), .C2 (n_145_86) );
AOI211_X1 g_126_92 (.ZN (n_126_92), .A (n_130_90), .B (n_136_87), .C1 (n_140_85), .C2 (n_143_85) );
AOI211_X1 g_128_93 (.ZN (n_128_93), .A (n_128_91), .B (n_134_88), .C1 (n_138_86), .C2 (n_141_86) );
AOI211_X1 g_127_91 (.ZN (n_127_91), .A (n_126_92), .B (n_132_89), .C1 (n_136_87), .C2 (n_139_87) );
AOI211_X1 g_125_92 (.ZN (n_125_92), .A (n_128_93), .B (n_130_90), .C1 (n_134_88), .C2 (n_140_85) );
AOI211_X1 g_123_93 (.ZN (n_123_93), .A (n_127_91), .B (n_128_91), .C1 (n_132_89), .C2 (n_138_86) );
AOI211_X1 g_121_94 (.ZN (n_121_94), .A (n_125_92), .B (n_126_92), .C1 (n_130_90), .C2 (n_136_87) );
AOI211_X1 g_119_95 (.ZN (n_119_95), .A (n_123_93), .B (n_128_93), .C1 (n_128_91), .C2 (n_134_88) );
AOI211_X1 g_117_96 (.ZN (n_117_96), .A (n_121_94), .B (n_127_91), .C1 (n_126_92), .C2 (n_132_89) );
AOI211_X1 g_115_97 (.ZN (n_115_97), .A (n_119_95), .B (n_125_92), .C1 (n_128_93), .C2 (n_130_90) );
AOI211_X1 g_113_98 (.ZN (n_113_98), .A (n_117_96), .B (n_123_93), .C1 (n_127_91), .C2 (n_128_91) );
AOI211_X1 g_111_99 (.ZN (n_111_99), .A (n_115_97), .B (n_121_94), .C1 (n_125_92), .C2 (n_126_92) );
AOI211_X1 g_109_100 (.ZN (n_109_100), .A (n_113_98), .B (n_119_95), .C1 (n_123_93), .C2 (n_128_93) );
AOI211_X1 g_107_101 (.ZN (n_107_101), .A (n_111_99), .B (n_117_96), .C1 (n_121_94), .C2 (n_127_91) );
AOI211_X1 g_105_102 (.ZN (n_105_102), .A (n_109_100), .B (n_115_97), .C1 (n_119_95), .C2 (n_125_92) );
AOI211_X1 g_103_101 (.ZN (n_103_101), .A (n_107_101), .B (n_113_98), .C1 (n_117_96), .C2 (n_123_93) );
AOI211_X1 g_101_102 (.ZN (n_101_102), .A (n_105_102), .B (n_111_99), .C1 (n_115_97), .C2 (n_121_94) );
AOI211_X1 g_99_103 (.ZN (n_99_103), .A (n_103_101), .B (n_109_100), .C1 (n_113_98), .C2 (n_119_95) );
AOI211_X1 g_97_104 (.ZN (n_97_104), .A (n_101_102), .B (n_107_101), .C1 (n_111_99), .C2 (n_117_96) );
AOI211_X1 g_95_105 (.ZN (n_95_105), .A (n_99_103), .B (n_105_102), .C1 (n_109_100), .C2 (n_115_97) );
AOI211_X1 g_93_104 (.ZN (n_93_104), .A (n_97_104), .B (n_103_101), .C1 (n_107_101), .C2 (n_113_98) );
AOI211_X1 g_91_105 (.ZN (n_91_105), .A (n_95_105), .B (n_101_102), .C1 (n_105_102), .C2 (n_111_99) );
AOI211_X1 g_92_103 (.ZN (n_92_103), .A (n_93_104), .B (n_99_103), .C1 (n_103_101), .C2 (n_109_100) );
AOI211_X1 g_90_104 (.ZN (n_90_104), .A (n_91_105), .B (n_97_104), .C1 (n_101_102), .C2 (n_107_101) );
AOI211_X1 g_88_105 (.ZN (n_88_105), .A (n_92_103), .B (n_95_105), .C1 (n_99_103), .C2 (n_105_102) );
AOI211_X1 g_86_106 (.ZN (n_86_106), .A (n_90_104), .B (n_93_104), .C1 (n_97_104), .C2 (n_103_101) );
AOI211_X1 g_84_107 (.ZN (n_84_107), .A (n_88_105), .B (n_91_105), .C1 (n_95_105), .C2 (n_101_102) );
AOI211_X1 g_82_108 (.ZN (n_82_108), .A (n_86_106), .B (n_92_103), .C1 (n_93_104), .C2 (n_99_103) );
AOI211_X1 g_80_109 (.ZN (n_80_109), .A (n_84_107), .B (n_90_104), .C1 (n_91_105), .C2 (n_97_104) );
AOI211_X1 g_78_110 (.ZN (n_78_110), .A (n_82_108), .B (n_88_105), .C1 (n_92_103), .C2 (n_95_105) );
AOI211_X1 g_76_111 (.ZN (n_76_111), .A (n_80_109), .B (n_86_106), .C1 (n_90_104), .C2 (n_93_104) );
AOI211_X1 g_74_112 (.ZN (n_74_112), .A (n_78_110), .B (n_84_107), .C1 (n_88_105), .C2 (n_91_105) );
AOI211_X1 g_72_113 (.ZN (n_72_113), .A (n_76_111), .B (n_82_108), .C1 (n_86_106), .C2 (n_92_103) );
AOI211_X1 g_70_114 (.ZN (n_70_114), .A (n_74_112), .B (n_80_109), .C1 (n_84_107), .C2 (n_90_104) );
AOI211_X1 g_68_115 (.ZN (n_68_115), .A (n_72_113), .B (n_78_110), .C1 (n_82_108), .C2 (n_88_105) );
AOI211_X1 g_66_116 (.ZN (n_66_116), .A (n_70_114), .B (n_76_111), .C1 (n_80_109), .C2 (n_86_106) );
AOI211_X1 g_64_117 (.ZN (n_64_117), .A (n_68_115), .B (n_74_112), .C1 (n_78_110), .C2 (n_84_107) );
AOI211_X1 g_62_118 (.ZN (n_62_118), .A (n_66_116), .B (n_72_113), .C1 (n_76_111), .C2 (n_82_108) );
AOI211_X1 g_60_119 (.ZN (n_60_119), .A (n_64_117), .B (n_70_114), .C1 (n_74_112), .C2 (n_80_109) );
AOI211_X1 g_58_120 (.ZN (n_58_120), .A (n_62_118), .B (n_68_115), .C1 (n_72_113), .C2 (n_78_110) );
AOI211_X1 g_56_121 (.ZN (n_56_121), .A (n_60_119), .B (n_66_116), .C1 (n_70_114), .C2 (n_76_111) );
AOI211_X1 g_54_122 (.ZN (n_54_122), .A (n_58_120), .B (n_64_117), .C1 (n_68_115), .C2 (n_74_112) );
AOI211_X1 g_52_123 (.ZN (n_52_123), .A (n_56_121), .B (n_62_118), .C1 (n_66_116), .C2 (n_72_113) );
AOI211_X1 g_51_125 (.ZN (n_51_125), .A (n_54_122), .B (n_60_119), .C1 (n_64_117), .C2 (n_70_114) );
AOI211_X1 g_50_123 (.ZN (n_50_123), .A (n_52_123), .B (n_58_120), .C1 (n_62_118), .C2 (n_68_115) );
AOI211_X1 g_52_122 (.ZN (n_52_122), .A (n_51_125), .B (n_56_121), .C1 (n_60_119), .C2 (n_66_116) );
AOI211_X1 g_54_121 (.ZN (n_54_121), .A (n_50_123), .B (n_54_122), .C1 (n_58_120), .C2 (n_64_117) );
AOI211_X1 g_56_120 (.ZN (n_56_120), .A (n_52_122), .B (n_52_123), .C1 (n_56_121), .C2 (n_62_118) );
AOI211_X1 g_55_122 (.ZN (n_55_122), .A (n_54_121), .B (n_51_125), .C1 (n_54_122), .C2 (n_60_119) );
AOI211_X1 g_57_121 (.ZN (n_57_121), .A (n_56_120), .B (n_50_123), .C1 (n_52_123), .C2 (n_58_120) );
AOI211_X1 g_56_123 (.ZN (n_56_123), .A (n_55_122), .B (n_52_122), .C1 (n_51_125), .C2 (n_56_121) );
AOI211_X1 g_55_121 (.ZN (n_55_121), .A (n_57_121), .B (n_54_121), .C1 (n_50_123), .C2 (n_54_122) );
AOI211_X1 g_57_120 (.ZN (n_57_120), .A (n_56_123), .B (n_56_120), .C1 (n_52_122), .C2 (n_52_123) );
AOI211_X1 g_59_119 (.ZN (n_59_119), .A (n_55_121), .B (n_55_122), .C1 (n_54_121), .C2 (n_51_125) );
AOI211_X1 g_61_118 (.ZN (n_61_118), .A (n_57_120), .B (n_57_121), .C1 (n_56_120), .C2 (n_50_123) );
AOI211_X1 g_63_117 (.ZN (n_63_117), .A (n_59_119), .B (n_56_123), .C1 (n_55_122), .C2 (n_52_122) );
AOI211_X1 g_64_119 (.ZN (n_64_119), .A (n_61_118), .B (n_55_121), .C1 (n_57_121), .C2 (n_54_121) );
AOI211_X1 g_62_120 (.ZN (n_62_120), .A (n_63_117), .B (n_57_120), .C1 (n_56_123), .C2 (n_56_120) );
AOI211_X1 g_60_121 (.ZN (n_60_121), .A (n_64_119), .B (n_59_119), .C1 (n_55_121), .C2 (n_55_122) );
AOI211_X1 g_58_122 (.ZN (n_58_122), .A (n_62_120), .B (n_61_118), .C1 (n_57_120), .C2 (n_57_121) );
AOI211_X1 g_57_124 (.ZN (n_57_124), .A (n_60_121), .B (n_63_117), .C1 (n_59_119), .C2 (n_56_123) );
AOI211_X1 g_56_122 (.ZN (n_56_122), .A (n_58_122), .B (n_64_119), .C1 (n_61_118), .C2 (n_55_121) );
AOI211_X1 g_58_121 (.ZN (n_58_121), .A (n_57_124), .B (n_62_120), .C1 (n_63_117), .C2 (n_57_120) );
AOI211_X1 g_60_120 (.ZN (n_60_120), .A (n_56_122), .B (n_60_121), .C1 (n_64_119), .C2 (n_59_119) );
AOI211_X1 g_62_119 (.ZN (n_62_119), .A (n_58_121), .B (n_58_122), .C1 (n_62_120), .C2 (n_61_118) );
AOI211_X1 g_64_118 (.ZN (n_64_118), .A (n_60_120), .B (n_57_124), .C1 (n_60_121), .C2 (n_63_117) );
AOI211_X1 g_66_117 (.ZN (n_66_117), .A (n_62_119), .B (n_56_122), .C1 (n_58_122), .C2 (n_64_119) );
AOI211_X1 g_68_116 (.ZN (n_68_116), .A (n_64_118), .B (n_58_121), .C1 (n_57_124), .C2 (n_62_120) );
AOI211_X1 g_70_115 (.ZN (n_70_115), .A (n_66_117), .B (n_60_120), .C1 (n_56_122), .C2 (n_60_121) );
AOI211_X1 g_72_114 (.ZN (n_72_114), .A (n_68_116), .B (n_62_119), .C1 (n_58_121), .C2 (n_58_122) );
AOI211_X1 g_74_113 (.ZN (n_74_113), .A (n_70_115), .B (n_64_118), .C1 (n_60_120), .C2 (n_57_124) );
AOI211_X1 g_76_112 (.ZN (n_76_112), .A (n_72_114), .B (n_66_117), .C1 (n_62_119), .C2 (n_56_122) );
AOI211_X1 g_78_111 (.ZN (n_78_111), .A (n_74_113), .B (n_68_116), .C1 (n_64_118), .C2 (n_58_121) );
AOI211_X1 g_80_110 (.ZN (n_80_110), .A (n_76_112), .B (n_70_115), .C1 (n_66_117), .C2 (n_60_120) );
AOI211_X1 g_79_112 (.ZN (n_79_112), .A (n_78_111), .B (n_72_114), .C1 (n_68_116), .C2 (n_62_119) );
AOI211_X1 g_81_111 (.ZN (n_81_111), .A (n_80_110), .B (n_74_113), .C1 (n_70_115), .C2 (n_64_118) );
AOI211_X1 g_83_110 (.ZN (n_83_110), .A (n_79_112), .B (n_76_112), .C1 (n_72_114), .C2 (n_66_117) );
AOI211_X1 g_85_109 (.ZN (n_85_109), .A (n_81_111), .B (n_78_111), .C1 (n_74_113), .C2 (n_68_116) );
AOI211_X1 g_87_108 (.ZN (n_87_108), .A (n_83_110), .B (n_80_110), .C1 (n_76_112), .C2 (n_70_115) );
AOI211_X1 g_89_107 (.ZN (n_89_107), .A (n_85_109), .B (n_79_112), .C1 (n_78_111), .C2 (n_72_114) );
AOI211_X1 g_91_106 (.ZN (n_91_106), .A (n_87_108), .B (n_81_111), .C1 (n_80_110), .C2 (n_74_113) );
AOI211_X1 g_93_105 (.ZN (n_93_105), .A (n_89_107), .B (n_83_110), .C1 (n_79_112), .C2 (n_76_112) );
AOI211_X1 g_95_106 (.ZN (n_95_106), .A (n_91_106), .B (n_85_109), .C1 (n_81_111), .C2 (n_78_111) );
AOI211_X1 g_94_104 (.ZN (n_94_104), .A (n_93_105), .B (n_87_108), .C1 (n_83_110), .C2 (n_80_110) );
AOI211_X1 g_92_105 (.ZN (n_92_105), .A (n_95_106), .B (n_89_107), .C1 (n_85_109), .C2 (n_79_112) );
AOI211_X1 g_90_106 (.ZN (n_90_106), .A (n_94_104), .B (n_91_106), .C1 (n_87_108), .C2 (n_81_111) );
AOI211_X1 g_88_107 (.ZN (n_88_107), .A (n_92_105), .B (n_93_105), .C1 (n_89_107), .C2 (n_83_110) );
AOI211_X1 g_86_108 (.ZN (n_86_108), .A (n_90_106), .B (n_95_106), .C1 (n_91_106), .C2 (n_85_109) );
AOI211_X1 g_84_109 (.ZN (n_84_109), .A (n_88_107), .B (n_94_104), .C1 (n_93_105), .C2 (n_87_108) );
AOI211_X1 g_82_110 (.ZN (n_82_110), .A (n_86_108), .B (n_92_105), .C1 (n_95_106), .C2 (n_89_107) );
AOI211_X1 g_80_111 (.ZN (n_80_111), .A (n_84_109), .B (n_90_106), .C1 (n_94_104), .C2 (n_91_106) );
AOI211_X1 g_78_112 (.ZN (n_78_112), .A (n_82_110), .B (n_88_107), .C1 (n_92_105), .C2 (n_93_105) );
AOI211_X1 g_76_113 (.ZN (n_76_113), .A (n_80_111), .B (n_86_108), .C1 (n_90_106), .C2 (n_95_106) );
AOI211_X1 g_74_114 (.ZN (n_74_114), .A (n_78_112), .B (n_84_109), .C1 (n_88_107), .C2 (n_94_104) );
AOI211_X1 g_72_115 (.ZN (n_72_115), .A (n_76_113), .B (n_82_110), .C1 (n_86_108), .C2 (n_92_105) );
AOI211_X1 g_70_116 (.ZN (n_70_116), .A (n_74_114), .B (n_80_111), .C1 (n_84_109), .C2 (n_90_106) );
AOI211_X1 g_68_117 (.ZN (n_68_117), .A (n_72_115), .B (n_78_112), .C1 (n_82_110), .C2 (n_88_107) );
AOI211_X1 g_67_119 (.ZN (n_67_119), .A (n_70_116), .B (n_76_113), .C1 (n_80_111), .C2 (n_86_108) );
AOI211_X1 g_65_118 (.ZN (n_65_118), .A (n_68_117), .B (n_74_114), .C1 (n_78_112), .C2 (n_84_109) );
AOI211_X1 g_67_117 (.ZN (n_67_117), .A (n_67_119), .B (n_72_115), .C1 (n_76_113), .C2 (n_82_110) );
AOI211_X1 g_69_116 (.ZN (n_69_116), .A (n_65_118), .B (n_70_116), .C1 (n_74_114), .C2 (n_80_111) );
AOI211_X1 g_71_115 (.ZN (n_71_115), .A (n_67_117), .B (n_68_117), .C1 (n_72_115), .C2 (n_78_112) );
AOI211_X1 g_73_114 (.ZN (n_73_114), .A (n_69_116), .B (n_67_119), .C1 (n_70_116), .C2 (n_76_113) );
AOI211_X1 g_75_113 (.ZN (n_75_113), .A (n_71_115), .B (n_65_118), .C1 (n_68_117), .C2 (n_74_114) );
AOI211_X1 g_77_112 (.ZN (n_77_112), .A (n_73_114), .B (n_67_117), .C1 (n_67_119), .C2 (n_72_115) );
AOI211_X1 g_79_111 (.ZN (n_79_111), .A (n_75_113), .B (n_69_116), .C1 (n_65_118), .C2 (n_70_116) );
AOI211_X1 g_81_110 (.ZN (n_81_110), .A (n_77_112), .B (n_71_115), .C1 (n_67_117), .C2 (n_68_117) );
AOI211_X1 g_83_109 (.ZN (n_83_109), .A (n_79_111), .B (n_73_114), .C1 (n_69_116), .C2 (n_67_119) );
AOI211_X1 g_85_108 (.ZN (n_85_108), .A (n_81_110), .B (n_75_113), .C1 (n_71_115), .C2 (n_65_118) );
AOI211_X1 g_87_107 (.ZN (n_87_107), .A (n_83_109), .B (n_77_112), .C1 (n_73_114), .C2 (n_67_117) );
AOI211_X1 g_89_106 (.ZN (n_89_106), .A (n_85_108), .B (n_79_111), .C1 (n_75_113), .C2 (n_69_116) );
AOI211_X1 g_88_108 (.ZN (n_88_108), .A (n_87_107), .B (n_81_110), .C1 (n_77_112), .C2 (n_71_115) );
AOI211_X1 g_90_107 (.ZN (n_90_107), .A (n_89_106), .B (n_83_109), .C1 (n_79_111), .C2 (n_73_114) );
AOI211_X1 g_92_106 (.ZN (n_92_106), .A (n_88_108), .B (n_85_108), .C1 (n_81_110), .C2 (n_75_113) );
AOI211_X1 g_94_105 (.ZN (n_94_105), .A (n_90_107), .B (n_87_107), .C1 (n_83_109), .C2 (n_77_112) );
AOI211_X1 g_93_107 (.ZN (n_93_107), .A (n_92_106), .B (n_89_106), .C1 (n_85_108), .C2 (n_79_111) );
AOI211_X1 g_91_108 (.ZN (n_91_108), .A (n_94_105), .B (n_88_108), .C1 (n_87_107), .C2 (n_81_110) );
AOI211_X1 g_89_109 (.ZN (n_89_109), .A (n_93_107), .B (n_90_107), .C1 (n_89_106), .C2 (n_83_109) );
AOI211_X1 g_87_110 (.ZN (n_87_110), .A (n_91_108), .B (n_92_106), .C1 (n_88_108), .C2 (n_85_108) );
AOI211_X1 g_85_111 (.ZN (n_85_111), .A (n_89_109), .B (n_94_105), .C1 (n_90_107), .C2 (n_87_107) );
AOI211_X1 g_86_109 (.ZN (n_86_109), .A (n_87_110), .B (n_93_107), .C1 (n_92_106), .C2 (n_89_106) );
AOI211_X1 g_84_110 (.ZN (n_84_110), .A (n_85_111), .B (n_91_108), .C1 (n_94_105), .C2 (n_88_108) );
AOI211_X1 g_82_111 (.ZN (n_82_111), .A (n_86_109), .B (n_89_109), .C1 (n_93_107), .C2 (n_90_107) );
AOI211_X1 g_80_112 (.ZN (n_80_112), .A (n_84_110), .B (n_87_110), .C1 (n_91_108), .C2 (n_92_106) );
AOI211_X1 g_78_113 (.ZN (n_78_113), .A (n_82_111), .B (n_85_111), .C1 (n_89_109), .C2 (n_94_105) );
AOI211_X1 g_76_114 (.ZN (n_76_114), .A (n_80_112), .B (n_86_109), .C1 (n_87_110), .C2 (n_93_107) );
AOI211_X1 g_74_115 (.ZN (n_74_115), .A (n_78_113), .B (n_84_110), .C1 (n_85_111), .C2 (n_91_108) );
AOI211_X1 g_72_116 (.ZN (n_72_116), .A (n_76_114), .B (n_82_111), .C1 (n_86_109), .C2 (n_89_109) );
AOI211_X1 g_70_117 (.ZN (n_70_117), .A (n_74_115), .B (n_80_112), .C1 (n_84_110), .C2 (n_87_110) );
AOI211_X1 g_68_118 (.ZN (n_68_118), .A (n_72_116), .B (n_78_113), .C1 (n_82_111), .C2 (n_85_111) );
AOI211_X1 g_66_119 (.ZN (n_66_119), .A (n_70_117), .B (n_76_114), .C1 (n_80_112), .C2 (n_86_109) );
AOI211_X1 g_64_120 (.ZN (n_64_120), .A (n_68_118), .B (n_74_115), .C1 (n_78_113), .C2 (n_84_110) );
AOI211_X1 g_62_121 (.ZN (n_62_121), .A (n_66_119), .B (n_72_116), .C1 (n_76_114), .C2 (n_82_111) );
AOI211_X1 g_63_119 (.ZN (n_63_119), .A (n_64_120), .B (n_70_117), .C1 (n_74_115), .C2 (n_80_112) );
AOI211_X1 g_61_120 (.ZN (n_61_120), .A (n_62_121), .B (n_68_118), .C1 (n_72_116), .C2 (n_78_113) );
AOI211_X1 g_59_121 (.ZN (n_59_121), .A (n_63_119), .B (n_66_119), .C1 (n_70_117), .C2 (n_76_114) );
AOI211_X1 g_57_122 (.ZN (n_57_122), .A (n_61_120), .B (n_64_120), .C1 (n_68_118), .C2 (n_74_115) );
AOI211_X1 g_55_123 (.ZN (n_55_123), .A (n_59_121), .B (n_62_121), .C1 (n_66_119), .C2 (n_72_116) );
AOI211_X1 g_53_122 (.ZN (n_53_122), .A (n_57_122), .B (n_63_119), .C1 (n_64_120), .C2 (n_70_117) );
AOI211_X1 g_51_123 (.ZN (n_51_123), .A (n_55_123), .B (n_61_120), .C1 (n_62_121), .C2 (n_68_118) );
AOI211_X1 g_53_124 (.ZN (n_53_124), .A (n_53_122), .B (n_59_121), .C1 (n_63_119), .C2 (n_66_119) );
AOI211_X1 g_55_125 (.ZN (n_55_125), .A (n_51_123), .B (n_57_122), .C1 (n_61_120), .C2 (n_64_120) );
AOI211_X1 g_54_123 (.ZN (n_54_123), .A (n_53_124), .B (n_55_123), .C1 (n_59_121), .C2 (n_62_121) );
AOI211_X1 g_52_124 (.ZN (n_52_124), .A (n_55_125), .B (n_53_122), .C1 (n_57_122), .C2 (n_63_119) );
AOI211_X1 g_50_125 (.ZN (n_50_125), .A (n_54_123), .B (n_51_123), .C1 (n_55_123), .C2 (n_61_120) );
AOI211_X1 g_48_124 (.ZN (n_48_124), .A (n_52_124), .B (n_53_124), .C1 (n_53_122), .C2 (n_59_121) );
AOI211_X1 g_46_125 (.ZN (n_46_125), .A (n_50_125), .B (n_55_125), .C1 (n_51_123), .C2 (n_57_122) );
AOI211_X1 g_47_123 (.ZN (n_47_123), .A (n_48_124), .B (n_54_123), .C1 (n_53_124), .C2 (n_55_123) );
AOI211_X1 g_49_124 (.ZN (n_49_124), .A (n_46_125), .B (n_52_124), .C1 (n_55_125), .C2 (n_53_122) );
AOI211_X1 g_48_126 (.ZN (n_48_126), .A (n_47_123), .B (n_50_125), .C1 (n_54_123), .C2 (n_51_123) );
AOI211_X1 g_46_127 (.ZN (n_46_127), .A (n_49_124), .B (n_48_124), .C1 (n_52_124), .C2 (n_53_124) );
AOI211_X1 g_47_125 (.ZN (n_47_125), .A (n_48_126), .B (n_46_125), .C1 (n_50_125), .C2 (n_55_125) );
AOI211_X1 g_45_124 (.ZN (n_45_124), .A (n_46_127), .B (n_47_123), .C1 (n_48_124), .C2 (n_54_123) );
AOI211_X1 g_44_126 (.ZN (n_44_126), .A (n_47_125), .B (n_49_124), .C1 (n_46_125), .C2 (n_52_124) );
AOI211_X1 g_42_127 (.ZN (n_42_127), .A (n_45_124), .B (n_48_126), .C1 (n_47_123), .C2 (n_50_125) );
AOI211_X1 g_43_125 (.ZN (n_43_125), .A (n_44_126), .B (n_46_127), .C1 (n_49_124), .C2 (n_48_124) );
AOI211_X1 g_41_126 (.ZN (n_41_126), .A (n_42_127), .B (n_47_125), .C1 (n_48_126), .C2 (n_46_125) );
AOI211_X1 g_39_127 (.ZN (n_39_127), .A (n_43_125), .B (n_45_124), .C1 (n_46_127), .C2 (n_47_123) );
AOI211_X1 g_37_128 (.ZN (n_37_128), .A (n_41_126), .B (n_44_126), .C1 (n_47_125), .C2 (n_49_124) );
AOI211_X1 g_35_129 (.ZN (n_35_129), .A (n_39_127), .B (n_42_127), .C1 (n_45_124), .C2 (n_48_126) );
AOI211_X1 g_33_130 (.ZN (n_33_130), .A (n_37_128), .B (n_43_125), .C1 (n_44_126), .C2 (n_46_127) );
AOI211_X1 g_31_131 (.ZN (n_31_131), .A (n_35_129), .B (n_41_126), .C1 (n_42_127), .C2 (n_47_125) );
AOI211_X1 g_29_132 (.ZN (n_29_132), .A (n_33_130), .B (n_39_127), .C1 (n_43_125), .C2 (n_45_124) );
AOI211_X1 g_27_133 (.ZN (n_27_133), .A (n_31_131), .B (n_37_128), .C1 (n_41_126), .C2 (n_44_126) );
AOI211_X1 g_25_134 (.ZN (n_25_134), .A (n_29_132), .B (n_35_129), .C1 (n_39_127), .C2 (n_42_127) );
AOI211_X1 g_23_135 (.ZN (n_23_135), .A (n_27_133), .B (n_33_130), .C1 (n_37_128), .C2 (n_43_125) );
AOI211_X1 g_21_136 (.ZN (n_21_136), .A (n_25_134), .B (n_31_131), .C1 (n_35_129), .C2 (n_41_126) );
AOI211_X1 g_19_137 (.ZN (n_19_137), .A (n_23_135), .B (n_29_132), .C1 (n_33_130), .C2 (n_39_127) );
AOI211_X1 g_17_138 (.ZN (n_17_138), .A (n_21_136), .B (n_27_133), .C1 (n_31_131), .C2 (n_37_128) );
AOI211_X1 g_15_139 (.ZN (n_15_139), .A (n_19_137), .B (n_25_134), .C1 (n_29_132), .C2 (n_35_129) );
AOI211_X1 g_13_140 (.ZN (n_13_140), .A (n_17_138), .B (n_23_135), .C1 (n_27_133), .C2 (n_33_130) );
AOI211_X1 g_12_142 (.ZN (n_12_142), .A (n_15_139), .B (n_21_136), .C1 (n_25_134), .C2 (n_31_131) );
AOI211_X1 g_11_140 (.ZN (n_11_140), .A (n_13_140), .B (n_19_137), .C1 (n_23_135), .C2 (n_29_132) );
AOI211_X1 g_9_141 (.ZN (n_9_141), .A (n_12_142), .B (n_17_138), .C1 (n_21_136), .C2 (n_27_133) );
AOI211_X1 g_10_143 (.ZN (n_10_143), .A (n_11_140), .B (n_15_139), .C1 (n_19_137), .C2 (n_25_134) );
AOI211_X1 g_9_145 (.ZN (n_9_145), .A (n_9_141), .B (n_13_140), .C1 (n_17_138), .C2 (n_23_135) );
AOI211_X1 g_8_147 (.ZN (n_8_147), .A (n_10_143), .B (n_12_142), .C1 (n_15_139), .C2 (n_21_136) );
AOI211_X1 g_7_145 (.ZN (n_7_145), .A (n_9_145), .B (n_11_140), .C1 (n_13_140), .C2 (n_19_137) );
AOI211_X1 g_8_143 (.ZN (n_8_143), .A (n_8_147), .B (n_9_141), .C1 (n_12_142), .C2 (n_17_138) );
AOI211_X1 g_10_142 (.ZN (n_10_142), .A (n_7_145), .B (n_10_143), .C1 (n_11_140), .C2 (n_15_139) );
AOI211_X1 g_9_144 (.ZN (n_9_144), .A (n_8_143), .B (n_9_145), .C1 (n_9_141), .C2 (n_13_140) );
AOI211_X1 g_11_143 (.ZN (n_11_143), .A (n_10_142), .B (n_8_147), .C1 (n_10_143), .C2 (n_12_142) );
AOI211_X1 g_12_141 (.ZN (n_12_141), .A (n_9_144), .B (n_7_145), .C1 (n_9_145), .C2 (n_11_140) );
AOI211_X1 g_13_139 (.ZN (n_13_139), .A (n_11_143), .B (n_8_143), .C1 (n_8_147), .C2 (n_9_141) );
AOI211_X1 g_15_138 (.ZN (n_15_138), .A (n_12_141), .B (n_10_142), .C1 (n_7_145), .C2 (n_10_143) );
AOI211_X1 g_17_137 (.ZN (n_17_137), .A (n_13_139), .B (n_9_144), .C1 (n_8_143), .C2 (n_9_145) );
AOI211_X1 g_19_136 (.ZN (n_19_136), .A (n_15_138), .B (n_11_143), .C1 (n_10_142), .C2 (n_8_147) );
AOI211_X1 g_21_135 (.ZN (n_21_135), .A (n_17_137), .B (n_12_141), .C1 (n_9_144), .C2 (n_7_145) );
AOI211_X1 g_23_134 (.ZN (n_23_134), .A (n_19_136), .B (n_13_139), .C1 (n_11_143), .C2 (n_8_143) );
AOI211_X1 g_25_135 (.ZN (n_25_135), .A (n_21_135), .B (n_15_138), .C1 (n_12_141), .C2 (n_10_142) );
AOI211_X1 g_23_136 (.ZN (n_23_136), .A (n_23_134), .B (n_17_137), .C1 (n_13_139), .C2 (n_9_144) );
AOI211_X1 g_21_137 (.ZN (n_21_137), .A (n_25_135), .B (n_19_136), .C1 (n_15_138), .C2 (n_11_143) );
AOI211_X1 g_19_138 (.ZN (n_19_138), .A (n_23_136), .B (n_21_135), .C1 (n_17_137), .C2 (n_12_141) );
AOI211_X1 g_17_139 (.ZN (n_17_139), .A (n_21_137), .B (n_23_134), .C1 (n_19_136), .C2 (n_13_139) );
AOI211_X1 g_15_140 (.ZN (n_15_140), .A (n_19_138), .B (n_25_135), .C1 (n_21_135), .C2 (n_15_138) );
AOI211_X1 g_13_141 (.ZN (n_13_141), .A (n_17_139), .B (n_23_136), .C1 (n_23_134), .C2 (n_17_137) );
AOI211_X1 g_11_142 (.ZN (n_11_142), .A (n_15_140), .B (n_21_137), .C1 (n_25_135), .C2 (n_19_136) );
AOI211_X1 g_10_144 (.ZN (n_10_144), .A (n_13_141), .B (n_19_138), .C1 (n_23_136), .C2 (n_21_135) );
AOI211_X1 g_9_146 (.ZN (n_9_146), .A (n_11_142), .B (n_17_139), .C1 (n_21_137), .C2 (n_23_134) );
AOI211_X1 g_10_148 (.ZN (n_10_148), .A (n_10_144), .B (n_15_140), .C1 (n_19_138), .C2 (n_25_135) );
AOI211_X1 g_11_146 (.ZN (n_11_146), .A (n_9_146), .B (n_13_141), .C1 (n_17_139), .C2 (n_23_136) );
AOI211_X1 g_12_144 (.ZN (n_12_144), .A (n_10_148), .B (n_11_142), .C1 (n_15_140), .C2 (n_21_137) );
AOI211_X1 g_13_142 (.ZN (n_13_142), .A (n_11_146), .B (n_10_144), .C1 (n_13_141), .C2 (n_19_138) );
AOI211_X1 g_14_140 (.ZN (n_14_140), .A (n_12_144), .B (n_9_146), .C1 (n_11_142), .C2 (n_17_139) );
AOI211_X1 g_16_139 (.ZN (n_16_139), .A (n_13_142), .B (n_10_148), .C1 (n_10_144), .C2 (n_15_140) );
AOI211_X1 g_18_138 (.ZN (n_18_138), .A (n_14_140), .B (n_11_146), .C1 (n_9_146), .C2 (n_13_141) );
AOI211_X1 g_20_137 (.ZN (n_20_137), .A (n_16_139), .B (n_12_144), .C1 (n_10_148), .C2 (n_11_142) );
AOI211_X1 g_22_136 (.ZN (n_22_136), .A (n_18_138), .B (n_13_142), .C1 (n_11_146), .C2 (n_10_144) );
AOI211_X1 g_24_135 (.ZN (n_24_135), .A (n_20_137), .B (n_14_140), .C1 (n_12_144), .C2 (n_9_146) );
AOI211_X1 g_26_134 (.ZN (n_26_134), .A (n_22_136), .B (n_16_139), .C1 (n_13_142), .C2 (n_10_148) );
AOI211_X1 g_25_136 (.ZN (n_25_136), .A (n_24_135), .B (n_18_138), .C1 (n_14_140), .C2 (n_11_146) );
AOI211_X1 g_27_135 (.ZN (n_27_135), .A (n_26_134), .B (n_20_137), .C1 (n_16_139), .C2 (n_12_144) );
AOI211_X1 g_29_134 (.ZN (n_29_134), .A (n_25_136), .B (n_22_136), .C1 (n_18_138), .C2 (n_13_142) );
AOI211_X1 g_31_133 (.ZN (n_31_133), .A (n_27_135), .B (n_24_135), .C1 (n_20_137), .C2 (n_14_140) );
AOI211_X1 g_33_132 (.ZN (n_33_132), .A (n_29_134), .B (n_26_134), .C1 (n_22_136), .C2 (n_16_139) );
AOI211_X1 g_35_131 (.ZN (n_35_131), .A (n_31_133), .B (n_25_136), .C1 (n_24_135), .C2 (n_18_138) );
AOI211_X1 g_37_130 (.ZN (n_37_130), .A (n_33_132), .B (n_27_135), .C1 (n_26_134), .C2 (n_20_137) );
AOI211_X1 g_39_129 (.ZN (n_39_129), .A (n_35_131), .B (n_29_134), .C1 (n_25_136), .C2 (n_22_136) );
AOI211_X1 g_41_128 (.ZN (n_41_128), .A (n_37_130), .B (n_31_133), .C1 (n_27_135), .C2 (n_24_135) );
AOI211_X1 g_43_127 (.ZN (n_43_127), .A (n_39_129), .B (n_33_132), .C1 (n_29_134), .C2 (n_26_134) );
AOI211_X1 g_45_126 (.ZN (n_45_126), .A (n_41_128), .B (n_35_131), .C1 (n_31_133), .C2 (n_25_136) );
AOI211_X1 g_44_128 (.ZN (n_44_128), .A (n_43_127), .B (n_37_130), .C1 (n_33_132), .C2 (n_27_135) );
AOI211_X1 g_42_129 (.ZN (n_42_129), .A (n_45_126), .B (n_39_129), .C1 (n_35_131), .C2 (n_29_134) );
AOI211_X1 g_40_128 (.ZN (n_40_128), .A (n_44_128), .B (n_41_128), .C1 (n_37_130), .C2 (n_31_133) );
AOI211_X1 g_38_129 (.ZN (n_38_129), .A (n_42_129), .B (n_43_127), .C1 (n_39_129), .C2 (n_33_132) );
AOI211_X1 g_36_130 (.ZN (n_36_130), .A (n_40_128), .B (n_45_126), .C1 (n_41_128), .C2 (n_35_131) );
AOI211_X1 g_34_131 (.ZN (n_34_131), .A (n_38_129), .B (n_44_128), .C1 (n_43_127), .C2 (n_37_130) );
AOI211_X1 g_32_132 (.ZN (n_32_132), .A (n_36_130), .B (n_42_129), .C1 (n_45_126), .C2 (n_39_129) );
AOI211_X1 g_30_133 (.ZN (n_30_133), .A (n_34_131), .B (n_40_128), .C1 (n_44_128), .C2 (n_41_128) );
AOI211_X1 g_28_134 (.ZN (n_28_134), .A (n_32_132), .B (n_38_129), .C1 (n_42_129), .C2 (n_43_127) );
AOI211_X1 g_26_135 (.ZN (n_26_135), .A (n_30_133), .B (n_36_130), .C1 (n_40_128), .C2 (n_45_126) );
AOI211_X1 g_24_136 (.ZN (n_24_136), .A (n_28_134), .B (n_34_131), .C1 (n_38_129), .C2 (n_44_128) );
AOI211_X1 g_22_137 (.ZN (n_22_137), .A (n_26_135), .B (n_32_132), .C1 (n_36_130), .C2 (n_42_129) );
AOI211_X1 g_20_138 (.ZN (n_20_138), .A (n_24_136), .B (n_30_133), .C1 (n_34_131), .C2 (n_40_128) );
AOI211_X1 g_18_139 (.ZN (n_18_139), .A (n_22_137), .B (n_28_134), .C1 (n_32_132), .C2 (n_38_129) );
AOI211_X1 g_16_140 (.ZN (n_16_140), .A (n_20_138), .B (n_26_135), .C1 (n_30_133), .C2 (n_36_130) );
AOI211_X1 g_14_141 (.ZN (n_14_141), .A (n_18_139), .B (n_24_136), .C1 (n_28_134), .C2 (n_34_131) );
AOI211_X1 g_13_143 (.ZN (n_13_143), .A (n_16_140), .B (n_22_137), .C1 (n_26_135), .C2 (n_32_132) );
AOI211_X1 g_11_144 (.ZN (n_11_144), .A (n_14_141), .B (n_20_138), .C1 (n_24_136), .C2 (n_30_133) );
AOI211_X1 g_13_145 (.ZN (n_13_145), .A (n_13_143), .B (n_18_139), .C1 (n_22_137), .C2 (n_28_134) );
AOI211_X1 g_12_143 (.ZN (n_12_143), .A (n_11_144), .B (n_16_140), .C1 (n_20_138), .C2 (n_26_135) );
AOI211_X1 g_11_145 (.ZN (n_11_145), .A (n_13_145), .B (n_14_141), .C1 (n_18_139), .C2 (n_24_136) );
AOI211_X1 g_12_147 (.ZN (n_12_147), .A (n_12_143), .B (n_13_143), .C1 (n_16_140), .C2 (n_22_137) );
AOI211_X1 g_14_148 (.ZN (n_14_148), .A (n_11_145), .B (n_11_144), .C1 (n_14_141), .C2 (n_20_138) );
AOI211_X1 g_12_149 (.ZN (n_12_149), .A (n_12_147), .B (n_13_145), .C1 (n_13_143), .C2 (n_18_139) );
AOI211_X1 g_11_147 (.ZN (n_11_147), .A (n_14_148), .B (n_12_143), .C1 (n_11_144), .C2 (n_16_140) );
AOI211_X1 g_13_146 (.ZN (n_13_146), .A (n_12_149), .B (n_11_145), .C1 (n_13_145), .C2 (n_14_141) );
AOI211_X1 g_14_144 (.ZN (n_14_144), .A (n_11_147), .B (n_12_147), .C1 (n_12_143), .C2 (n_13_143) );
AOI211_X1 g_12_145 (.ZN (n_12_145), .A (n_13_146), .B (n_14_148), .C1 (n_11_145), .C2 (n_11_144) );
AOI211_X1 g_13_147 (.ZN (n_13_147), .A (n_14_144), .B (n_12_149), .C1 (n_12_147), .C2 (n_13_145) );
AOI211_X1 g_15_146 (.ZN (n_15_146), .A (n_12_145), .B (n_11_147), .C1 (n_14_148), .C2 (n_12_143) );
AOI211_X1 g_17_145 (.ZN (n_17_145), .A (n_13_147), .B (n_13_146), .C1 (n_12_149), .C2 (n_11_145) );
AOI211_X1 g_16_147 (.ZN (n_16_147), .A (n_15_146), .B (n_14_144), .C1 (n_11_147), .C2 (n_12_147) );
AOI211_X1 g_15_145 (.ZN (n_15_145), .A (n_17_145), .B (n_12_145), .C1 (n_13_146), .C2 (n_14_148) );
AOI211_X1 g_14_143 (.ZN (n_14_143), .A (n_16_147), .B (n_13_147), .C1 (n_14_144), .C2 (n_12_149) );
AOI211_X1 g_15_141 (.ZN (n_15_141), .A (n_15_145), .B (n_15_146), .C1 (n_12_145), .C2 (n_11_147) );
AOI211_X1 g_17_140 (.ZN (n_17_140), .A (n_14_143), .B (n_17_145), .C1 (n_13_147), .C2 (n_13_146) );
AOI211_X1 g_19_139 (.ZN (n_19_139), .A (n_15_141), .B (n_16_147), .C1 (n_15_146), .C2 (n_14_144) );
AOI211_X1 g_21_138 (.ZN (n_21_138), .A (n_17_140), .B (n_15_145), .C1 (n_17_145), .C2 (n_12_145) );
AOI211_X1 g_23_137 (.ZN (n_23_137), .A (n_19_139), .B (n_14_143), .C1 (n_16_147), .C2 (n_13_147) );
AOI211_X1 g_22_139 (.ZN (n_22_139), .A (n_21_138), .B (n_15_141), .C1 (n_15_145), .C2 (n_15_146) );
AOI211_X1 g_24_138 (.ZN (n_24_138), .A (n_23_137), .B (n_17_140), .C1 (n_14_143), .C2 (n_17_145) );
AOI211_X1 g_26_137 (.ZN (n_26_137), .A (n_22_139), .B (n_19_139), .C1 (n_15_141), .C2 (n_16_147) );
AOI211_X1 g_28_136 (.ZN (n_28_136), .A (n_24_138), .B (n_21_138), .C1 (n_17_140), .C2 (n_15_145) );
AOI211_X1 g_30_135 (.ZN (n_30_135), .A (n_26_137), .B (n_23_137), .C1 (n_19_139), .C2 (n_14_143) );
AOI211_X1 g_32_134 (.ZN (n_32_134), .A (n_28_136), .B (n_22_139), .C1 (n_21_138), .C2 (n_15_141) );
AOI211_X1 g_34_133 (.ZN (n_34_133), .A (n_30_135), .B (n_24_138), .C1 (n_23_137), .C2 (n_17_140) );
AOI211_X1 g_36_132 (.ZN (n_36_132), .A (n_32_134), .B (n_26_137), .C1 (n_22_139), .C2 (n_19_139) );
AOI211_X1 g_38_131 (.ZN (n_38_131), .A (n_34_133), .B (n_28_136), .C1 (n_24_138), .C2 (n_21_138) );
AOI211_X1 g_40_130 (.ZN (n_40_130), .A (n_36_132), .B (n_30_135), .C1 (n_26_137), .C2 (n_23_137) );
AOI211_X1 g_39_132 (.ZN (n_39_132), .A (n_38_131), .B (n_32_134), .C1 (n_28_136), .C2 (n_22_139) );
AOI211_X1 g_38_130 (.ZN (n_38_130), .A (n_40_130), .B (n_34_133), .C1 (n_30_135), .C2 (n_24_138) );
AOI211_X1 g_40_129 (.ZN (n_40_129), .A (n_39_132), .B (n_36_132), .C1 (n_32_134), .C2 (n_26_137) );
AOI211_X1 g_42_128 (.ZN (n_42_128), .A (n_38_130), .B (n_38_131), .C1 (n_34_133), .C2 (n_28_136) );
AOI211_X1 g_44_127 (.ZN (n_44_127), .A (n_40_129), .B (n_40_130), .C1 (n_36_132), .C2 (n_30_135) );
AOI211_X1 g_46_126 (.ZN (n_46_126), .A (n_42_128), .B (n_39_132), .C1 (n_38_131), .C2 (n_32_134) );
AOI211_X1 g_48_125 (.ZN (n_48_125), .A (n_44_127), .B (n_38_130), .C1 (n_40_130), .C2 (n_34_133) );
AOI211_X1 g_47_127 (.ZN (n_47_127), .A (n_46_126), .B (n_40_129), .C1 (n_39_132), .C2 (n_36_132) );
AOI211_X1 g_49_126 (.ZN (n_49_126), .A (n_48_125), .B (n_42_128), .C1 (n_38_130), .C2 (n_38_131) );
AOI211_X1 g_48_128 (.ZN (n_48_128), .A (n_47_127), .B (n_44_127), .C1 (n_40_129), .C2 (n_40_130) );
AOI211_X1 g_47_126 (.ZN (n_47_126), .A (n_49_126), .B (n_46_126), .C1 (n_42_128), .C2 (n_39_132) );
AOI211_X1 g_49_125 (.ZN (n_49_125), .A (n_48_128), .B (n_48_125), .C1 (n_44_127), .C2 (n_38_130) );
AOI211_X1 g_51_124 (.ZN (n_51_124), .A (n_47_126), .B (n_47_127), .C1 (n_46_126), .C2 (n_40_129) );
AOI211_X1 g_53_123 (.ZN (n_53_123), .A (n_49_125), .B (n_49_126), .C1 (n_48_125), .C2 (n_42_128) );
AOI211_X1 g_52_125 (.ZN (n_52_125), .A (n_51_124), .B (n_48_128), .C1 (n_47_127), .C2 (n_44_127) );
AOI211_X1 g_54_124 (.ZN (n_54_124), .A (n_53_123), .B (n_47_126), .C1 (n_49_126), .C2 (n_46_126) );
AOI211_X1 g_53_126 (.ZN (n_53_126), .A (n_52_125), .B (n_49_125), .C1 (n_48_128), .C2 (n_48_125) );
AOI211_X1 g_51_127 (.ZN (n_51_127), .A (n_54_124), .B (n_51_124), .C1 (n_47_126), .C2 (n_47_127) );
AOI211_X1 g_49_128 (.ZN (n_49_128), .A (n_53_126), .B (n_53_123), .C1 (n_49_125), .C2 (n_49_126) );
AOI211_X1 g_50_126 (.ZN (n_50_126), .A (n_51_127), .B (n_52_125), .C1 (n_51_124), .C2 (n_48_128) );
AOI211_X1 g_48_127 (.ZN (n_48_127), .A (n_49_128), .B (n_54_124), .C1 (n_53_123), .C2 (n_47_126) );
AOI211_X1 g_46_128 (.ZN (n_46_128), .A (n_50_126), .B (n_53_126), .C1 (n_52_125), .C2 (n_49_125) );
AOI211_X1 g_44_129 (.ZN (n_44_129), .A (n_48_127), .B (n_51_127), .C1 (n_54_124), .C2 (n_51_124) );
AOI211_X1 g_45_127 (.ZN (n_45_127), .A (n_46_128), .B (n_49_128), .C1 (n_53_126), .C2 (n_53_123) );
AOI211_X1 g_43_128 (.ZN (n_43_128), .A (n_44_129), .B (n_50_126), .C1 (n_51_127), .C2 (n_52_125) );
AOI211_X1 g_41_129 (.ZN (n_41_129), .A (n_45_127), .B (n_48_127), .C1 (n_49_128), .C2 (n_54_124) );
AOI211_X1 g_39_130 (.ZN (n_39_130), .A (n_43_128), .B (n_46_128), .C1 (n_50_126), .C2 (n_53_126) );
AOI211_X1 g_37_131 (.ZN (n_37_131), .A (n_41_129), .B (n_44_129), .C1 (n_48_127), .C2 (n_51_127) );
AOI211_X1 g_35_132 (.ZN (n_35_132), .A (n_39_130), .B (n_45_127), .C1 (n_46_128), .C2 (n_49_128) );
AOI211_X1 g_33_133 (.ZN (n_33_133), .A (n_37_131), .B (n_43_128), .C1 (n_44_129), .C2 (n_50_126) );
AOI211_X1 g_31_134 (.ZN (n_31_134), .A (n_35_132), .B (n_41_129), .C1 (n_45_127), .C2 (n_48_127) );
AOI211_X1 g_29_135 (.ZN (n_29_135), .A (n_33_133), .B (n_39_130), .C1 (n_43_128), .C2 (n_46_128) );
AOI211_X1 g_27_136 (.ZN (n_27_136), .A (n_31_134), .B (n_37_131), .C1 (n_41_129), .C2 (n_44_129) );
AOI211_X1 g_25_137 (.ZN (n_25_137), .A (n_29_135), .B (n_35_132), .C1 (n_39_130), .C2 (n_45_127) );
AOI211_X1 g_23_138 (.ZN (n_23_138), .A (n_27_136), .B (n_33_133), .C1 (n_37_131), .C2 (n_43_128) );
AOI211_X1 g_21_139 (.ZN (n_21_139), .A (n_25_137), .B (n_31_134), .C1 (n_35_132), .C2 (n_41_129) );
AOI211_X1 g_19_140 (.ZN (n_19_140), .A (n_23_138), .B (n_29_135), .C1 (n_33_133), .C2 (n_39_130) );
AOI211_X1 g_17_141 (.ZN (n_17_141), .A (n_21_139), .B (n_27_136), .C1 (n_31_134), .C2 (n_37_131) );
AOI211_X1 g_15_142 (.ZN (n_15_142), .A (n_19_140), .B (n_25_137), .C1 (n_29_135), .C2 (n_35_132) );
AOI211_X1 g_16_144 (.ZN (n_16_144), .A (n_17_141), .B (n_23_138), .C1 (n_27_136), .C2 (n_33_133) );
AOI211_X1 g_14_145 (.ZN (n_14_145), .A (n_15_142), .B (n_21_139), .C1 (n_25_137), .C2 (n_31_134) );
AOI211_X1 g_15_143 (.ZN (n_15_143), .A (n_16_144), .B (n_19_140), .C1 (n_23_138), .C2 (n_29_135) );
AOI211_X1 g_13_144 (.ZN (n_13_144), .A (n_14_145), .B (n_17_141), .C1 (n_21_139), .C2 (n_27_136) );
AOI211_X1 g_14_142 (.ZN (n_14_142), .A (n_15_143), .B (n_15_142), .C1 (n_19_140), .C2 (n_25_137) );
AOI211_X1 g_16_143 (.ZN (n_16_143), .A (n_13_144), .B (n_16_144), .C1 (n_17_141), .C2 (n_23_138) );
AOI211_X1 g_18_142 (.ZN (n_18_142), .A (n_14_142), .B (n_14_145), .C1 (n_15_142), .C2 (n_21_139) );
AOI211_X1 g_16_141 (.ZN (n_16_141), .A (n_16_143), .B (n_15_143), .C1 (n_16_144), .C2 (n_19_140) );
AOI211_X1 g_18_140 (.ZN (n_18_140), .A (n_18_142), .B (n_13_144), .C1 (n_14_145), .C2 (n_17_141) );
AOI211_X1 g_17_142 (.ZN (n_17_142), .A (n_16_141), .B (n_14_142), .C1 (n_15_143), .C2 (n_15_142) );
AOI211_X1 g_19_141 (.ZN (n_19_141), .A (n_18_140), .B (n_16_143), .C1 (n_13_144), .C2 (n_16_144) );
AOI211_X1 g_20_139 (.ZN (n_20_139), .A (n_17_142), .B (n_18_142), .C1 (n_14_142), .C2 (n_14_145) );
AOI211_X1 g_22_138 (.ZN (n_22_138), .A (n_19_141), .B (n_16_141), .C1 (n_16_143), .C2 (n_15_143) );
AOI211_X1 g_24_137 (.ZN (n_24_137), .A (n_20_139), .B (n_18_140), .C1 (n_18_142), .C2 (n_13_144) );
AOI211_X1 g_26_136 (.ZN (n_26_136), .A (n_22_138), .B (n_17_142), .C1 (n_16_141), .C2 (n_14_142) );
AOI211_X1 g_28_135 (.ZN (n_28_135), .A (n_24_137), .B (n_19_141), .C1 (n_18_140), .C2 (n_16_143) );
AOI211_X1 g_30_134 (.ZN (n_30_134), .A (n_26_136), .B (n_20_139), .C1 (n_17_142), .C2 (n_18_142) );
AOI211_X1 g_32_133 (.ZN (n_32_133), .A (n_28_135), .B (n_22_138), .C1 (n_19_141), .C2 (n_16_141) );
AOI211_X1 g_34_132 (.ZN (n_34_132), .A (n_30_134), .B (n_24_137), .C1 (n_20_139), .C2 (n_18_140) );
AOI211_X1 g_36_131 (.ZN (n_36_131), .A (n_32_133), .B (n_26_136), .C1 (n_22_138), .C2 (n_17_142) );
AOI211_X1 g_37_133 (.ZN (n_37_133), .A (n_34_132), .B (n_28_135), .C1 (n_24_137), .C2 (n_19_141) );
AOI211_X1 g_35_134 (.ZN (n_35_134), .A (n_36_131), .B (n_30_134), .C1 (n_26_136), .C2 (n_20_139) );
AOI211_X1 g_33_135 (.ZN (n_33_135), .A (n_37_133), .B (n_32_133), .C1 (n_28_135), .C2 (n_22_138) );
AOI211_X1 g_31_136 (.ZN (n_31_136), .A (n_35_134), .B (n_34_132), .C1 (n_30_134), .C2 (n_24_137) );
AOI211_X1 g_29_137 (.ZN (n_29_137), .A (n_33_135), .B (n_36_131), .C1 (n_32_133), .C2 (n_26_136) );
AOI211_X1 g_27_138 (.ZN (n_27_138), .A (n_31_136), .B (n_37_133), .C1 (n_34_132), .C2 (n_28_135) );
AOI211_X1 g_25_139 (.ZN (n_25_139), .A (n_29_137), .B (n_35_134), .C1 (n_36_131), .C2 (n_30_134) );
AOI211_X1 g_23_140 (.ZN (n_23_140), .A (n_27_138), .B (n_33_135), .C1 (n_37_133), .C2 (n_32_133) );
AOI211_X1 g_21_141 (.ZN (n_21_141), .A (n_25_139), .B (n_31_136), .C1 (n_35_134), .C2 (n_34_132) );
AOI211_X1 g_19_142 (.ZN (n_19_142), .A (n_23_140), .B (n_29_137), .C1 (n_33_135), .C2 (n_36_131) );
AOI211_X1 g_20_140 (.ZN (n_20_140), .A (n_21_141), .B (n_27_138), .C1 (n_31_136), .C2 (n_37_133) );
AOI211_X1 g_18_141 (.ZN (n_18_141), .A (n_19_142), .B (n_25_139), .C1 (n_29_137), .C2 (n_35_134) );
AOI211_X1 g_16_142 (.ZN (n_16_142), .A (n_20_140), .B (n_23_140), .C1 (n_27_138), .C2 (n_33_135) );
AOI211_X1 g_15_144 (.ZN (n_15_144), .A (n_18_141), .B (n_21_141), .C1 (n_25_139), .C2 (n_31_136) );
AOI211_X1 g_17_143 (.ZN (n_17_143), .A (n_16_142), .B (n_19_142), .C1 (n_23_140), .C2 (n_29_137) );
AOI211_X1 g_16_145 (.ZN (n_16_145), .A (n_15_144), .B (n_20_140), .C1 (n_21_141), .C2 (n_27_138) );
AOI211_X1 g_14_146 (.ZN (n_14_146), .A (n_17_143), .B (n_18_141), .C1 (n_19_142), .C2 (n_25_139) );
AOI211_X1 g_13_148 (.ZN (n_13_148), .A (n_16_145), .B (n_16_142), .C1 (n_20_140), .C2 (n_23_140) );
AOI211_X1 g_14_150 (.ZN (n_14_150), .A (n_14_146), .B (n_15_144), .C1 (n_18_141), .C2 (n_21_141) );
AOI211_X1 g_15_148 (.ZN (n_15_148), .A (n_13_148), .B (n_17_143), .C1 (n_16_142), .C2 (n_19_142) );
AOI211_X1 g_16_146 (.ZN (n_16_146), .A (n_14_150), .B (n_16_145), .C1 (n_15_144), .C2 (n_20_140) );
AOI211_X1 g_17_144 (.ZN (n_17_144), .A (n_15_148), .B (n_14_146), .C1 (n_17_143), .C2 (n_18_141) );
AOI211_X1 g_19_143 (.ZN (n_19_143), .A (n_16_146), .B (n_13_148), .C1 (n_16_145), .C2 (n_16_142) );
AOI211_X1 g_20_141 (.ZN (n_20_141), .A (n_17_144), .B (n_14_150), .C1 (n_14_146), .C2 (n_15_144) );
AOI211_X1 g_22_140 (.ZN (n_22_140), .A (n_19_143), .B (n_15_148), .C1 (n_13_148), .C2 (n_17_143) );
AOI211_X1 g_24_139 (.ZN (n_24_139), .A (n_20_141), .B (n_16_146), .C1 (n_14_150), .C2 (n_16_145) );
AOI211_X1 g_26_138 (.ZN (n_26_138), .A (n_22_140), .B (n_17_144), .C1 (n_15_148), .C2 (n_14_146) );
AOI211_X1 g_28_137 (.ZN (n_28_137), .A (n_24_139), .B (n_19_143), .C1 (n_16_146), .C2 (n_13_148) );
AOI211_X1 g_30_136 (.ZN (n_30_136), .A (n_26_138), .B (n_20_141), .C1 (n_17_144), .C2 (n_14_150) );
AOI211_X1 g_32_135 (.ZN (n_32_135), .A (n_28_137), .B (n_22_140), .C1 (n_19_143), .C2 (n_15_148) );
AOI211_X1 g_34_134 (.ZN (n_34_134), .A (n_30_136), .B (n_24_139), .C1 (n_20_141), .C2 (n_16_146) );
AOI211_X1 g_36_133 (.ZN (n_36_133), .A (n_32_135), .B (n_26_138), .C1 (n_22_140), .C2 (n_17_144) );
AOI211_X1 g_38_132 (.ZN (n_38_132), .A (n_34_134), .B (n_28_137), .C1 (n_24_139), .C2 (n_19_143) );
AOI211_X1 g_40_131 (.ZN (n_40_131), .A (n_36_133), .B (n_30_136), .C1 (n_26_138), .C2 (n_20_141) );
AOI211_X1 g_42_130 (.ZN (n_42_130), .A (n_38_132), .B (n_32_135), .C1 (n_28_137), .C2 (n_22_140) );
AOI211_X1 g_41_132 (.ZN (n_41_132), .A (n_40_131), .B (n_34_134), .C1 (n_30_136), .C2 (n_24_139) );
AOI211_X1 g_39_131 (.ZN (n_39_131), .A (n_42_130), .B (n_36_133), .C1 (n_32_135), .C2 (n_26_138) );
AOI211_X1 g_41_130 (.ZN (n_41_130), .A (n_41_132), .B (n_38_132), .C1 (n_34_134), .C2 (n_28_137) );
AOI211_X1 g_43_129 (.ZN (n_43_129), .A (n_39_131), .B (n_40_131), .C1 (n_36_133), .C2 (n_30_136) );
AOI211_X1 g_45_128 (.ZN (n_45_128), .A (n_41_130), .B (n_42_130), .C1 (n_38_132), .C2 (n_32_135) );
AOI211_X1 g_47_129 (.ZN (n_47_129), .A (n_43_129), .B (n_41_132), .C1 (n_40_131), .C2 (n_34_134) );
AOI211_X1 g_45_130 (.ZN (n_45_130), .A (n_45_128), .B (n_39_131), .C1 (n_42_130), .C2 (n_36_133) );
AOI211_X1 g_43_131 (.ZN (n_43_131), .A (n_47_129), .B (n_41_130), .C1 (n_41_132), .C2 (n_38_132) );
AOI211_X1 g_42_133 (.ZN (n_42_133), .A (n_45_130), .B (n_43_129), .C1 (n_39_131), .C2 (n_40_131) );
AOI211_X1 g_41_131 (.ZN (n_41_131), .A (n_43_131), .B (n_45_128), .C1 (n_41_130), .C2 (n_42_130) );
AOI211_X1 g_43_130 (.ZN (n_43_130), .A (n_42_133), .B (n_47_129), .C1 (n_43_129), .C2 (n_41_132) );
AOI211_X1 g_45_129 (.ZN (n_45_129), .A (n_41_131), .B (n_45_130), .C1 (n_45_128), .C2 (n_39_131) );
AOI211_X1 g_47_128 (.ZN (n_47_128), .A (n_43_130), .B (n_43_131), .C1 (n_47_129), .C2 (n_41_130) );
AOI211_X1 g_49_127 (.ZN (n_49_127), .A (n_45_129), .B (n_42_133), .C1 (n_45_130), .C2 (n_43_129) );
AOI211_X1 g_51_126 (.ZN (n_51_126), .A (n_47_128), .B (n_41_131), .C1 (n_43_131), .C2 (n_45_128) );
AOI211_X1 g_53_125 (.ZN (n_53_125), .A (n_49_127), .B (n_43_130), .C1 (n_42_133), .C2 (n_47_129) );
AOI211_X1 g_55_124 (.ZN (n_55_124), .A (n_51_126), .B (n_45_129), .C1 (n_41_131), .C2 (n_45_130) );
AOI211_X1 g_57_123 (.ZN (n_57_123), .A (n_53_125), .B (n_47_128), .C1 (n_43_130), .C2 (n_43_131) );
AOI211_X1 g_59_122 (.ZN (n_59_122), .A (n_55_124), .B (n_49_127), .C1 (n_45_129), .C2 (n_42_133) );
AOI211_X1 g_61_121 (.ZN (n_61_121), .A (n_57_123), .B (n_51_126), .C1 (n_47_128), .C2 (n_41_131) );
AOI211_X1 g_63_120 (.ZN (n_63_120), .A (n_59_122), .B (n_53_125), .C1 (n_49_127), .C2 (n_43_130) );
AOI211_X1 g_65_119 (.ZN (n_65_119), .A (n_61_121), .B (n_55_124), .C1 (n_51_126), .C2 (n_45_129) );
AOI211_X1 g_67_118 (.ZN (n_67_118), .A (n_63_120), .B (n_57_123), .C1 (n_53_125), .C2 (n_47_128) );
AOI211_X1 g_69_117 (.ZN (n_69_117), .A (n_65_119), .B (n_59_122), .C1 (n_55_124), .C2 (n_49_127) );
AOI211_X1 g_71_116 (.ZN (n_71_116), .A (n_67_118), .B (n_61_121), .C1 (n_57_123), .C2 (n_51_126) );
AOI211_X1 g_73_115 (.ZN (n_73_115), .A (n_69_117), .B (n_63_120), .C1 (n_59_122), .C2 (n_53_125) );
AOI211_X1 g_75_114 (.ZN (n_75_114), .A (n_71_116), .B (n_65_119), .C1 (n_61_121), .C2 (n_55_124) );
AOI211_X1 g_77_113 (.ZN (n_77_113), .A (n_73_115), .B (n_67_118), .C1 (n_63_120), .C2 (n_57_123) );
AOI211_X1 g_76_115 (.ZN (n_76_115), .A (n_75_114), .B (n_69_117), .C1 (n_65_119), .C2 (n_59_122) );
AOI211_X1 g_78_114 (.ZN (n_78_114), .A (n_77_113), .B (n_71_116), .C1 (n_67_118), .C2 (n_61_121) );
AOI211_X1 g_80_113 (.ZN (n_80_113), .A (n_76_115), .B (n_73_115), .C1 (n_69_117), .C2 (n_63_120) );
AOI211_X1 g_82_112 (.ZN (n_82_112), .A (n_78_114), .B (n_75_114), .C1 (n_71_116), .C2 (n_65_119) );
AOI211_X1 g_84_111 (.ZN (n_84_111), .A (n_80_113), .B (n_77_113), .C1 (n_73_115), .C2 (n_67_118) );
AOI211_X1 g_86_110 (.ZN (n_86_110), .A (n_82_112), .B (n_76_115), .C1 (n_75_114), .C2 (n_69_117) );
AOI211_X1 g_88_109 (.ZN (n_88_109), .A (n_84_111), .B (n_78_114), .C1 (n_77_113), .C2 (n_71_116) );
AOI211_X1 g_90_108 (.ZN (n_90_108), .A (n_86_110), .B (n_80_113), .C1 (n_76_115), .C2 (n_73_115) );
AOI211_X1 g_92_107 (.ZN (n_92_107), .A (n_88_109), .B (n_82_112), .C1 (n_78_114), .C2 (n_75_114) );
AOI211_X1 g_94_106 (.ZN (n_94_106), .A (n_90_108), .B (n_84_111), .C1 (n_80_113), .C2 (n_77_113) );
AOI211_X1 g_96_105 (.ZN (n_96_105), .A (n_92_107), .B (n_86_110), .C1 (n_82_112), .C2 (n_76_115) );
AOI211_X1 g_98_104 (.ZN (n_98_104), .A (n_94_106), .B (n_88_109), .C1 (n_84_111), .C2 (n_78_114) );
AOI211_X1 g_100_103 (.ZN (n_100_103), .A (n_96_105), .B (n_90_108), .C1 (n_86_110), .C2 (n_80_113) );
AOI211_X1 g_102_102 (.ZN (n_102_102), .A (n_98_104), .B (n_92_107), .C1 (n_88_109), .C2 (n_82_112) );
AOI211_X1 g_101_104 (.ZN (n_101_104), .A (n_100_103), .B (n_94_106), .C1 (n_90_108), .C2 (n_84_111) );
AOI211_X1 g_103_103 (.ZN (n_103_103), .A (n_102_102), .B (n_96_105), .C1 (n_92_107), .C2 (n_86_110) );
AOI211_X1 g_102_105 (.ZN (n_102_105), .A (n_101_104), .B (n_98_104), .C1 (n_94_106), .C2 (n_88_109) );
AOI211_X1 g_100_104 (.ZN (n_100_104), .A (n_103_103), .B (n_100_103), .C1 (n_96_105), .C2 (n_90_108) );
AOI211_X1 g_102_103 (.ZN (n_102_103), .A (n_102_105), .B (n_102_102), .C1 (n_98_104), .C2 (n_92_107) );
AOI211_X1 g_104_104 (.ZN (n_104_104), .A (n_100_104), .B (n_101_104), .C1 (n_100_103), .C2 (n_94_106) );
AOI211_X1 g_106_103 (.ZN (n_106_103), .A (n_102_103), .B (n_103_103), .C1 (n_102_102), .C2 (n_96_105) );
AOI211_X1 g_108_102 (.ZN (n_108_102), .A (n_104_104), .B (n_102_105), .C1 (n_101_104), .C2 (n_98_104) );
AOI211_X1 g_110_101 (.ZN (n_110_101), .A (n_106_103), .B (n_100_104), .C1 (n_103_103), .C2 (n_100_103) );
AOI211_X1 g_112_100 (.ZN (n_112_100), .A (n_108_102), .B (n_102_103), .C1 (n_102_105), .C2 (n_102_102) );
AOI211_X1 g_114_99 (.ZN (n_114_99), .A (n_110_101), .B (n_104_104), .C1 (n_100_104), .C2 (n_101_104) );
AOI211_X1 g_116_98 (.ZN (n_116_98), .A (n_112_100), .B (n_106_103), .C1 (n_102_103), .C2 (n_103_103) );
AOI211_X1 g_118_97 (.ZN (n_118_97), .A (n_114_99), .B (n_108_102), .C1 (n_104_104), .C2 (n_102_105) );
AOI211_X1 g_120_96 (.ZN (n_120_96), .A (n_116_98), .B (n_110_101), .C1 (n_106_103), .C2 (n_100_104) );
AOI211_X1 g_122_95 (.ZN (n_122_95), .A (n_118_97), .B (n_112_100), .C1 (n_108_102), .C2 (n_102_103) );
AOI211_X1 g_124_94 (.ZN (n_124_94), .A (n_120_96), .B (n_114_99), .C1 (n_110_101), .C2 (n_104_104) );
AOI211_X1 g_126_93 (.ZN (n_126_93), .A (n_122_95), .B (n_116_98), .C1 (n_112_100), .C2 (n_106_103) );
AOI211_X1 g_128_92 (.ZN (n_128_92), .A (n_124_94), .B (n_118_97), .C1 (n_114_99), .C2 (n_108_102) );
AOI211_X1 g_130_91 (.ZN (n_130_91), .A (n_126_93), .B (n_120_96), .C1 (n_116_98), .C2 (n_110_101) );
AOI211_X1 g_132_90 (.ZN (n_132_90), .A (n_128_92), .B (n_122_95), .C1 (n_118_97), .C2 (n_112_100) );
AOI211_X1 g_134_89 (.ZN (n_134_89), .A (n_130_91), .B (n_124_94), .C1 (n_120_96), .C2 (n_114_99) );
AOI211_X1 g_136_88 (.ZN (n_136_88), .A (n_132_90), .B (n_126_93), .C1 (n_122_95), .C2 (n_116_98) );
AOI211_X1 g_138_87 (.ZN (n_138_87), .A (n_134_89), .B (n_128_92), .C1 (n_124_94), .C2 (n_118_97) );
AOI211_X1 g_140_86 (.ZN (n_140_86), .A (n_136_88), .B (n_130_91), .C1 (n_126_93), .C2 (n_120_96) );
AOI211_X1 g_142_85 (.ZN (n_142_85), .A (n_138_87), .B (n_132_90), .C1 (n_128_92), .C2 (n_122_95) );
AOI211_X1 g_141_87 (.ZN (n_141_87), .A (n_140_86), .B (n_134_89), .C1 (n_130_91), .C2 (n_124_94) );
AOI211_X1 g_139_88 (.ZN (n_139_88), .A (n_142_85), .B (n_136_88), .C1 (n_132_90), .C2 (n_126_93) );
AOI211_X1 g_137_89 (.ZN (n_137_89), .A (n_141_87), .B (n_138_87), .C1 (n_134_89), .C2 (n_128_92) );
AOI211_X1 g_135_90 (.ZN (n_135_90), .A (n_139_88), .B (n_140_86), .C1 (n_136_88), .C2 (n_130_91) );
AOI211_X1 g_133_91 (.ZN (n_133_91), .A (n_137_89), .B (n_142_85), .C1 (n_138_87), .C2 (n_132_90) );
AOI211_X1 g_131_92 (.ZN (n_131_92), .A (n_135_90), .B (n_141_87), .C1 (n_140_86), .C2 (n_134_89) );
AOI211_X1 g_129_93 (.ZN (n_129_93), .A (n_133_91), .B (n_139_88), .C1 (n_142_85), .C2 (n_136_88) );
AOI211_X1 g_127_94 (.ZN (n_127_94), .A (n_131_92), .B (n_137_89), .C1 (n_141_87), .C2 (n_138_87) );
AOI211_X1 g_125_95 (.ZN (n_125_95), .A (n_129_93), .B (n_135_90), .C1 (n_139_88), .C2 (n_140_86) );
AOI211_X1 g_123_96 (.ZN (n_123_96), .A (n_127_94), .B (n_133_91), .C1 (n_137_89), .C2 (n_142_85) );
AOI211_X1 g_122_94 (.ZN (n_122_94), .A (n_125_95), .B (n_131_92), .C1 (n_135_90), .C2 (n_141_87) );
AOI211_X1 g_120_95 (.ZN (n_120_95), .A (n_123_96), .B (n_129_93), .C1 (n_133_91), .C2 (n_139_88) );
AOI211_X1 g_118_96 (.ZN (n_118_96), .A (n_122_94), .B (n_127_94), .C1 (n_131_92), .C2 (n_137_89) );
AOI211_X1 g_116_97 (.ZN (n_116_97), .A (n_120_95), .B (n_125_95), .C1 (n_129_93), .C2 (n_135_90) );
AOI211_X1 g_114_98 (.ZN (n_114_98), .A (n_118_96), .B (n_123_96), .C1 (n_127_94), .C2 (n_133_91) );
AOI211_X1 g_112_99 (.ZN (n_112_99), .A (n_116_97), .B (n_122_94), .C1 (n_125_95), .C2 (n_131_92) );
AOI211_X1 g_110_100 (.ZN (n_110_100), .A (n_114_98), .B (n_120_95), .C1 (n_123_96), .C2 (n_129_93) );
AOI211_X1 g_108_101 (.ZN (n_108_101), .A (n_112_99), .B (n_118_96), .C1 (n_122_94), .C2 (n_127_94) );
AOI211_X1 g_106_102 (.ZN (n_106_102), .A (n_110_100), .B (n_116_97), .C1 (n_120_95), .C2 (n_125_95) );
AOI211_X1 g_104_103 (.ZN (n_104_103), .A (n_108_101), .B (n_114_98), .C1 (n_118_96), .C2 (n_123_96) );
AOI211_X1 g_102_104 (.ZN (n_102_104), .A (n_106_102), .B (n_112_99), .C1 (n_116_97), .C2 (n_122_94) );
AOI211_X1 g_100_105 (.ZN (n_100_105), .A (n_104_103), .B (n_110_100), .C1 (n_114_98), .C2 (n_120_95) );
AOI211_X1 g_98_106 (.ZN (n_98_106), .A (n_102_104), .B (n_108_101), .C1 (n_112_99), .C2 (n_118_96) );
AOI211_X1 g_96_107 (.ZN (n_96_107), .A (n_100_105), .B (n_106_102), .C1 (n_110_100), .C2 (n_116_97) );
AOI211_X1 g_94_108 (.ZN (n_94_108), .A (n_98_106), .B (n_104_103), .C1 (n_108_101), .C2 (n_114_98) );
AOI211_X1 g_93_106 (.ZN (n_93_106), .A (n_96_107), .B (n_102_104), .C1 (n_106_102), .C2 (n_112_99) );
AOI211_X1 g_91_107 (.ZN (n_91_107), .A (n_94_108), .B (n_100_105), .C1 (n_104_103), .C2 (n_110_100) );
AOI211_X1 g_89_108 (.ZN (n_89_108), .A (n_93_106), .B (n_98_106), .C1 (n_102_104), .C2 (n_108_101) );
AOI211_X1 g_87_109 (.ZN (n_87_109), .A (n_91_107), .B (n_96_107), .C1 (n_100_105), .C2 (n_106_102) );
AOI211_X1 g_85_110 (.ZN (n_85_110), .A (n_89_108), .B (n_94_108), .C1 (n_98_106), .C2 (n_104_103) );
AOI211_X1 g_83_111 (.ZN (n_83_111), .A (n_87_109), .B (n_93_106), .C1 (n_96_107), .C2 (n_102_104) );
AOI211_X1 g_81_112 (.ZN (n_81_112), .A (n_85_110), .B (n_91_107), .C1 (n_94_108), .C2 (n_100_105) );
AOI211_X1 g_79_113 (.ZN (n_79_113), .A (n_83_111), .B (n_89_108), .C1 (n_93_106), .C2 (n_98_106) );
AOI211_X1 g_77_114 (.ZN (n_77_114), .A (n_81_112), .B (n_87_109), .C1 (n_91_107), .C2 (n_96_107) );
AOI211_X1 g_75_115 (.ZN (n_75_115), .A (n_79_113), .B (n_85_110), .C1 (n_89_108), .C2 (n_94_108) );
AOI211_X1 g_73_116 (.ZN (n_73_116), .A (n_77_114), .B (n_83_111), .C1 (n_87_109), .C2 (n_93_106) );
AOI211_X1 g_71_117 (.ZN (n_71_117), .A (n_75_115), .B (n_81_112), .C1 (n_85_110), .C2 (n_91_107) );
AOI211_X1 g_69_118 (.ZN (n_69_118), .A (n_73_116), .B (n_79_113), .C1 (n_83_111), .C2 (n_89_108) );
AOI211_X1 g_68_120 (.ZN (n_68_120), .A (n_71_117), .B (n_77_114), .C1 (n_81_112), .C2 (n_87_109) );
AOI211_X1 g_70_119 (.ZN (n_70_119), .A (n_69_118), .B (n_75_115), .C1 (n_79_113), .C2 (n_85_110) );
AOI211_X1 g_72_118 (.ZN (n_72_118), .A (n_68_120), .B (n_73_116), .C1 (n_77_114), .C2 (n_83_111) );
AOI211_X1 g_74_117 (.ZN (n_74_117), .A (n_70_119), .B (n_71_117), .C1 (n_75_115), .C2 (n_81_112) );
AOI211_X1 g_76_116 (.ZN (n_76_116), .A (n_72_118), .B (n_69_118), .C1 (n_73_116), .C2 (n_79_113) );
AOI211_X1 g_78_115 (.ZN (n_78_115), .A (n_74_117), .B (n_68_120), .C1 (n_71_117), .C2 (n_77_114) );
AOI211_X1 g_80_114 (.ZN (n_80_114), .A (n_76_116), .B (n_70_119), .C1 (n_69_118), .C2 (n_75_115) );
AOI211_X1 g_82_113 (.ZN (n_82_113), .A (n_78_115), .B (n_72_118), .C1 (n_68_120), .C2 (n_73_116) );
AOI211_X1 g_84_112 (.ZN (n_84_112), .A (n_80_114), .B (n_74_117), .C1 (n_70_119), .C2 (n_71_117) );
AOI211_X1 g_86_111 (.ZN (n_86_111), .A (n_82_113), .B (n_76_116), .C1 (n_72_118), .C2 (n_69_118) );
AOI211_X1 g_88_110 (.ZN (n_88_110), .A (n_84_112), .B (n_78_115), .C1 (n_74_117), .C2 (n_68_120) );
AOI211_X1 g_90_109 (.ZN (n_90_109), .A (n_86_111), .B (n_80_114), .C1 (n_76_116), .C2 (n_70_119) );
AOI211_X1 g_92_108 (.ZN (n_92_108), .A (n_88_110), .B (n_82_113), .C1 (n_78_115), .C2 (n_72_118) );
AOI211_X1 g_94_107 (.ZN (n_94_107), .A (n_90_109), .B (n_84_112), .C1 (n_80_114), .C2 (n_74_117) );
AOI211_X1 g_96_106 (.ZN (n_96_106), .A (n_92_108), .B (n_86_111), .C1 (n_82_113), .C2 (n_76_116) );
AOI211_X1 g_98_105 (.ZN (n_98_105), .A (n_94_107), .B (n_88_110), .C1 (n_84_112), .C2 (n_78_115) );
AOI211_X1 g_100_106 (.ZN (n_100_106), .A (n_96_106), .B (n_90_109), .C1 (n_86_111), .C2 (n_80_114) );
AOI211_X1 g_98_107 (.ZN (n_98_107), .A (n_98_105), .B (n_92_108), .C1 (n_88_110), .C2 (n_82_113) );
AOI211_X1 g_99_105 (.ZN (n_99_105), .A (n_100_106), .B (n_94_107), .C1 (n_90_109), .C2 (n_84_112) );
AOI211_X1 g_97_106 (.ZN (n_97_106), .A (n_98_107), .B (n_96_106), .C1 (n_92_108), .C2 (n_86_111) );
AOI211_X1 g_95_107 (.ZN (n_95_107), .A (n_99_105), .B (n_98_105), .C1 (n_94_107), .C2 (n_88_110) );
AOI211_X1 g_93_108 (.ZN (n_93_108), .A (n_97_106), .B (n_100_106), .C1 (n_96_106), .C2 (n_90_109) );
AOI211_X1 g_91_109 (.ZN (n_91_109), .A (n_95_107), .B (n_98_107), .C1 (n_98_105), .C2 (n_92_108) );
AOI211_X1 g_89_110 (.ZN (n_89_110), .A (n_93_108), .B (n_99_105), .C1 (n_100_106), .C2 (n_94_107) );
AOI211_X1 g_87_111 (.ZN (n_87_111), .A (n_91_109), .B (n_97_106), .C1 (n_98_107), .C2 (n_96_106) );
AOI211_X1 g_85_112 (.ZN (n_85_112), .A (n_89_110), .B (n_95_107), .C1 (n_99_105), .C2 (n_98_105) );
AOI211_X1 g_83_113 (.ZN (n_83_113), .A (n_87_111), .B (n_93_108), .C1 (n_97_106), .C2 (n_100_106) );
AOI211_X1 g_81_114 (.ZN (n_81_114), .A (n_85_112), .B (n_91_109), .C1 (n_95_107), .C2 (n_98_107) );
AOI211_X1 g_79_115 (.ZN (n_79_115), .A (n_83_113), .B (n_89_110), .C1 (n_93_108), .C2 (n_99_105) );
AOI211_X1 g_77_116 (.ZN (n_77_116), .A (n_81_114), .B (n_87_111), .C1 (n_91_109), .C2 (n_97_106) );
AOI211_X1 g_75_117 (.ZN (n_75_117), .A (n_79_115), .B (n_85_112), .C1 (n_89_110), .C2 (n_95_107) );
AOI211_X1 g_73_118 (.ZN (n_73_118), .A (n_77_116), .B (n_83_113), .C1 (n_87_111), .C2 (n_93_108) );
AOI211_X1 g_74_116 (.ZN (n_74_116), .A (n_75_117), .B (n_81_114), .C1 (n_85_112), .C2 (n_91_109) );
AOI211_X1 g_72_117 (.ZN (n_72_117), .A (n_73_118), .B (n_79_115), .C1 (n_83_113), .C2 (n_89_110) );
AOI211_X1 g_70_118 (.ZN (n_70_118), .A (n_74_116), .B (n_77_116), .C1 (n_81_114), .C2 (n_87_111) );
AOI211_X1 g_68_119 (.ZN (n_68_119), .A (n_72_117), .B (n_75_117), .C1 (n_79_115), .C2 (n_85_112) );
AOI211_X1 g_66_120 (.ZN (n_66_120), .A (n_70_118), .B (n_73_118), .C1 (n_77_116), .C2 (n_83_113) );
AOI211_X1 g_64_121 (.ZN (n_64_121), .A (n_68_119), .B (n_74_116), .C1 (n_75_117), .C2 (n_81_114) );
AOI211_X1 g_62_122 (.ZN (n_62_122), .A (n_66_120), .B (n_72_117), .C1 (n_73_118), .C2 (n_79_115) );
AOI211_X1 g_60_123 (.ZN (n_60_123), .A (n_64_121), .B (n_70_118), .C1 (n_74_116), .C2 (n_77_116) );
AOI211_X1 g_58_124 (.ZN (n_58_124), .A (n_62_122), .B (n_68_119), .C1 (n_72_117), .C2 (n_75_117) );
AOI211_X1 g_56_125 (.ZN (n_56_125), .A (n_60_123), .B (n_66_120), .C1 (n_70_118), .C2 (n_73_118) );
AOI211_X1 g_54_126 (.ZN (n_54_126), .A (n_58_124), .B (n_64_121), .C1 (n_68_119), .C2 (n_74_116) );
AOI211_X1 g_52_127 (.ZN (n_52_127), .A (n_56_125), .B (n_62_122), .C1 (n_66_120), .C2 (n_72_117) );
AOI211_X1 g_50_128 (.ZN (n_50_128), .A (n_54_126), .B (n_60_123), .C1 (n_64_121), .C2 (n_70_118) );
AOI211_X1 g_48_129 (.ZN (n_48_129), .A (n_52_127), .B (n_58_124), .C1 (n_62_122), .C2 (n_68_119) );
AOI211_X1 g_46_130 (.ZN (n_46_130), .A (n_50_128), .B (n_56_125), .C1 (n_60_123), .C2 (n_66_120) );
AOI211_X1 g_44_131 (.ZN (n_44_131), .A (n_48_129), .B (n_54_126), .C1 (n_58_124), .C2 (n_64_121) );
AOI211_X1 g_42_132 (.ZN (n_42_132), .A (n_46_130), .B (n_52_127), .C1 (n_56_125), .C2 (n_62_122) );
AOI211_X1 g_40_133 (.ZN (n_40_133), .A (n_44_131), .B (n_50_128), .C1 (n_54_126), .C2 (n_60_123) );
AOI211_X1 g_38_134 (.ZN (n_38_134), .A (n_42_132), .B (n_48_129), .C1 (n_52_127), .C2 (n_58_124) );
AOI211_X1 g_37_132 (.ZN (n_37_132), .A (n_40_133), .B (n_46_130), .C1 (n_50_128), .C2 (n_56_125) );
AOI211_X1 g_35_133 (.ZN (n_35_133), .A (n_38_134), .B (n_44_131), .C1 (n_48_129), .C2 (n_54_126) );
AOI211_X1 g_33_134 (.ZN (n_33_134), .A (n_37_132), .B (n_42_132), .C1 (n_46_130), .C2 (n_52_127) );
AOI211_X1 g_31_135 (.ZN (n_31_135), .A (n_35_133), .B (n_40_133), .C1 (n_44_131), .C2 (n_50_128) );
AOI211_X1 g_29_136 (.ZN (n_29_136), .A (n_33_134), .B (n_38_134), .C1 (n_42_132), .C2 (n_48_129) );
AOI211_X1 g_27_137 (.ZN (n_27_137), .A (n_31_135), .B (n_37_132), .C1 (n_40_133), .C2 (n_46_130) );
AOI211_X1 g_25_138 (.ZN (n_25_138), .A (n_29_136), .B (n_35_133), .C1 (n_38_134), .C2 (n_44_131) );
AOI211_X1 g_23_139 (.ZN (n_23_139), .A (n_27_137), .B (n_33_134), .C1 (n_37_132), .C2 (n_42_132) );
AOI211_X1 g_21_140 (.ZN (n_21_140), .A (n_25_138), .B (n_31_135), .C1 (n_35_133), .C2 (n_40_133) );
AOI211_X1 g_20_142 (.ZN (n_20_142), .A (n_23_139), .B (n_29_136), .C1 (n_33_134), .C2 (n_38_134) );
AOI211_X1 g_18_143 (.ZN (n_18_143), .A (n_21_140), .B (n_27_137), .C1 (n_31_135), .C2 (n_37_132) );
AOI211_X1 g_19_145 (.ZN (n_19_145), .A (n_20_142), .B (n_25_138), .C1 (n_29_136), .C2 (n_35_133) );
AOI211_X1 g_20_143 (.ZN (n_20_143), .A (n_18_143), .B (n_23_139), .C1 (n_27_137), .C2 (n_33_134) );
AOI211_X1 g_18_144 (.ZN (n_18_144), .A (n_19_145), .B (n_21_140), .C1 (n_25_138), .C2 (n_31_135) );
AOI211_X1 g_17_146 (.ZN (n_17_146), .A (n_20_143), .B (n_20_142), .C1 (n_23_139), .C2 (n_29_136) );
AOI211_X1 g_15_147 (.ZN (n_15_147), .A (n_18_144), .B (n_18_143), .C1 (n_21_140), .C2 (n_27_137) );
AOI211_X1 g_16_149 (.ZN (n_16_149), .A (n_17_146), .B (n_19_145), .C1 (n_20_142), .C2 (n_25_138) );
AOI211_X1 g_18_148 (.ZN (n_18_148), .A (n_15_147), .B (n_20_143), .C1 (n_18_143), .C2 (n_23_139) );
AOI211_X1 g_20_147 (.ZN (n_20_147), .A (n_16_149), .B (n_18_144), .C1 (n_19_145), .C2 (n_21_140) );
AOI211_X1 g_18_146 (.ZN (n_18_146), .A (n_18_148), .B (n_17_146), .C1 (n_20_143), .C2 (n_20_142) );
AOI211_X1 g_17_148 (.ZN (n_17_148), .A (n_20_147), .B (n_15_147), .C1 (n_18_144), .C2 (n_18_143) );
AOI211_X1 g_18_150 (.ZN (n_18_150), .A (n_18_146), .B (n_16_149), .C1 (n_17_146), .C2 (n_19_145) );
AOI211_X1 g_19_148 (.ZN (n_19_148), .A (n_17_148), .B (n_18_148), .C1 (n_15_147), .C2 (n_20_143) );
AOI211_X1 g_17_147 (.ZN (n_17_147), .A (n_18_150), .B (n_20_147), .C1 (n_16_149), .C2 (n_18_144) );
AOI211_X1 g_19_146 (.ZN (n_19_146), .A (n_19_148), .B (n_18_146), .C1 (n_18_148), .C2 (n_17_146) );
AOI211_X1 g_21_145 (.ZN (n_21_145), .A (n_17_147), .B (n_17_148), .C1 (n_20_147), .C2 (n_15_147) );
AOI211_X1 g_19_144 (.ZN (n_19_144), .A (n_19_146), .B (n_18_150), .C1 (n_18_146), .C2 (n_16_149) );
AOI211_X1 g_20_146 (.ZN (n_20_146), .A (n_21_145), .B (n_19_148), .C1 (n_17_148), .C2 (n_18_148) );
AOI211_X1 g_18_145 (.ZN (n_18_145), .A (n_19_144), .B (n_17_147), .C1 (n_18_150), .C2 (n_20_147) );
AOI211_X1 g_20_144 (.ZN (n_20_144), .A (n_20_146), .B (n_19_146), .C1 (n_19_148), .C2 (n_18_146) );
AOI211_X1 g_21_142 (.ZN (n_21_142), .A (n_18_145), .B (n_21_145), .C1 (n_17_147), .C2 (n_17_148) );
AOI211_X1 g_23_141 (.ZN (n_23_141), .A (n_20_144), .B (n_19_144), .C1 (n_19_146), .C2 (n_18_150) );
AOI211_X1 g_22_143 (.ZN (n_22_143), .A (n_21_142), .B (n_20_146), .C1 (n_21_145), .C2 (n_19_148) );
AOI211_X1 g_24_142 (.ZN (n_24_142), .A (n_23_141), .B (n_18_145), .C1 (n_19_144), .C2 (n_17_147) );
AOI211_X1 g_25_140 (.ZN (n_25_140), .A (n_22_143), .B (n_20_144), .C1 (n_20_146), .C2 (n_19_146) );
AOI211_X1 g_27_139 (.ZN (n_27_139), .A (n_24_142), .B (n_21_142), .C1 (n_18_145), .C2 (n_21_145) );
AOI211_X1 g_29_138 (.ZN (n_29_138), .A (n_25_140), .B (n_23_141), .C1 (n_20_144), .C2 (n_19_144) );
AOI211_X1 g_31_137 (.ZN (n_31_137), .A (n_27_139), .B (n_22_143), .C1 (n_21_142), .C2 (n_20_146) );
AOI211_X1 g_33_136 (.ZN (n_33_136), .A (n_29_138), .B (n_24_142), .C1 (n_23_141), .C2 (n_18_145) );
AOI211_X1 g_35_135 (.ZN (n_35_135), .A (n_31_137), .B (n_25_140), .C1 (n_22_143), .C2 (n_20_144) );
AOI211_X1 g_37_134 (.ZN (n_37_134), .A (n_33_136), .B (n_27_139), .C1 (n_24_142), .C2 (n_21_142) );
AOI211_X1 g_39_133 (.ZN (n_39_133), .A (n_35_135), .B (n_29_138), .C1 (n_25_140), .C2 (n_23_141) );
AOI211_X1 g_38_135 (.ZN (n_38_135), .A (n_37_134), .B (n_31_137), .C1 (n_27_139), .C2 (n_22_143) );
AOI211_X1 g_40_134 (.ZN (n_40_134), .A (n_39_133), .B (n_33_136), .C1 (n_29_138), .C2 (n_24_142) );
AOI211_X1 g_38_133 (.ZN (n_38_133), .A (n_38_135), .B (n_35_135), .C1 (n_31_137), .C2 (n_25_140) );
AOI211_X1 g_40_132 (.ZN (n_40_132), .A (n_40_134), .B (n_37_134), .C1 (n_33_136), .C2 (n_27_139) );
AOI211_X1 g_42_131 (.ZN (n_42_131), .A (n_38_133), .B (n_39_133), .C1 (n_35_135), .C2 (n_29_138) );
AOI211_X1 g_44_130 (.ZN (n_44_130), .A (n_40_132), .B (n_38_135), .C1 (n_37_134), .C2 (n_31_137) );
AOI211_X1 g_46_129 (.ZN (n_46_129), .A (n_42_131), .B (n_40_134), .C1 (n_39_133), .C2 (n_33_136) );
AOI211_X1 g_45_131 (.ZN (n_45_131), .A (n_44_130), .B (n_38_133), .C1 (n_38_135), .C2 (n_35_135) );
AOI211_X1 g_47_130 (.ZN (n_47_130), .A (n_46_129), .B (n_40_132), .C1 (n_40_134), .C2 (n_37_134) );
AOI211_X1 g_49_129 (.ZN (n_49_129), .A (n_45_131), .B (n_42_131), .C1 (n_38_133), .C2 (n_39_133) );
AOI211_X1 g_50_127 (.ZN (n_50_127), .A (n_47_130), .B (n_44_130), .C1 (n_40_132), .C2 (n_38_135) );
AOI211_X1 g_52_126 (.ZN (n_52_126), .A (n_49_129), .B (n_46_129), .C1 (n_42_131), .C2 (n_40_134) );
AOI211_X1 g_54_125 (.ZN (n_54_125), .A (n_50_127), .B (n_45_131), .C1 (n_44_130), .C2 (n_38_133) );
AOI211_X1 g_56_124 (.ZN (n_56_124), .A (n_52_126), .B (n_47_130), .C1 (n_46_129), .C2 (n_40_132) );
AOI211_X1 g_58_123 (.ZN (n_58_123), .A (n_54_125), .B (n_49_129), .C1 (n_45_131), .C2 (n_42_131) );
AOI211_X1 g_60_122 (.ZN (n_60_122), .A (n_56_124), .B (n_50_127), .C1 (n_47_130), .C2 (n_44_130) );
AOI211_X1 g_59_124 (.ZN (n_59_124), .A (n_58_123), .B (n_52_126), .C1 (n_49_129), .C2 (n_46_129) );
AOI211_X1 g_61_123 (.ZN (n_61_123), .A (n_60_122), .B (n_54_125), .C1 (n_50_127), .C2 (n_45_131) );
AOI211_X1 g_63_122 (.ZN (n_63_122), .A (n_59_124), .B (n_56_124), .C1 (n_52_126), .C2 (n_47_130) );
AOI211_X1 g_65_121 (.ZN (n_65_121), .A (n_61_123), .B (n_58_123), .C1 (n_54_125), .C2 (n_49_129) );
AOI211_X1 g_67_120 (.ZN (n_67_120), .A (n_63_122), .B (n_60_122), .C1 (n_56_124), .C2 (n_50_127) );
AOI211_X1 g_69_119 (.ZN (n_69_119), .A (n_65_121), .B (n_59_124), .C1 (n_58_123), .C2 (n_52_126) );
AOI211_X1 g_71_118 (.ZN (n_71_118), .A (n_67_120), .B (n_61_123), .C1 (n_60_122), .C2 (n_54_125) );
AOI211_X1 g_73_117 (.ZN (n_73_117), .A (n_69_119), .B (n_63_122), .C1 (n_59_124), .C2 (n_56_124) );
AOI211_X1 g_75_116 (.ZN (n_75_116), .A (n_71_118), .B (n_65_121), .C1 (n_61_123), .C2 (n_58_123) );
AOI211_X1 g_77_115 (.ZN (n_77_115), .A (n_73_117), .B (n_67_120), .C1 (n_63_122), .C2 (n_60_122) );
AOI211_X1 g_79_114 (.ZN (n_79_114), .A (n_75_116), .B (n_69_119), .C1 (n_65_121), .C2 (n_59_124) );
AOI211_X1 g_81_113 (.ZN (n_81_113), .A (n_77_115), .B (n_71_118), .C1 (n_67_120), .C2 (n_61_123) );
AOI211_X1 g_83_112 (.ZN (n_83_112), .A (n_79_114), .B (n_73_117), .C1 (n_69_119), .C2 (n_63_122) );
AOI211_X1 g_82_114 (.ZN (n_82_114), .A (n_81_113), .B (n_75_116), .C1 (n_71_118), .C2 (n_65_121) );
AOI211_X1 g_84_113 (.ZN (n_84_113), .A (n_83_112), .B (n_77_115), .C1 (n_73_117), .C2 (n_67_120) );
AOI211_X1 g_86_112 (.ZN (n_86_112), .A (n_82_114), .B (n_79_114), .C1 (n_75_116), .C2 (n_69_119) );
AOI211_X1 g_88_111 (.ZN (n_88_111), .A (n_84_113), .B (n_81_113), .C1 (n_77_115), .C2 (n_71_118) );
AOI211_X1 g_90_110 (.ZN (n_90_110), .A (n_86_112), .B (n_83_112), .C1 (n_79_114), .C2 (n_73_117) );
AOI211_X1 g_92_109 (.ZN (n_92_109), .A (n_88_111), .B (n_82_114), .C1 (n_81_113), .C2 (n_75_116) );
AOI211_X1 g_91_111 (.ZN (n_91_111), .A (n_90_110), .B (n_84_113), .C1 (n_83_112), .C2 (n_77_115) );
AOI211_X1 g_93_110 (.ZN (n_93_110), .A (n_92_109), .B (n_86_112), .C1 (n_82_114), .C2 (n_79_114) );
AOI211_X1 g_95_109 (.ZN (n_95_109), .A (n_91_111), .B (n_88_111), .C1 (n_84_113), .C2 (n_81_113) );
AOI211_X1 g_97_108 (.ZN (n_97_108), .A (n_93_110), .B (n_90_110), .C1 (n_86_112), .C2 (n_83_112) );
AOI211_X1 g_99_107 (.ZN (n_99_107), .A (n_95_109), .B (n_92_109), .C1 (n_88_111), .C2 (n_82_114) );
AOI211_X1 g_101_106 (.ZN (n_101_106), .A (n_97_108), .B (n_91_111), .C1 (n_90_110), .C2 (n_84_113) );
AOI211_X1 g_103_105 (.ZN (n_103_105), .A (n_99_107), .B (n_93_110), .C1 (n_92_109), .C2 (n_86_112) );
AOI211_X1 g_105_104 (.ZN (n_105_104), .A (n_101_106), .B (n_95_109), .C1 (n_91_111), .C2 (n_88_111) );
AOI211_X1 g_107_103 (.ZN (n_107_103), .A (n_103_105), .B (n_97_108), .C1 (n_93_110), .C2 (n_90_110) );
AOI211_X1 g_109_102 (.ZN (n_109_102), .A (n_105_104), .B (n_99_107), .C1 (n_95_109), .C2 (n_92_109) );
AOI211_X1 g_111_101 (.ZN (n_111_101), .A (n_107_103), .B (n_101_106), .C1 (n_97_108), .C2 (n_91_111) );
AOI211_X1 g_113_100 (.ZN (n_113_100), .A (n_109_102), .B (n_103_105), .C1 (n_99_107), .C2 (n_93_110) );
AOI211_X1 g_115_99 (.ZN (n_115_99), .A (n_111_101), .B (n_105_104), .C1 (n_101_106), .C2 (n_95_109) );
AOI211_X1 g_117_98 (.ZN (n_117_98), .A (n_113_100), .B (n_107_103), .C1 (n_103_105), .C2 (n_97_108) );
AOI211_X1 g_119_97 (.ZN (n_119_97), .A (n_115_99), .B (n_109_102), .C1 (n_105_104), .C2 (n_99_107) );
AOI211_X1 g_121_96 (.ZN (n_121_96), .A (n_117_98), .B (n_111_101), .C1 (n_107_103), .C2 (n_101_106) );
AOI211_X1 g_123_95 (.ZN (n_123_95), .A (n_119_97), .B (n_113_100), .C1 (n_109_102), .C2 (n_103_105) );
AOI211_X1 g_125_94 (.ZN (n_125_94), .A (n_121_96), .B (n_115_99), .C1 (n_111_101), .C2 (n_105_104) );
AOI211_X1 g_127_93 (.ZN (n_127_93), .A (n_123_95), .B (n_117_98), .C1 (n_113_100), .C2 (n_107_103) );
AOI211_X1 g_129_92 (.ZN (n_129_92), .A (n_125_94), .B (n_119_97), .C1 (n_115_99), .C2 (n_109_102) );
AOI211_X1 g_131_91 (.ZN (n_131_91), .A (n_127_93), .B (n_121_96), .C1 (n_117_98), .C2 (n_111_101) );
AOI211_X1 g_133_90 (.ZN (n_133_90), .A (n_129_92), .B (n_123_95), .C1 (n_119_97), .C2 (n_113_100) );
AOI211_X1 g_135_89 (.ZN (n_135_89), .A (n_131_91), .B (n_125_94), .C1 (n_121_96), .C2 (n_115_99) );
AOI211_X1 g_137_88 (.ZN (n_137_88), .A (n_133_90), .B (n_127_93), .C1 (n_123_95), .C2 (n_117_98) );
AOI211_X1 g_136_90 (.ZN (n_136_90), .A (n_135_89), .B (n_129_92), .C1 (n_125_94), .C2 (n_119_97) );
AOI211_X1 g_138_89 (.ZN (n_138_89), .A (n_137_88), .B (n_131_91), .C1 (n_127_93), .C2 (n_121_96) );
AOI211_X1 g_140_88 (.ZN (n_140_88), .A (n_136_90), .B (n_133_90), .C1 (n_129_92), .C2 (n_123_95) );
AOI211_X1 g_142_87 (.ZN (n_142_87), .A (n_138_89), .B (n_135_89), .C1 (n_131_91), .C2 (n_125_94) );
AOI211_X1 g_144_86 (.ZN (n_144_86), .A (n_140_88), .B (n_137_88), .C1 (n_133_90), .C2 (n_127_93) );
AOI211_X1 g_146_87 (.ZN (n_146_87), .A (n_142_87), .B (n_136_90), .C1 (n_135_89), .C2 (n_129_92) );
AOI211_X1 g_144_88 (.ZN (n_144_88), .A (n_144_86), .B (n_138_89), .C1 (n_137_88), .C2 (n_131_91) );
AOI211_X1 g_142_89 (.ZN (n_142_89), .A (n_146_87), .B (n_140_88), .C1 (n_136_90), .C2 (n_133_90) );
AOI211_X1 g_143_87 (.ZN (n_143_87), .A (n_144_88), .B (n_142_87), .C1 (n_138_89), .C2 (n_135_89) );
AOI211_X1 g_144_89 (.ZN (n_144_89), .A (n_142_89), .B (n_144_86), .C1 (n_140_88), .C2 (n_137_88) );
AOI211_X1 g_146_90 (.ZN (n_146_90), .A (n_143_87), .B (n_146_87), .C1 (n_142_87), .C2 (n_136_90) );
AOI211_X1 g_145_88 (.ZN (n_145_88), .A (n_144_89), .B (n_144_88), .C1 (n_144_86), .C2 (n_138_89) );
AOI211_X1 g_147_89 (.ZN (n_147_89), .A (n_146_90), .B (n_142_89), .C1 (n_146_87), .C2 (n_140_88) );
AOI211_X1 g_148_91 (.ZN (n_148_91), .A (n_145_88), .B (n_143_87), .C1 (n_144_88), .C2 (n_142_87) );
AOI211_X1 g_146_92 (.ZN (n_146_92), .A (n_147_89), .B (n_144_89), .C1 (n_142_89), .C2 (n_144_86) );
AOI211_X1 g_145_90 (.ZN (n_145_90), .A (n_148_91), .B (n_146_90), .C1 (n_143_87), .C2 (n_146_87) );
AOI211_X1 g_143_89 (.ZN (n_143_89), .A (n_146_92), .B (n_145_88), .C1 (n_144_89), .C2 (n_144_88) );
AOI211_X1 g_144_87 (.ZN (n_144_87), .A (n_145_90), .B (n_147_89), .C1 (n_146_90), .C2 (n_142_89) );
AOI211_X1 g_142_86 (.ZN (n_142_86), .A (n_143_89), .B (n_148_91), .C1 (n_145_88), .C2 (n_143_87) );
AOI211_X1 g_141_88 (.ZN (n_141_88), .A (n_144_87), .B (n_146_92), .C1 (n_147_89), .C2 (n_144_89) );
AOI211_X1 g_140_90 (.ZN (n_140_90), .A (n_142_86), .B (n_145_90), .C1 (n_148_91), .C2 (n_146_90) );
AOI211_X1 g_138_91 (.ZN (n_138_91), .A (n_141_88), .B (n_143_89), .C1 (n_146_92), .C2 (n_145_88) );
AOI211_X1 g_139_89 (.ZN (n_139_89), .A (n_140_90), .B (n_144_87), .C1 (n_145_90), .C2 (n_147_89) );
AOI211_X1 g_140_87 (.ZN (n_140_87), .A (n_138_91), .B (n_142_86), .C1 (n_143_89), .C2 (n_148_91) );
AOI211_X1 g_142_88 (.ZN (n_142_88), .A (n_139_89), .B (n_141_88), .C1 (n_144_87), .C2 (n_146_92) );
AOI211_X1 g_141_90 (.ZN (n_141_90), .A (n_140_87), .B (n_140_90), .C1 (n_142_86), .C2 (n_145_90) );
AOI211_X1 g_143_91 (.ZN (n_143_91), .A (n_142_88), .B (n_138_91), .C1 (n_141_88), .C2 (n_143_89) );
AOI211_X1 g_144_93 (.ZN (n_144_93), .A (n_141_90), .B (n_139_89), .C1 (n_140_90), .C2 (n_144_87) );
AOI211_X1 g_146_94 (.ZN (n_146_94), .A (n_143_91), .B (n_140_87), .C1 (n_138_91), .C2 (n_142_86) );
AOI211_X1 g_148_95 (.ZN (n_148_95), .A (n_144_93), .B (n_142_88), .C1 (n_139_89), .C2 (n_141_88) );
AOI211_X1 g_147_93 (.ZN (n_147_93), .A (n_146_94), .B (n_141_90), .C1 (n_140_87), .C2 (n_140_90) );
AOI211_X1 g_145_92 (.ZN (n_145_92), .A (n_148_95), .B (n_143_91), .C1 (n_142_88), .C2 (n_138_91) );
AOI211_X1 g_144_90 (.ZN (n_144_90), .A (n_147_93), .B (n_144_93), .C1 (n_141_90), .C2 (n_139_89) );
AOI211_X1 g_143_88 (.ZN (n_143_88), .A (n_145_92), .B (n_146_94), .C1 (n_143_91), .C2 (n_140_87) );
AOI211_X1 g_145_89 (.ZN (n_145_89), .A (n_144_90), .B (n_148_95), .C1 (n_144_93), .C2 (n_142_88) );
AOI211_X1 g_146_91 (.ZN (n_146_91), .A (n_143_88), .B (n_147_93), .C1 (n_146_94), .C2 (n_141_90) );
AOI211_X1 g_144_92 (.ZN (n_144_92), .A (n_145_89), .B (n_145_92), .C1 (n_148_95), .C2 (n_143_91) );
AOI211_X1 g_143_90 (.ZN (n_143_90), .A (n_146_91), .B (n_144_90), .C1 (n_147_93), .C2 (n_144_93) );
AOI211_X1 g_141_89 (.ZN (n_141_89), .A (n_144_92), .B (n_143_88), .C1 (n_145_92), .C2 (n_146_94) );
AOI211_X1 g_142_91 (.ZN (n_142_91), .A (n_143_90), .B (n_145_89), .C1 (n_144_90), .C2 (n_148_95) );
AOI211_X1 g_140_92 (.ZN (n_140_92), .A (n_141_89), .B (n_146_91), .C1 (n_143_88), .C2 (n_147_93) );
AOI211_X1 g_139_90 (.ZN (n_139_90), .A (n_142_91), .B (n_144_92), .C1 (n_145_89), .C2 (n_145_92) );
AOI211_X1 g_138_88 (.ZN (n_138_88), .A (n_140_92), .B (n_143_90), .C1 (n_146_91), .C2 (n_144_90) );
AOI211_X1 g_136_89 (.ZN (n_136_89), .A (n_139_90), .B (n_141_89), .C1 (n_144_92), .C2 (n_143_88) );
AOI211_X1 g_134_90 (.ZN (n_134_90), .A (n_138_88), .B (n_142_91), .C1 (n_143_90), .C2 (n_145_89) );
AOI211_X1 g_132_91 (.ZN (n_132_91), .A (n_136_89), .B (n_140_92), .C1 (n_141_89), .C2 (n_146_91) );
AOI211_X1 g_131_93 (.ZN (n_131_93), .A (n_134_90), .B (n_139_90), .C1 (n_142_91), .C2 (n_144_92) );
AOI211_X1 g_133_92 (.ZN (n_133_92), .A (n_132_91), .B (n_138_88), .C1 (n_140_92), .C2 (n_143_90) );
AOI211_X1 g_135_91 (.ZN (n_135_91), .A (n_131_93), .B (n_136_89), .C1 (n_139_90), .C2 (n_141_89) );
AOI211_X1 g_137_90 (.ZN (n_137_90), .A (n_133_92), .B (n_134_90), .C1 (n_138_88), .C2 (n_142_91) );
AOI211_X1 g_136_92 (.ZN (n_136_92), .A (n_135_91), .B (n_132_91), .C1 (n_136_89), .C2 (n_140_92) );
AOI211_X1 g_134_91 (.ZN (n_134_91), .A (n_137_90), .B (n_131_93), .C1 (n_134_90), .C2 (n_139_90) );
AOI211_X1 g_132_92 (.ZN (n_132_92), .A (n_136_92), .B (n_133_92), .C1 (n_132_91), .C2 (n_138_88) );
AOI211_X1 g_130_93 (.ZN (n_130_93), .A (n_134_91), .B (n_135_91), .C1 (n_131_93), .C2 (n_136_89) );
AOI211_X1 g_128_94 (.ZN (n_128_94), .A (n_132_92), .B (n_137_90), .C1 (n_133_92), .C2 (n_134_90) );
AOI211_X1 g_126_95 (.ZN (n_126_95), .A (n_130_93), .B (n_136_92), .C1 (n_135_91), .C2 (n_132_91) );
AOI211_X1 g_124_96 (.ZN (n_124_96), .A (n_128_94), .B (n_134_91), .C1 (n_137_90), .C2 (n_131_93) );
AOI211_X1 g_122_97 (.ZN (n_122_97), .A (n_126_95), .B (n_132_92), .C1 (n_136_92), .C2 (n_133_92) );
AOI211_X1 g_120_98 (.ZN (n_120_98), .A (n_124_96), .B (n_130_93), .C1 (n_134_91), .C2 (n_135_91) );
AOI211_X1 g_118_99 (.ZN (n_118_99), .A (n_122_97), .B (n_128_94), .C1 (n_132_92), .C2 (n_137_90) );
AOI211_X1 g_116_100 (.ZN (n_116_100), .A (n_120_98), .B (n_126_95), .C1 (n_130_93), .C2 (n_136_92) );
AOI211_X1 g_115_98 (.ZN (n_115_98), .A (n_118_99), .B (n_124_96), .C1 (n_128_94), .C2 (n_134_91) );
AOI211_X1 g_113_99 (.ZN (n_113_99), .A (n_116_100), .B (n_122_97), .C1 (n_126_95), .C2 (n_132_92) );
AOI211_X1 g_114_101 (.ZN (n_114_101), .A (n_115_98), .B (n_120_98), .C1 (n_124_96), .C2 (n_130_93) );
AOI211_X1 g_112_102 (.ZN (n_112_102), .A (n_113_99), .B (n_118_99), .C1 (n_122_97), .C2 (n_128_94) );
AOI211_X1 g_110_103 (.ZN (n_110_103), .A (n_114_101), .B (n_116_100), .C1 (n_120_98), .C2 (n_126_95) );
AOI211_X1 g_108_104 (.ZN (n_108_104), .A (n_112_102), .B (n_115_98), .C1 (n_118_99), .C2 (n_124_96) );
AOI211_X1 g_106_105 (.ZN (n_106_105), .A (n_110_103), .B (n_113_99), .C1 (n_116_100), .C2 (n_122_97) );
AOI211_X1 g_105_103 (.ZN (n_105_103), .A (n_108_104), .B (n_114_101), .C1 (n_115_98), .C2 (n_120_98) );
AOI211_X1 g_103_104 (.ZN (n_103_104), .A (n_106_105), .B (n_112_102), .C1 (n_113_99), .C2 (n_118_99) );
AOI211_X1 g_101_105 (.ZN (n_101_105), .A (n_105_103), .B (n_110_103), .C1 (n_114_101), .C2 (n_116_100) );
AOI211_X1 g_99_106 (.ZN (n_99_106), .A (n_103_104), .B (n_108_104), .C1 (n_112_102), .C2 (n_115_98) );
AOI211_X1 g_97_107 (.ZN (n_97_107), .A (n_101_105), .B (n_106_105), .C1 (n_110_103), .C2 (n_113_99) );
AOI211_X1 g_95_108 (.ZN (n_95_108), .A (n_99_106), .B (n_105_103), .C1 (n_108_104), .C2 (n_114_101) );
AOI211_X1 g_93_109 (.ZN (n_93_109), .A (n_97_107), .B (n_103_104), .C1 (n_106_105), .C2 (n_112_102) );
AOI211_X1 g_91_110 (.ZN (n_91_110), .A (n_95_108), .B (n_101_105), .C1 (n_105_103), .C2 (n_110_103) );
AOI211_X1 g_89_111 (.ZN (n_89_111), .A (n_93_109), .B (n_99_106), .C1 (n_103_104), .C2 (n_108_104) );
AOI211_X1 g_87_112 (.ZN (n_87_112), .A (n_91_110), .B (n_97_107), .C1 (n_101_105), .C2 (n_106_105) );
AOI211_X1 g_85_113 (.ZN (n_85_113), .A (n_89_111), .B (n_95_108), .C1 (n_99_106), .C2 (n_105_103) );
AOI211_X1 g_83_114 (.ZN (n_83_114), .A (n_87_112), .B (n_93_109), .C1 (n_97_107), .C2 (n_103_104) );
AOI211_X1 g_81_115 (.ZN (n_81_115), .A (n_85_113), .B (n_91_110), .C1 (n_95_108), .C2 (n_101_105) );
AOI211_X1 g_79_116 (.ZN (n_79_116), .A (n_83_114), .B (n_89_111), .C1 (n_93_109), .C2 (n_99_106) );
AOI211_X1 g_77_117 (.ZN (n_77_117), .A (n_81_115), .B (n_87_112), .C1 (n_91_110), .C2 (n_97_107) );
AOI211_X1 g_75_118 (.ZN (n_75_118), .A (n_79_116), .B (n_85_113), .C1 (n_89_111), .C2 (n_95_108) );
AOI211_X1 g_73_119 (.ZN (n_73_119), .A (n_77_117), .B (n_83_114), .C1 (n_87_112), .C2 (n_93_109) );
AOI211_X1 g_71_120 (.ZN (n_71_120), .A (n_75_118), .B (n_81_115), .C1 (n_85_113), .C2 (n_91_110) );
AOI211_X1 g_69_121 (.ZN (n_69_121), .A (n_73_119), .B (n_79_116), .C1 (n_83_114), .C2 (n_89_111) );
AOI211_X1 g_67_122 (.ZN (n_67_122), .A (n_71_120), .B (n_77_117), .C1 (n_81_115), .C2 (n_87_112) );
AOI211_X1 g_65_123 (.ZN (n_65_123), .A (n_69_121), .B (n_75_118), .C1 (n_79_116), .C2 (n_85_113) );
AOI211_X1 g_66_121 (.ZN (n_66_121), .A (n_67_122), .B (n_73_119), .C1 (n_77_117), .C2 (n_83_114) );
AOI211_X1 g_64_122 (.ZN (n_64_122), .A (n_65_123), .B (n_71_120), .C1 (n_75_118), .C2 (n_81_115) );
AOI211_X1 g_65_120 (.ZN (n_65_120), .A (n_66_121), .B (n_69_121), .C1 (n_73_119), .C2 (n_79_116) );
AOI211_X1 g_63_121 (.ZN (n_63_121), .A (n_64_122), .B (n_67_122), .C1 (n_71_120), .C2 (n_77_117) );
AOI211_X1 g_61_122 (.ZN (n_61_122), .A (n_65_120), .B (n_65_123), .C1 (n_69_121), .C2 (n_75_118) );
AOI211_X1 g_59_123 (.ZN (n_59_123), .A (n_63_121), .B (n_66_121), .C1 (n_67_122), .C2 (n_73_119) );
AOI211_X1 g_58_125 (.ZN (n_58_125), .A (n_61_122), .B (n_64_122), .C1 (n_65_123), .C2 (n_71_120) );
AOI211_X1 g_60_124 (.ZN (n_60_124), .A (n_59_123), .B (n_65_120), .C1 (n_66_121), .C2 (n_69_121) );
AOI211_X1 g_62_123 (.ZN (n_62_123), .A (n_58_125), .B (n_63_121), .C1 (n_64_122), .C2 (n_67_122) );
AOI211_X1 g_61_125 (.ZN (n_61_125), .A (n_60_124), .B (n_61_122), .C1 (n_65_120), .C2 (n_65_123) );
AOI211_X1 g_63_124 (.ZN (n_63_124), .A (n_62_123), .B (n_59_123), .C1 (n_63_121), .C2 (n_66_121) );
AOI211_X1 g_62_126 (.ZN (n_62_126), .A (n_61_125), .B (n_58_125), .C1 (n_61_122), .C2 (n_64_122) );
AOI211_X1 g_61_124 (.ZN (n_61_124), .A (n_63_124), .B (n_60_124), .C1 (n_59_123), .C2 (n_65_120) );
AOI211_X1 g_63_123 (.ZN (n_63_123), .A (n_62_126), .B (n_62_123), .C1 (n_58_125), .C2 (n_63_121) );
AOI211_X1 g_65_122 (.ZN (n_65_122), .A (n_61_124), .B (n_61_125), .C1 (n_60_124), .C2 (n_61_122) );
AOI211_X1 g_67_121 (.ZN (n_67_121), .A (n_63_123), .B (n_63_124), .C1 (n_62_123), .C2 (n_59_123) );
AOI211_X1 g_69_120 (.ZN (n_69_120), .A (n_65_122), .B (n_62_126), .C1 (n_61_125), .C2 (n_58_125) );
AOI211_X1 g_71_119 (.ZN (n_71_119), .A (n_67_121), .B (n_61_124), .C1 (n_63_124), .C2 (n_60_124) );
AOI211_X1 g_70_121 (.ZN (n_70_121), .A (n_69_120), .B (n_63_123), .C1 (n_62_126), .C2 (n_62_123) );
AOI211_X1 g_72_120 (.ZN (n_72_120), .A (n_71_119), .B (n_65_122), .C1 (n_61_124), .C2 (n_61_125) );
AOI211_X1 g_74_119 (.ZN (n_74_119), .A (n_70_121), .B (n_67_121), .C1 (n_63_123), .C2 (n_63_124) );
AOI211_X1 g_76_118 (.ZN (n_76_118), .A (n_72_120), .B (n_69_120), .C1 (n_65_122), .C2 (n_62_126) );
AOI211_X1 g_78_117 (.ZN (n_78_117), .A (n_74_119), .B (n_71_119), .C1 (n_67_121), .C2 (n_61_124) );
AOI211_X1 g_80_116 (.ZN (n_80_116), .A (n_76_118), .B (n_70_121), .C1 (n_69_120), .C2 (n_63_123) );
AOI211_X1 g_82_115 (.ZN (n_82_115), .A (n_78_117), .B (n_72_120), .C1 (n_71_119), .C2 (n_65_122) );
AOI211_X1 g_84_114 (.ZN (n_84_114), .A (n_80_116), .B (n_74_119), .C1 (n_70_121), .C2 (n_67_121) );
AOI211_X1 g_86_113 (.ZN (n_86_113), .A (n_82_115), .B (n_76_118), .C1 (n_72_120), .C2 (n_69_120) );
AOI211_X1 g_88_112 (.ZN (n_88_112), .A (n_84_114), .B (n_78_117), .C1 (n_74_119), .C2 (n_71_119) );
AOI211_X1 g_90_111 (.ZN (n_90_111), .A (n_86_113), .B (n_80_116), .C1 (n_76_118), .C2 (n_70_121) );
AOI211_X1 g_92_110 (.ZN (n_92_110), .A (n_88_112), .B (n_82_115), .C1 (n_78_117), .C2 (n_72_120) );
AOI211_X1 g_94_109 (.ZN (n_94_109), .A (n_90_111), .B (n_84_114), .C1 (n_80_116), .C2 (n_74_119) );
AOI211_X1 g_96_108 (.ZN (n_96_108), .A (n_92_110), .B (n_86_113), .C1 (n_82_115), .C2 (n_76_118) );
AOI211_X1 g_95_110 (.ZN (n_95_110), .A (n_94_109), .B (n_88_112), .C1 (n_84_114), .C2 (n_78_117) );
AOI211_X1 g_97_109 (.ZN (n_97_109), .A (n_96_108), .B (n_90_111), .C1 (n_86_113), .C2 (n_80_116) );
AOI211_X1 g_99_108 (.ZN (n_99_108), .A (n_95_110), .B (n_92_110), .C1 (n_88_112), .C2 (n_82_115) );
AOI211_X1 g_101_107 (.ZN (n_101_107), .A (n_97_109), .B (n_94_109), .C1 (n_90_111), .C2 (n_84_114) );
AOI211_X1 g_103_106 (.ZN (n_103_106), .A (n_99_108), .B (n_96_108), .C1 (n_92_110), .C2 (n_86_113) );
AOI211_X1 g_105_105 (.ZN (n_105_105), .A (n_101_107), .B (n_95_110), .C1 (n_94_109), .C2 (n_88_112) );
AOI211_X1 g_107_104 (.ZN (n_107_104), .A (n_103_106), .B (n_97_109), .C1 (n_96_108), .C2 (n_90_111) );
AOI211_X1 g_109_103 (.ZN (n_109_103), .A (n_105_105), .B (n_99_108), .C1 (n_95_110), .C2 (n_92_110) );
AOI211_X1 g_111_102 (.ZN (n_111_102), .A (n_107_104), .B (n_101_107), .C1 (n_97_109), .C2 (n_94_109) );
AOI211_X1 g_113_101 (.ZN (n_113_101), .A (n_109_103), .B (n_103_106), .C1 (n_99_108), .C2 (n_96_108) );
AOI211_X1 g_115_100 (.ZN (n_115_100), .A (n_111_102), .B (n_105_105), .C1 (n_101_107), .C2 (n_95_110) );
AOI211_X1 g_117_99 (.ZN (n_117_99), .A (n_113_101), .B (n_107_104), .C1 (n_103_106), .C2 (n_97_109) );
AOI211_X1 g_119_98 (.ZN (n_119_98), .A (n_115_100), .B (n_109_103), .C1 (n_105_105), .C2 (n_99_108) );
AOI211_X1 g_121_97 (.ZN (n_121_97), .A (n_117_99), .B (n_111_102), .C1 (n_107_104), .C2 (n_101_107) );
AOI211_X1 g_120_99 (.ZN (n_120_99), .A (n_119_98), .B (n_113_101), .C1 (n_109_103), .C2 (n_103_106) );
AOI211_X1 g_118_98 (.ZN (n_118_98), .A (n_121_97), .B (n_115_100), .C1 (n_111_102), .C2 (n_105_105) );
AOI211_X1 g_120_97 (.ZN (n_120_97), .A (n_120_99), .B (n_117_99), .C1 (n_113_101), .C2 (n_107_104) );
AOI211_X1 g_122_96 (.ZN (n_122_96), .A (n_118_98), .B (n_119_98), .C1 (n_115_100), .C2 (n_109_103) );
AOI211_X1 g_124_95 (.ZN (n_124_95), .A (n_120_97), .B (n_121_97), .C1 (n_117_99), .C2 (n_111_102) );
AOI211_X1 g_126_94 (.ZN (n_126_94), .A (n_122_96), .B (n_120_99), .C1 (n_119_98), .C2 (n_113_101) );
AOI211_X1 g_125_96 (.ZN (n_125_96), .A (n_124_95), .B (n_118_98), .C1 (n_121_97), .C2 (n_115_100) );
AOI211_X1 g_127_95 (.ZN (n_127_95), .A (n_126_94), .B (n_120_97), .C1 (n_120_99), .C2 (n_117_99) );
AOI211_X1 g_129_94 (.ZN (n_129_94), .A (n_125_96), .B (n_122_96), .C1 (n_118_98), .C2 (n_119_98) );
AOI211_X1 g_128_96 (.ZN (n_128_96), .A (n_127_95), .B (n_124_95), .C1 (n_120_97), .C2 (n_121_97) );
AOI211_X1 g_130_95 (.ZN (n_130_95), .A (n_129_94), .B (n_126_94), .C1 (n_122_96), .C2 (n_120_99) );
AOI211_X1 g_132_94 (.ZN (n_132_94), .A (n_128_96), .B (n_125_96), .C1 (n_124_95), .C2 (n_118_98) );
AOI211_X1 g_134_93 (.ZN (n_134_93), .A (n_130_95), .B (n_127_95), .C1 (n_126_94), .C2 (n_120_97) );
AOI211_X1 g_133_95 (.ZN (n_133_95), .A (n_132_94), .B (n_129_94), .C1 (n_125_96), .C2 (n_122_96) );
AOI211_X1 g_132_93 (.ZN (n_132_93), .A (n_134_93), .B (n_128_96), .C1 (n_127_95), .C2 (n_124_95) );
AOI211_X1 g_134_92 (.ZN (n_134_92), .A (n_133_95), .B (n_130_95), .C1 (n_129_94), .C2 (n_126_94) );
AOI211_X1 g_136_91 (.ZN (n_136_91), .A (n_132_93), .B (n_132_94), .C1 (n_128_96), .C2 (n_125_96) );
AOI211_X1 g_138_90 (.ZN (n_138_90), .A (n_134_92), .B (n_134_93), .C1 (n_130_95), .C2 (n_127_95) );
AOI211_X1 g_140_89 (.ZN (n_140_89), .A (n_136_91), .B (n_133_95), .C1 (n_132_94), .C2 (n_129_94) );
AOI211_X1 g_139_91 (.ZN (n_139_91), .A (n_138_90), .B (n_132_93), .C1 (n_134_93), .C2 (n_128_96) );
AOI211_X1 g_137_92 (.ZN (n_137_92), .A (n_140_89), .B (n_134_92), .C1 (n_133_95), .C2 (n_130_95) );
AOI211_X1 g_135_93 (.ZN (n_135_93), .A (n_139_91), .B (n_136_91), .C1 (n_132_93), .C2 (n_132_94) );
AOI211_X1 g_133_94 (.ZN (n_133_94), .A (n_137_92), .B (n_138_90), .C1 (n_134_92), .C2 (n_134_93) );
AOI211_X1 g_131_95 (.ZN (n_131_95), .A (n_135_93), .B (n_140_89), .C1 (n_136_91), .C2 (n_133_95) );
AOI211_X1 g_129_96 (.ZN (n_129_96), .A (n_133_94), .B (n_139_91), .C1 (n_138_90), .C2 (n_132_93) );
AOI211_X1 g_130_94 (.ZN (n_130_94), .A (n_131_95), .B (n_137_92), .C1 (n_140_89), .C2 (n_134_92) );
AOI211_X1 g_128_95 (.ZN (n_128_95), .A (n_129_96), .B (n_135_93), .C1 (n_139_91), .C2 (n_136_91) );
AOI211_X1 g_126_96 (.ZN (n_126_96), .A (n_130_94), .B (n_133_94), .C1 (n_137_92), .C2 (n_138_90) );
AOI211_X1 g_124_97 (.ZN (n_124_97), .A (n_128_95), .B (n_131_95), .C1 (n_135_93), .C2 (n_140_89) );
AOI211_X1 g_122_98 (.ZN (n_122_98), .A (n_126_96), .B (n_129_96), .C1 (n_133_94), .C2 (n_139_91) );
AOI211_X1 g_121_100 (.ZN (n_121_100), .A (n_124_97), .B (n_130_94), .C1 (n_131_95), .C2 (n_137_92) );
AOI211_X1 g_119_99 (.ZN (n_119_99), .A (n_122_98), .B (n_128_95), .C1 (n_129_96), .C2 (n_135_93) );
AOI211_X1 g_121_98 (.ZN (n_121_98), .A (n_121_100), .B (n_126_96), .C1 (n_130_94), .C2 (n_133_94) );
AOI211_X1 g_123_97 (.ZN (n_123_97), .A (n_119_99), .B (n_124_97), .C1 (n_128_95), .C2 (n_131_95) );
AOI211_X1 g_122_99 (.ZN (n_122_99), .A (n_121_98), .B (n_122_98), .C1 (n_126_96), .C2 (n_129_96) );
AOI211_X1 g_124_98 (.ZN (n_124_98), .A (n_123_97), .B (n_121_100), .C1 (n_124_97), .C2 (n_130_94) );
AOI211_X1 g_126_97 (.ZN (n_126_97), .A (n_122_99), .B (n_119_99), .C1 (n_122_98), .C2 (n_128_95) );
AOI211_X1 g_125_99 (.ZN (n_125_99), .A (n_124_98), .B (n_121_98), .C1 (n_121_100), .C2 (n_126_96) );
AOI211_X1 g_123_98 (.ZN (n_123_98), .A (n_126_97), .B (n_123_97), .C1 (n_119_99), .C2 (n_124_97) );
AOI211_X1 g_125_97 (.ZN (n_125_97), .A (n_125_99), .B (n_122_99), .C1 (n_121_98), .C2 (n_122_98) );
AOI211_X1 g_127_96 (.ZN (n_127_96), .A (n_123_98), .B (n_124_98), .C1 (n_123_97), .C2 (n_121_100) );
AOI211_X1 g_129_95 (.ZN (n_129_95), .A (n_125_97), .B (n_126_97), .C1 (n_122_99), .C2 (n_119_99) );
AOI211_X1 g_131_94 (.ZN (n_131_94), .A (n_127_96), .B (n_125_99), .C1 (n_124_98), .C2 (n_121_98) );
AOI211_X1 g_133_93 (.ZN (n_133_93), .A (n_129_95), .B (n_123_98), .C1 (n_126_97), .C2 (n_123_97) );
AOI211_X1 g_135_92 (.ZN (n_135_92), .A (n_131_94), .B (n_125_97), .C1 (n_125_99), .C2 (n_122_99) );
AOI211_X1 g_137_91 (.ZN (n_137_91), .A (n_133_93), .B (n_127_96), .C1 (n_123_98), .C2 (n_124_98) );
AOI211_X1 g_138_93 (.ZN (n_138_93), .A (n_135_92), .B (n_129_95), .C1 (n_125_97), .C2 (n_126_97) );
AOI211_X1 g_136_94 (.ZN (n_136_94), .A (n_137_91), .B (n_131_94), .C1 (n_127_96), .C2 (n_125_99) );
AOI211_X1 g_134_95 (.ZN (n_134_95), .A (n_138_93), .B (n_133_93), .C1 (n_129_95), .C2 (n_123_98) );
AOI211_X1 g_132_96 (.ZN (n_132_96), .A (n_136_94), .B (n_135_92), .C1 (n_131_94), .C2 (n_125_97) );
AOI211_X1 g_130_97 (.ZN (n_130_97), .A (n_134_95), .B (n_137_91), .C1 (n_133_93), .C2 (n_127_96) );
AOI211_X1 g_128_98 (.ZN (n_128_98), .A (n_132_96), .B (n_138_93), .C1 (n_135_92), .C2 (n_129_95) );
AOI211_X1 g_126_99 (.ZN (n_126_99), .A (n_130_97), .B (n_136_94), .C1 (n_137_91), .C2 (n_131_94) );
AOI211_X1 g_127_97 (.ZN (n_127_97), .A (n_128_98), .B (n_134_95), .C1 (n_138_93), .C2 (n_133_93) );
AOI211_X1 g_125_98 (.ZN (n_125_98), .A (n_126_99), .B (n_132_96), .C1 (n_136_94), .C2 (n_135_92) );
AOI211_X1 g_123_99 (.ZN (n_123_99), .A (n_127_97), .B (n_130_97), .C1 (n_134_95), .C2 (n_137_91) );
AOI211_X1 g_124_101 (.ZN (n_124_101), .A (n_125_98), .B (n_128_98), .C1 (n_132_96), .C2 (n_138_93) );
AOI211_X1 g_122_100 (.ZN (n_122_100), .A (n_123_99), .B (n_126_99), .C1 (n_130_97), .C2 (n_136_94) );
AOI211_X1 g_124_99 (.ZN (n_124_99), .A (n_124_101), .B (n_127_97), .C1 (n_128_98), .C2 (n_134_95) );
AOI211_X1 g_126_98 (.ZN (n_126_98), .A (n_122_100), .B (n_125_98), .C1 (n_126_99), .C2 (n_132_96) );
AOI211_X1 g_128_97 (.ZN (n_128_97), .A (n_124_99), .B (n_123_99), .C1 (n_127_97), .C2 (n_130_97) );
AOI211_X1 g_130_96 (.ZN (n_130_96), .A (n_126_98), .B (n_124_101), .C1 (n_125_98), .C2 (n_128_98) );
AOI211_X1 g_132_95 (.ZN (n_132_95), .A (n_128_97), .B (n_122_100), .C1 (n_123_99), .C2 (n_126_99) );
AOI211_X1 g_134_94 (.ZN (n_134_94), .A (n_130_96), .B (n_124_99), .C1 (n_124_101), .C2 (n_127_97) );
AOI211_X1 g_136_93 (.ZN (n_136_93), .A (n_132_95), .B (n_126_98), .C1 (n_122_100), .C2 (n_125_98) );
AOI211_X1 g_138_92 (.ZN (n_138_92), .A (n_134_94), .B (n_128_97), .C1 (n_124_99), .C2 (n_123_99) );
AOI211_X1 g_140_91 (.ZN (n_140_91), .A (n_136_93), .B (n_130_96), .C1 (n_126_98), .C2 (n_124_101) );
AOI211_X1 g_142_90 (.ZN (n_142_90), .A (n_138_92), .B (n_132_95), .C1 (n_128_97), .C2 (n_122_100) );
AOI211_X1 g_144_91 (.ZN (n_144_91), .A (n_140_91), .B (n_134_94), .C1 (n_130_96), .C2 (n_124_99) );
AOI211_X1 g_142_92 (.ZN (n_142_92), .A (n_142_90), .B (n_136_93), .C1 (n_132_95), .C2 (n_126_98) );
AOI211_X1 g_140_93 (.ZN (n_140_93), .A (n_144_91), .B (n_138_92), .C1 (n_134_94), .C2 (n_128_97) );
AOI211_X1 g_141_91 (.ZN (n_141_91), .A (n_142_92), .B (n_140_91), .C1 (n_136_93), .C2 (n_130_96) );
AOI211_X1 g_139_92 (.ZN (n_139_92), .A (n_140_93), .B (n_142_90), .C1 (n_138_92), .C2 (n_132_95) );
AOI211_X1 g_137_93 (.ZN (n_137_93), .A (n_141_91), .B (n_144_91), .C1 (n_140_91), .C2 (n_134_94) );
AOI211_X1 g_135_94 (.ZN (n_135_94), .A (n_139_92), .B (n_142_92), .C1 (n_142_90), .C2 (n_136_93) );
AOI211_X1 g_134_96 (.ZN (n_134_96), .A (n_137_93), .B (n_140_93), .C1 (n_144_91), .C2 (n_138_92) );
AOI211_X1 g_136_95 (.ZN (n_136_95), .A (n_135_94), .B (n_141_91), .C1 (n_142_92), .C2 (n_140_91) );
AOI211_X1 g_138_94 (.ZN (n_138_94), .A (n_134_96), .B (n_139_92), .C1 (n_140_93), .C2 (n_142_90) );
AOI211_X1 g_137_96 (.ZN (n_137_96), .A (n_136_95), .B (n_137_93), .C1 (n_141_91), .C2 (n_144_91) );
AOI211_X1 g_135_95 (.ZN (n_135_95), .A (n_138_94), .B (n_135_94), .C1 (n_139_92), .C2 (n_142_92) );
AOI211_X1 g_137_94 (.ZN (n_137_94), .A (n_137_96), .B (n_134_96), .C1 (n_137_93), .C2 (n_140_93) );
AOI211_X1 g_139_93 (.ZN (n_139_93), .A (n_135_95), .B (n_136_95), .C1 (n_135_94), .C2 (n_141_91) );
AOI211_X1 g_141_92 (.ZN (n_141_92), .A (n_137_94), .B (n_138_94), .C1 (n_134_96), .C2 (n_139_92) );
AOI211_X1 g_143_93 (.ZN (n_143_93), .A (n_139_93), .B (n_137_96), .C1 (n_136_95), .C2 (n_137_93) );
AOI211_X1 g_145_94 (.ZN (n_145_94), .A (n_141_92), .B (n_135_95), .C1 (n_138_94), .C2 (n_135_94) );
AOI211_X1 g_146_96 (.ZN (n_146_96), .A (n_143_93), .B (n_137_94), .C1 (n_137_96), .C2 (n_134_96) );
AOI211_X1 g_144_95 (.ZN (n_144_95), .A (n_145_94), .B (n_139_93), .C1 (n_135_95), .C2 (n_136_95) );
AOI211_X1 g_145_93 (.ZN (n_145_93), .A (n_146_96), .B (n_141_92), .C1 (n_137_94), .C2 (n_138_94) );
AOI211_X1 g_143_92 (.ZN (n_143_92), .A (n_144_95), .B (n_143_93), .C1 (n_139_93), .C2 (n_137_96) );
AOI211_X1 g_142_94 (.ZN (n_142_94), .A (n_145_93), .B (n_145_94), .C1 (n_141_92), .C2 (n_135_95) );
AOI211_X1 g_140_95 (.ZN (n_140_95), .A (n_143_92), .B (n_146_96), .C1 (n_143_93), .C2 (n_137_94) );
AOI211_X1 g_141_93 (.ZN (n_141_93), .A (n_142_94), .B (n_144_95), .C1 (n_145_94), .C2 (n_139_93) );
AOI211_X1 g_143_94 (.ZN (n_143_94), .A (n_140_95), .B (n_145_93), .C1 (n_146_96), .C2 (n_141_92) );
AOI211_X1 g_142_96 (.ZN (n_142_96), .A (n_141_93), .B (n_143_92), .C1 (n_144_95), .C2 (n_143_93) );
AOI211_X1 g_141_94 (.ZN (n_141_94), .A (n_143_94), .B (n_142_94), .C1 (n_145_93), .C2 (n_145_94) );
AOI211_X1 g_139_95 (.ZN (n_139_95), .A (n_142_96), .B (n_140_95), .C1 (n_143_92), .C2 (n_146_96) );
AOI211_X1 g_140_97 (.ZN (n_140_97), .A (n_141_94), .B (n_141_93), .C1 (n_142_94), .C2 (n_144_95) );
AOI211_X1 g_138_96 (.ZN (n_138_96), .A (n_139_95), .B (n_143_94), .C1 (n_140_95), .C2 (n_145_93) );
AOI211_X1 g_139_94 (.ZN (n_139_94), .A (n_140_97), .B (n_142_96), .C1 (n_141_93), .C2 (n_143_92) );
AOI211_X1 g_137_95 (.ZN (n_137_95), .A (n_138_96), .B (n_141_94), .C1 (n_143_94), .C2 (n_142_94) );
AOI211_X1 g_135_96 (.ZN (n_135_96), .A (n_139_94), .B (n_139_95), .C1 (n_142_96), .C2 (n_140_95) );
AOI211_X1 g_133_97 (.ZN (n_133_97), .A (n_137_95), .B (n_140_97), .C1 (n_141_94), .C2 (n_141_93) );
AOI211_X1 g_131_96 (.ZN (n_131_96), .A (n_135_96), .B (n_138_96), .C1 (n_139_95), .C2 (n_143_94) );
AOI211_X1 g_129_97 (.ZN (n_129_97), .A (n_133_97), .B (n_139_94), .C1 (n_140_97), .C2 (n_142_96) );
AOI211_X1 g_127_98 (.ZN (n_127_98), .A (n_131_96), .B (n_137_95), .C1 (n_138_96), .C2 (n_141_94) );
AOI211_X1 g_126_100 (.ZN (n_126_100), .A (n_129_97), .B (n_135_96), .C1 (n_139_94), .C2 (n_139_95) );
AOI211_X1 g_128_99 (.ZN (n_128_99), .A (n_127_98), .B (n_133_97), .C1 (n_137_95), .C2 (n_140_97) );
AOI211_X1 g_130_98 (.ZN (n_130_98), .A (n_126_100), .B (n_131_96), .C1 (n_135_96), .C2 (n_138_96) );
AOI211_X1 g_132_97 (.ZN (n_132_97), .A (n_128_99), .B (n_129_97), .C1 (n_133_97), .C2 (n_139_94) );
AOI211_X1 g_131_99 (.ZN (n_131_99), .A (n_130_98), .B (n_127_98), .C1 (n_131_96), .C2 (n_137_95) );
AOI211_X1 g_129_98 (.ZN (n_129_98), .A (n_132_97), .B (n_126_100), .C1 (n_129_97), .C2 (n_135_96) );
AOI211_X1 g_131_97 (.ZN (n_131_97), .A (n_131_99), .B (n_128_99), .C1 (n_127_98), .C2 (n_133_97) );
AOI211_X1 g_133_96 (.ZN (n_133_96), .A (n_129_98), .B (n_130_98), .C1 (n_126_100), .C2 (n_131_96) );
AOI211_X1 g_135_97 (.ZN (n_135_97), .A (n_131_97), .B (n_132_97), .C1 (n_128_99), .C2 (n_129_97) );
AOI211_X1 g_133_98 (.ZN (n_133_98), .A (n_133_96), .B (n_131_99), .C1 (n_130_98), .C2 (n_127_98) );
AOI211_X1 g_132_100 (.ZN (n_132_100), .A (n_135_97), .B (n_129_98), .C1 (n_132_97), .C2 (n_126_100) );
AOI211_X1 g_131_98 (.ZN (n_131_98), .A (n_133_98), .B (n_131_97), .C1 (n_131_99), .C2 (n_128_99) );
AOI211_X1 g_129_99 (.ZN (n_129_99), .A (n_132_100), .B (n_133_96), .C1 (n_129_98), .C2 (n_130_98) );
AOI211_X1 g_127_100 (.ZN (n_127_100), .A (n_131_98), .B (n_135_97), .C1 (n_131_97), .C2 (n_132_97) );
AOI211_X1 g_125_101 (.ZN (n_125_101), .A (n_129_99), .B (n_133_98), .C1 (n_133_96), .C2 (n_131_99) );
AOI211_X1 g_123_100 (.ZN (n_123_100), .A (n_127_100), .B (n_132_100), .C1 (n_135_97), .C2 (n_129_98) );
AOI211_X1 g_121_99 (.ZN (n_121_99), .A (n_125_101), .B (n_131_98), .C1 (n_133_98), .C2 (n_131_97) );
AOI211_X1 g_119_100 (.ZN (n_119_100), .A (n_123_100), .B (n_129_99), .C1 (n_132_100), .C2 (n_133_96) );
AOI211_X1 g_121_101 (.ZN (n_121_101), .A (n_121_99), .B (n_127_100), .C1 (n_131_98), .C2 (n_135_97) );
AOI211_X1 g_123_102 (.ZN (n_123_102), .A (n_119_100), .B (n_125_101), .C1 (n_129_99), .C2 (n_133_98) );
AOI211_X1 g_124_100 (.ZN (n_124_100), .A (n_121_101), .B (n_123_100), .C1 (n_127_100), .C2 (n_132_100) );
AOI211_X1 g_122_101 (.ZN (n_122_101), .A (n_123_102), .B (n_121_99), .C1 (n_125_101), .C2 (n_131_98) );
AOI211_X1 g_120_100 (.ZN (n_120_100), .A (n_124_100), .B (n_119_100), .C1 (n_123_100), .C2 (n_129_99) );
AOI211_X1 g_118_101 (.ZN (n_118_101), .A (n_122_101), .B (n_121_101), .C1 (n_121_99), .C2 (n_127_100) );
AOI211_X1 g_120_102 (.ZN (n_120_102), .A (n_120_100), .B (n_123_102), .C1 (n_119_100), .C2 (n_125_101) );
AOI211_X1 g_122_103 (.ZN (n_122_103), .A (n_118_101), .B (n_124_100), .C1 (n_121_101), .C2 (n_123_100) );
AOI211_X1 g_123_101 (.ZN (n_123_101), .A (n_120_102), .B (n_122_101), .C1 (n_123_102), .C2 (n_121_99) );
AOI211_X1 g_125_100 (.ZN (n_125_100), .A (n_122_103), .B (n_120_100), .C1 (n_124_100), .C2 (n_119_100) );
AOI211_X1 g_127_99 (.ZN (n_127_99), .A (n_123_101), .B (n_118_101), .C1 (n_122_101), .C2 (n_121_101) );
AOI211_X1 g_129_100 (.ZN (n_129_100), .A (n_125_100), .B (n_120_102), .C1 (n_120_100), .C2 (n_123_102) );
AOI211_X1 g_127_101 (.ZN (n_127_101), .A (n_127_99), .B (n_122_103), .C1 (n_118_101), .C2 (n_124_100) );
AOI211_X1 g_125_102 (.ZN (n_125_102), .A (n_129_100), .B (n_123_101), .C1 (n_120_102), .C2 (n_122_101) );
AOI211_X1 g_123_103 (.ZN (n_123_103), .A (n_127_101), .B (n_125_100), .C1 (n_122_103), .C2 (n_120_100) );
AOI211_X1 g_121_102 (.ZN (n_121_102), .A (n_125_102), .B (n_127_99), .C1 (n_123_101), .C2 (n_118_101) );
AOI211_X1 g_119_101 (.ZN (n_119_101), .A (n_123_103), .B (n_129_100), .C1 (n_125_100), .C2 (n_120_102) );
AOI211_X1 g_117_100 (.ZN (n_117_100), .A (n_121_102), .B (n_127_101), .C1 (n_127_99), .C2 (n_122_103) );
AOI211_X1 g_116_102 (.ZN (n_116_102), .A (n_119_101), .B (n_125_102), .C1 (n_129_100), .C2 (n_123_101) );
AOI211_X1 g_114_103 (.ZN (n_114_103), .A (n_117_100), .B (n_123_103), .C1 (n_127_101), .C2 (n_125_100) );
AOI211_X1 g_115_101 (.ZN (n_115_101), .A (n_116_102), .B (n_121_102), .C1 (n_125_102), .C2 (n_127_99) );
AOI211_X1 g_116_99 (.ZN (n_116_99), .A (n_114_103), .B (n_119_101), .C1 (n_123_103), .C2 (n_129_100) );
AOI211_X1 g_114_100 (.ZN (n_114_100), .A (n_115_101), .B (n_117_100), .C1 (n_121_102), .C2 (n_127_101) );
AOI211_X1 g_112_101 (.ZN (n_112_101), .A (n_116_99), .B (n_116_102), .C1 (n_119_101), .C2 (n_125_102) );
AOI211_X1 g_110_102 (.ZN (n_110_102), .A (n_114_100), .B (n_114_103), .C1 (n_117_100), .C2 (n_123_103) );
AOI211_X1 g_108_103 (.ZN (n_108_103), .A (n_112_101), .B (n_115_101), .C1 (n_116_102), .C2 (n_121_102) );
AOI211_X1 g_106_104 (.ZN (n_106_104), .A (n_110_102), .B (n_116_99), .C1 (n_114_103), .C2 (n_119_101) );
AOI211_X1 g_104_105 (.ZN (n_104_105), .A (n_108_103), .B (n_114_100), .C1 (n_115_101), .C2 (n_117_100) );
AOI211_X1 g_102_106 (.ZN (n_102_106), .A (n_106_104), .B (n_112_101), .C1 (n_116_99), .C2 (n_116_102) );
AOI211_X1 g_100_107 (.ZN (n_100_107), .A (n_104_105), .B (n_110_102), .C1 (n_114_100), .C2 (n_114_103) );
AOI211_X1 g_98_108 (.ZN (n_98_108), .A (n_102_106), .B (n_108_103), .C1 (n_112_101), .C2 (n_115_101) );
AOI211_X1 g_96_109 (.ZN (n_96_109), .A (n_100_107), .B (n_106_104), .C1 (n_110_102), .C2 (n_116_99) );
AOI211_X1 g_94_110 (.ZN (n_94_110), .A (n_98_108), .B (n_104_105), .C1 (n_108_103), .C2 (n_114_100) );
AOI211_X1 g_92_111 (.ZN (n_92_111), .A (n_96_109), .B (n_102_106), .C1 (n_106_104), .C2 (n_112_101) );
AOI211_X1 g_90_112 (.ZN (n_90_112), .A (n_94_110), .B (n_100_107), .C1 (n_104_105), .C2 (n_110_102) );
AOI211_X1 g_88_113 (.ZN (n_88_113), .A (n_92_111), .B (n_98_108), .C1 (n_102_106), .C2 (n_108_103) );
AOI211_X1 g_86_114 (.ZN (n_86_114), .A (n_90_112), .B (n_96_109), .C1 (n_100_107), .C2 (n_106_104) );
AOI211_X1 g_84_115 (.ZN (n_84_115), .A (n_88_113), .B (n_94_110), .C1 (n_98_108), .C2 (n_104_105) );
AOI211_X1 g_82_116 (.ZN (n_82_116), .A (n_86_114), .B (n_92_111), .C1 (n_96_109), .C2 (n_102_106) );
AOI211_X1 g_80_115 (.ZN (n_80_115), .A (n_84_115), .B (n_90_112), .C1 (n_94_110), .C2 (n_100_107) );
AOI211_X1 g_78_116 (.ZN (n_78_116), .A (n_82_116), .B (n_88_113), .C1 (n_92_111), .C2 (n_98_108) );
AOI211_X1 g_76_117 (.ZN (n_76_117), .A (n_80_115), .B (n_86_114), .C1 (n_90_112), .C2 (n_96_109) );
AOI211_X1 g_74_118 (.ZN (n_74_118), .A (n_78_116), .B (n_84_115), .C1 (n_88_113), .C2 (n_94_110) );
AOI211_X1 g_72_119 (.ZN (n_72_119), .A (n_76_117), .B (n_82_116), .C1 (n_86_114), .C2 (n_92_111) );
AOI211_X1 g_70_120 (.ZN (n_70_120), .A (n_74_118), .B (n_80_115), .C1 (n_84_115), .C2 (n_90_112) );
AOI211_X1 g_68_121 (.ZN (n_68_121), .A (n_72_119), .B (n_78_116), .C1 (n_82_116), .C2 (n_88_113) );
AOI211_X1 g_66_122 (.ZN (n_66_122), .A (n_70_120), .B (n_76_117), .C1 (n_80_115), .C2 (n_86_114) );
AOI211_X1 g_64_123 (.ZN (n_64_123), .A (n_68_121), .B (n_74_118), .C1 (n_78_116), .C2 (n_84_115) );
AOI211_X1 g_62_124 (.ZN (n_62_124), .A (n_66_122), .B (n_72_119), .C1 (n_76_117), .C2 (n_82_116) );
AOI211_X1 g_60_125 (.ZN (n_60_125), .A (n_64_123), .B (n_70_120), .C1 (n_74_118), .C2 (n_80_115) );
AOI211_X1 g_58_126 (.ZN (n_58_126), .A (n_62_124), .B (n_68_121), .C1 (n_72_119), .C2 (n_78_116) );
AOI211_X1 g_56_127 (.ZN (n_56_127), .A (n_60_125), .B (n_66_122), .C1 (n_70_120), .C2 (n_76_117) );
AOI211_X1 g_57_125 (.ZN (n_57_125), .A (n_58_126), .B (n_64_123), .C1 (n_68_121), .C2 (n_74_118) );
AOI211_X1 g_55_126 (.ZN (n_55_126), .A (n_56_127), .B (n_62_124), .C1 (n_66_122), .C2 (n_72_119) );
AOI211_X1 g_53_127 (.ZN (n_53_127), .A (n_57_125), .B (n_60_125), .C1 (n_64_123), .C2 (n_70_120) );
AOI211_X1 g_51_128 (.ZN (n_51_128), .A (n_55_126), .B (n_58_126), .C1 (n_62_124), .C2 (n_68_121) );
AOI211_X1 g_50_130 (.ZN (n_50_130), .A (n_53_127), .B (n_56_127), .C1 (n_60_125), .C2 (n_66_122) );
AOI211_X1 g_52_129 (.ZN (n_52_129), .A (n_51_128), .B (n_57_125), .C1 (n_58_126), .C2 (n_64_123) );
AOI211_X1 g_54_128 (.ZN (n_54_128), .A (n_50_130), .B (n_55_126), .C1 (n_56_127), .C2 (n_62_124) );
AOI211_X1 g_53_130 (.ZN (n_53_130), .A (n_52_129), .B (n_53_127), .C1 (n_57_125), .C2 (n_60_125) );
AOI211_X1 g_52_128 (.ZN (n_52_128), .A (n_54_128), .B (n_51_128), .C1 (n_55_126), .C2 (n_58_126) );
AOI211_X1 g_54_127 (.ZN (n_54_127), .A (n_53_130), .B (n_50_130), .C1 (n_53_127), .C2 (n_56_127) );
AOI211_X1 g_56_126 (.ZN (n_56_126), .A (n_52_128), .B (n_52_129), .C1 (n_51_128), .C2 (n_57_125) );
AOI211_X1 g_55_128 (.ZN (n_55_128), .A (n_54_127), .B (n_54_128), .C1 (n_50_130), .C2 (n_55_126) );
AOI211_X1 g_57_127 (.ZN (n_57_127), .A (n_56_126), .B (n_53_130), .C1 (n_52_129), .C2 (n_53_127) );
AOI211_X1 g_59_126 (.ZN (n_59_126), .A (n_55_128), .B (n_52_128), .C1 (n_54_128), .C2 (n_51_128) );
AOI211_X1 g_58_128 (.ZN (n_58_128), .A (n_57_127), .B (n_54_127), .C1 (n_53_130), .C2 (n_50_130) );
AOI211_X1 g_60_127 (.ZN (n_60_127), .A (n_59_126), .B (n_56_126), .C1 (n_52_128), .C2 (n_52_129) );
AOI211_X1 g_59_125 (.ZN (n_59_125), .A (n_58_128), .B (n_55_128), .C1 (n_54_127), .C2 (n_54_128) );
AOI211_X1 g_57_126 (.ZN (n_57_126), .A (n_60_127), .B (n_57_127), .C1 (n_56_126), .C2 (n_53_130) );
AOI211_X1 g_55_127 (.ZN (n_55_127), .A (n_59_125), .B (n_59_126), .C1 (n_55_128), .C2 (n_52_128) );
AOI211_X1 g_53_128 (.ZN (n_53_128), .A (n_57_126), .B (n_58_128), .C1 (n_57_127), .C2 (n_54_127) );
AOI211_X1 g_51_129 (.ZN (n_51_129), .A (n_55_127), .B (n_60_127), .C1 (n_59_126), .C2 (n_56_126) );
AOI211_X1 g_49_130 (.ZN (n_49_130), .A (n_53_128), .B (n_59_125), .C1 (n_58_128), .C2 (n_55_128) );
AOI211_X1 g_47_131 (.ZN (n_47_131), .A (n_51_129), .B (n_57_126), .C1 (n_60_127), .C2 (n_57_127) );
AOI211_X1 g_45_132 (.ZN (n_45_132), .A (n_49_130), .B (n_55_127), .C1 (n_59_125), .C2 (n_59_126) );
AOI211_X1 g_43_133 (.ZN (n_43_133), .A (n_47_131), .B (n_53_128), .C1 (n_57_126), .C2 (n_58_128) );
AOI211_X1 g_41_134 (.ZN (n_41_134), .A (n_45_132), .B (n_51_129), .C1 (n_55_127), .C2 (n_60_127) );
AOI211_X1 g_39_135 (.ZN (n_39_135), .A (n_43_133), .B (n_49_130), .C1 (n_53_128), .C2 (n_59_125) );
AOI211_X1 g_37_136 (.ZN (n_37_136), .A (n_41_134), .B (n_47_131), .C1 (n_51_129), .C2 (n_57_126) );
AOI211_X1 g_36_134 (.ZN (n_36_134), .A (n_39_135), .B (n_45_132), .C1 (n_49_130), .C2 (n_55_127) );
AOI211_X1 g_34_135 (.ZN (n_34_135), .A (n_37_136), .B (n_43_133), .C1 (n_47_131), .C2 (n_53_128) );
AOI211_X1 g_32_136 (.ZN (n_32_136), .A (n_36_134), .B (n_41_134), .C1 (n_45_132), .C2 (n_51_129) );
AOI211_X1 g_30_137 (.ZN (n_30_137), .A (n_34_135), .B (n_39_135), .C1 (n_43_133), .C2 (n_49_130) );
AOI211_X1 g_28_138 (.ZN (n_28_138), .A (n_32_136), .B (n_37_136), .C1 (n_41_134), .C2 (n_47_131) );
AOI211_X1 g_26_139 (.ZN (n_26_139), .A (n_30_137), .B (n_36_134), .C1 (n_39_135), .C2 (n_45_132) );
AOI211_X1 g_24_140 (.ZN (n_24_140), .A (n_28_138), .B (n_34_135), .C1 (n_37_136), .C2 (n_43_133) );
AOI211_X1 g_22_141 (.ZN (n_22_141), .A (n_26_139), .B (n_32_136), .C1 (n_36_134), .C2 (n_41_134) );
AOI211_X1 g_21_143 (.ZN (n_21_143), .A (n_24_140), .B (n_30_137), .C1 (n_34_135), .C2 (n_39_135) );
AOI211_X1 g_23_142 (.ZN (n_23_142), .A (n_22_141), .B (n_28_138), .C1 (n_32_136), .C2 (n_37_136) );
AOI211_X1 g_25_141 (.ZN (n_25_141), .A (n_21_143), .B (n_26_139), .C1 (n_30_137), .C2 (n_36_134) );
AOI211_X1 g_27_140 (.ZN (n_27_140), .A (n_23_142), .B (n_24_140), .C1 (n_28_138), .C2 (n_34_135) );
AOI211_X1 g_29_139 (.ZN (n_29_139), .A (n_25_141), .B (n_22_141), .C1 (n_26_139), .C2 (n_32_136) );
AOI211_X1 g_31_138 (.ZN (n_31_138), .A (n_27_140), .B (n_21_143), .C1 (n_24_140), .C2 (n_30_137) );
AOI211_X1 g_33_137 (.ZN (n_33_137), .A (n_29_139), .B (n_23_142), .C1 (n_22_141), .C2 (n_28_138) );
AOI211_X1 g_35_136 (.ZN (n_35_136), .A (n_31_138), .B (n_25_141), .C1 (n_21_143), .C2 (n_26_139) );
AOI211_X1 g_37_135 (.ZN (n_37_135), .A (n_33_137), .B (n_27_140), .C1 (n_23_142), .C2 (n_24_140) );
AOI211_X1 g_39_134 (.ZN (n_39_134), .A (n_35_136), .B (n_29_139), .C1 (n_25_141), .C2 (n_22_141) );
AOI211_X1 g_41_133 (.ZN (n_41_133), .A (n_37_135), .B (n_31_138), .C1 (n_27_140), .C2 (n_21_143) );
AOI211_X1 g_43_132 (.ZN (n_43_132), .A (n_39_134), .B (n_33_137), .C1 (n_29_139), .C2 (n_23_142) );
AOI211_X1 g_42_134 (.ZN (n_42_134), .A (n_41_133), .B (n_35_136), .C1 (n_31_138), .C2 (n_25_141) );
AOI211_X1 g_44_133 (.ZN (n_44_133), .A (n_43_132), .B (n_37_135), .C1 (n_33_137), .C2 (n_27_140) );
AOI211_X1 g_46_132 (.ZN (n_46_132), .A (n_42_134), .B (n_39_134), .C1 (n_35_136), .C2 (n_29_139) );
AOI211_X1 g_48_131 (.ZN (n_48_131), .A (n_44_133), .B (n_41_133), .C1 (n_37_135), .C2 (n_31_138) );
AOI211_X1 g_47_133 (.ZN (n_47_133), .A (n_46_132), .B (n_43_132), .C1 (n_39_134), .C2 (n_33_137) );
AOI211_X1 g_46_131 (.ZN (n_46_131), .A (n_48_131), .B (n_42_134), .C1 (n_41_133), .C2 (n_35_136) );
AOI211_X1 g_44_132 (.ZN (n_44_132), .A (n_47_133), .B (n_44_133), .C1 (n_43_132), .C2 (n_37_135) );
AOI211_X1 g_45_134 (.ZN (n_45_134), .A (n_46_131), .B (n_46_132), .C1 (n_42_134), .C2 (n_39_134) );
AOI211_X1 g_43_135 (.ZN (n_43_135), .A (n_44_132), .B (n_48_131), .C1 (n_44_133), .C2 (n_41_133) );
AOI211_X1 g_41_136 (.ZN (n_41_136), .A (n_45_134), .B (n_47_133), .C1 (n_46_132), .C2 (n_43_132) );
AOI211_X1 g_39_137 (.ZN (n_39_137), .A (n_43_135), .B (n_46_131), .C1 (n_48_131), .C2 (n_42_134) );
AOI211_X1 g_40_135 (.ZN (n_40_135), .A (n_41_136), .B (n_44_132), .C1 (n_47_133), .C2 (n_44_133) );
AOI211_X1 g_38_136 (.ZN (n_38_136), .A (n_39_137), .B (n_45_134), .C1 (n_46_131), .C2 (n_46_132) );
AOI211_X1 g_36_135 (.ZN (n_36_135), .A (n_40_135), .B (n_43_135), .C1 (n_44_132), .C2 (n_48_131) );
AOI211_X1 g_34_136 (.ZN (n_34_136), .A (n_38_136), .B (n_41_136), .C1 (n_45_134), .C2 (n_47_133) );
AOI211_X1 g_32_137 (.ZN (n_32_137), .A (n_36_135), .B (n_39_137), .C1 (n_43_135), .C2 (n_46_131) );
AOI211_X1 g_30_138 (.ZN (n_30_138), .A (n_34_136), .B (n_40_135), .C1 (n_41_136), .C2 (n_44_132) );
AOI211_X1 g_28_139 (.ZN (n_28_139), .A (n_32_137), .B (n_38_136), .C1 (n_39_137), .C2 (n_45_134) );
AOI211_X1 g_26_140 (.ZN (n_26_140), .A (n_30_138), .B (n_36_135), .C1 (n_40_135), .C2 (n_43_135) );
AOI211_X1 g_24_141 (.ZN (n_24_141), .A (n_28_139), .B (n_34_136), .C1 (n_38_136), .C2 (n_41_136) );
AOI211_X1 g_22_142 (.ZN (n_22_142), .A (n_26_140), .B (n_32_137), .C1 (n_36_135), .C2 (n_39_137) );
AOI211_X1 g_21_144 (.ZN (n_21_144), .A (n_24_141), .B (n_30_138), .C1 (n_34_136), .C2 (n_40_135) );
AOI211_X1 g_23_143 (.ZN (n_23_143), .A (n_22_142), .B (n_28_139), .C1 (n_32_137), .C2 (n_38_136) );
AOI211_X1 g_25_142 (.ZN (n_25_142), .A (n_21_144), .B (n_26_140), .C1 (n_30_138), .C2 (n_36_135) );
AOI211_X1 g_27_141 (.ZN (n_27_141), .A (n_23_143), .B (n_24_141), .C1 (n_28_139), .C2 (n_34_136) );
AOI211_X1 g_29_140 (.ZN (n_29_140), .A (n_25_142), .B (n_22_142), .C1 (n_26_140), .C2 (n_32_137) );
AOI211_X1 g_31_139 (.ZN (n_31_139), .A (n_27_141), .B (n_21_144), .C1 (n_24_141), .C2 (n_30_138) );
AOI211_X1 g_33_138 (.ZN (n_33_138), .A (n_29_140), .B (n_23_143), .C1 (n_22_142), .C2 (n_28_139) );
AOI211_X1 g_35_137 (.ZN (n_35_137), .A (n_31_139), .B (n_25_142), .C1 (n_21_144), .C2 (n_26_140) );
AOI211_X1 g_37_138 (.ZN (n_37_138), .A (n_33_138), .B (n_27_141), .C1 (n_23_143), .C2 (n_24_141) );
AOI211_X1 g_36_136 (.ZN (n_36_136), .A (n_35_137), .B (n_29_140), .C1 (n_25_142), .C2 (n_22_142) );
AOI211_X1 g_34_137 (.ZN (n_34_137), .A (n_37_138), .B (n_31_139), .C1 (n_27_141), .C2 (n_21_144) );
AOI211_X1 g_32_138 (.ZN (n_32_138), .A (n_36_136), .B (n_33_138), .C1 (n_29_140), .C2 (n_23_143) );
AOI211_X1 g_30_139 (.ZN (n_30_139), .A (n_34_137), .B (n_35_137), .C1 (n_31_139), .C2 (n_25_142) );
AOI211_X1 g_28_140 (.ZN (n_28_140), .A (n_32_138), .B (n_37_138), .C1 (n_33_138), .C2 (n_27_141) );
AOI211_X1 g_26_141 (.ZN (n_26_141), .A (n_30_139), .B (n_36_136), .C1 (n_35_137), .C2 (n_29_140) );
AOI211_X1 g_25_143 (.ZN (n_25_143), .A (n_28_140), .B (n_34_137), .C1 (n_37_138), .C2 (n_31_139) );
AOI211_X1 g_23_144 (.ZN (n_23_144), .A (n_26_141), .B (n_32_138), .C1 (n_36_136), .C2 (n_33_138) );
AOI211_X1 g_22_146 (.ZN (n_22_146), .A (n_25_143), .B (n_30_139), .C1 (n_34_137), .C2 (n_35_137) );
AOI211_X1 g_20_145 (.ZN (n_20_145), .A (n_23_144), .B (n_28_140), .C1 (n_32_138), .C2 (n_37_138) );
AOI211_X1 g_19_147 (.ZN (n_19_147), .A (n_22_146), .B (n_26_141), .C1 (n_30_139), .C2 (n_36_136) );
AOI211_X1 g_21_148 (.ZN (n_21_148), .A (n_20_145), .B (n_25_143), .C1 (n_28_140), .C2 (n_34_137) );
AOI211_X1 g_22_150 (.ZN (n_22_150), .A (n_19_147), .B (n_23_144), .C1 (n_26_141), .C2 (n_32_138) );
AOI211_X1 g_20_149 (.ZN (n_20_149), .A (n_21_148), .B (n_22_146), .C1 (n_25_143), .C2 (n_30_139) );
AOI211_X1 g_21_147 (.ZN (n_21_147), .A (n_22_150), .B (n_20_145), .C1 (n_23_144), .C2 (n_28_140) );
AOI211_X1 g_23_148 (.ZN (n_23_148), .A (n_20_149), .B (n_19_147), .C1 (n_22_146), .C2 (n_26_141) );
AOI211_X1 g_24_146 (.ZN (n_24_146), .A (n_21_147), .B (n_21_148), .C1 (n_20_145), .C2 (n_25_143) );
AOI211_X1 g_22_145 (.ZN (n_22_145), .A (n_23_148), .B (n_22_150), .C1 (n_19_147), .C2 (n_23_144) );
AOI211_X1 g_24_144 (.ZN (n_24_144), .A (n_24_146), .B (n_20_149), .C1 (n_21_148), .C2 (n_22_146) );
AOI211_X1 g_26_143 (.ZN (n_26_143), .A (n_22_145), .B (n_21_147), .C1 (n_22_150), .C2 (n_20_145) );
AOI211_X1 g_28_142 (.ZN (n_28_142), .A (n_24_144), .B (n_23_148), .C1 (n_20_149), .C2 (n_19_147) );
AOI211_X1 g_30_141 (.ZN (n_30_141), .A (n_26_143), .B (n_24_146), .C1 (n_21_147), .C2 (n_21_148) );
AOI211_X1 g_32_140 (.ZN (n_32_140), .A (n_28_142), .B (n_22_145), .C1 (n_23_148), .C2 (n_22_150) );
AOI211_X1 g_34_139 (.ZN (n_34_139), .A (n_30_141), .B (n_24_144), .C1 (n_24_146), .C2 (n_20_149) );
AOI211_X1 g_36_138 (.ZN (n_36_138), .A (n_32_140), .B (n_26_143), .C1 (n_22_145), .C2 (n_21_147) );
AOI211_X1 g_38_137 (.ZN (n_38_137), .A (n_34_139), .B (n_28_142), .C1 (n_24_144), .C2 (n_23_148) );
AOI211_X1 g_40_136 (.ZN (n_40_136), .A (n_36_138), .B (n_30_141), .C1 (n_26_143), .C2 (n_24_146) );
AOI211_X1 g_42_135 (.ZN (n_42_135), .A (n_38_137), .B (n_32_140), .C1 (n_28_142), .C2 (n_22_145) );
AOI211_X1 g_44_134 (.ZN (n_44_134), .A (n_40_136), .B (n_34_139), .C1 (n_30_141), .C2 (n_24_144) );
AOI211_X1 g_46_133 (.ZN (n_46_133), .A (n_42_135), .B (n_36_138), .C1 (n_32_140), .C2 (n_26_143) );
AOI211_X1 g_48_132 (.ZN (n_48_132), .A (n_44_134), .B (n_38_137), .C1 (n_34_139), .C2 (n_28_142) );
AOI211_X1 g_50_131 (.ZN (n_50_131), .A (n_46_133), .B (n_40_136), .C1 (n_36_138), .C2 (n_30_141) );
AOI211_X1 g_48_130 (.ZN (n_48_130), .A (n_48_132), .B (n_42_135), .C1 (n_38_137), .C2 (n_32_140) );
AOI211_X1 g_50_129 (.ZN (n_50_129), .A (n_50_131), .B (n_44_134), .C1 (n_40_136), .C2 (n_34_139) );
AOI211_X1 g_51_131 (.ZN (n_51_131), .A (n_48_130), .B (n_46_133), .C1 (n_42_135), .C2 (n_36_138) );
AOI211_X1 g_49_132 (.ZN (n_49_132), .A (n_50_129), .B (n_48_132), .C1 (n_44_134), .C2 (n_38_137) );
AOI211_X1 g_48_134 (.ZN (n_48_134), .A (n_51_131), .B (n_50_131), .C1 (n_46_133), .C2 (n_40_136) );
AOI211_X1 g_47_132 (.ZN (n_47_132), .A (n_49_132), .B (n_48_130), .C1 (n_48_132), .C2 (n_42_135) );
AOI211_X1 g_49_131 (.ZN (n_49_131), .A (n_48_134), .B (n_50_129), .C1 (n_50_131), .C2 (n_44_134) );
AOI211_X1 g_51_130 (.ZN (n_51_130), .A (n_47_132), .B (n_51_131), .C1 (n_48_130), .C2 (n_46_133) );
AOI211_X1 g_53_129 (.ZN (n_53_129), .A (n_49_131), .B (n_49_132), .C1 (n_50_129), .C2 (n_48_132) );
AOI211_X1 g_52_131 (.ZN (n_52_131), .A (n_51_130), .B (n_48_134), .C1 (n_51_131), .C2 (n_50_131) );
AOI211_X1 g_54_130 (.ZN (n_54_130), .A (n_53_129), .B (n_47_132), .C1 (n_49_132), .C2 (n_48_130) );
AOI211_X1 g_56_129 (.ZN (n_56_129), .A (n_52_131), .B (n_49_131), .C1 (n_48_134), .C2 (n_50_129) );
AOI211_X1 g_55_131 (.ZN (n_55_131), .A (n_54_130), .B (n_51_130), .C1 (n_47_132), .C2 (n_51_131) );
AOI211_X1 g_54_129 (.ZN (n_54_129), .A (n_56_129), .B (n_53_129), .C1 (n_49_131), .C2 (n_49_132) );
AOI211_X1 g_52_130 (.ZN (n_52_130), .A (n_55_131), .B (n_52_131), .C1 (n_51_130), .C2 (n_48_134) );
AOI211_X1 g_53_132 (.ZN (n_53_132), .A (n_54_129), .B (n_54_130), .C1 (n_53_129), .C2 (n_47_132) );
AOI211_X1 g_51_133 (.ZN (n_51_133), .A (n_52_130), .B (n_56_129), .C1 (n_52_131), .C2 (n_49_131) );
AOI211_X1 g_49_134 (.ZN (n_49_134), .A (n_53_132), .B (n_55_131), .C1 (n_54_130), .C2 (n_51_130) );
AOI211_X1 g_50_132 (.ZN (n_50_132), .A (n_51_133), .B (n_54_129), .C1 (n_56_129), .C2 (n_53_129) );
AOI211_X1 g_48_133 (.ZN (n_48_133), .A (n_49_134), .B (n_52_130), .C1 (n_55_131), .C2 (n_52_131) );
AOI211_X1 g_46_134 (.ZN (n_46_134), .A (n_50_132), .B (n_53_132), .C1 (n_54_129), .C2 (n_54_130) );
AOI211_X1 g_44_135 (.ZN (n_44_135), .A (n_48_133), .B (n_51_133), .C1 (n_52_130), .C2 (n_56_129) );
AOI211_X1 g_45_133 (.ZN (n_45_133), .A (n_46_134), .B (n_49_134), .C1 (n_53_132), .C2 (n_55_131) );
AOI211_X1 g_43_134 (.ZN (n_43_134), .A (n_44_135), .B (n_50_132), .C1 (n_51_133), .C2 (n_54_129) );
AOI211_X1 g_41_135 (.ZN (n_41_135), .A (n_45_133), .B (n_48_133), .C1 (n_49_134), .C2 (n_52_130) );
AOI211_X1 g_39_136 (.ZN (n_39_136), .A (n_43_134), .B (n_46_134), .C1 (n_50_132), .C2 (n_53_132) );
AOI211_X1 g_37_137 (.ZN (n_37_137), .A (n_41_135), .B (n_44_135), .C1 (n_48_133), .C2 (n_51_133) );
AOI211_X1 g_35_138 (.ZN (n_35_138), .A (n_39_136), .B (n_45_133), .C1 (n_46_134), .C2 (n_49_134) );
AOI211_X1 g_33_139 (.ZN (n_33_139), .A (n_37_137), .B (n_43_134), .C1 (n_44_135), .C2 (n_50_132) );
AOI211_X1 g_31_140 (.ZN (n_31_140), .A (n_35_138), .B (n_41_135), .C1 (n_45_133), .C2 (n_48_133) );
AOI211_X1 g_29_141 (.ZN (n_29_141), .A (n_33_139), .B (n_39_136), .C1 (n_43_134), .C2 (n_46_134) );
AOI211_X1 g_27_142 (.ZN (n_27_142), .A (n_31_140), .B (n_37_137), .C1 (n_41_135), .C2 (n_44_135) );
AOI211_X1 g_26_144 (.ZN (n_26_144), .A (n_29_141), .B (n_35_138), .C1 (n_39_136), .C2 (n_45_133) );
AOI211_X1 g_24_143 (.ZN (n_24_143), .A (n_27_142), .B (n_33_139), .C1 (n_37_137), .C2 (n_43_134) );
AOI211_X1 g_22_144 (.ZN (n_22_144), .A (n_26_144), .B (n_31_140), .C1 (n_35_138), .C2 (n_41_135) );
AOI211_X1 g_21_146 (.ZN (n_21_146), .A (n_24_143), .B (n_29_141), .C1 (n_33_139), .C2 (n_39_136) );
AOI211_X1 g_23_145 (.ZN (n_23_145), .A (n_22_144), .B (n_27_142), .C1 (n_31_140), .C2 (n_37_137) );
AOI211_X1 g_25_144 (.ZN (n_25_144), .A (n_21_146), .B (n_26_144), .C1 (n_29_141), .C2 (n_35_138) );
AOI211_X1 g_26_142 (.ZN (n_26_142), .A (n_23_145), .B (n_24_143), .C1 (n_27_142), .C2 (n_33_139) );
AOI211_X1 g_28_141 (.ZN (n_28_141), .A (n_25_144), .B (n_22_144), .C1 (n_26_144), .C2 (n_31_140) );
AOI211_X1 g_30_140 (.ZN (n_30_140), .A (n_26_142), .B (n_21_146), .C1 (n_24_143), .C2 (n_29_141) );
AOI211_X1 g_32_139 (.ZN (n_32_139), .A (n_28_141), .B (n_23_145), .C1 (n_22_144), .C2 (n_27_142) );
AOI211_X1 g_34_138 (.ZN (n_34_138), .A (n_30_140), .B (n_25_144), .C1 (n_21_146), .C2 (n_26_144) );
AOI211_X1 g_36_137 (.ZN (n_36_137), .A (n_32_139), .B (n_26_142), .C1 (n_23_145), .C2 (n_24_143) );
AOI211_X1 g_35_139 (.ZN (n_35_139), .A (n_34_138), .B (n_28_141), .C1 (n_25_144), .C2 (n_22_144) );
AOI211_X1 g_33_140 (.ZN (n_33_140), .A (n_36_137), .B (n_30_140), .C1 (n_26_142), .C2 (n_21_146) );
AOI211_X1 g_31_141 (.ZN (n_31_141), .A (n_35_139), .B (n_32_139), .C1 (n_28_141), .C2 (n_23_145) );
AOI211_X1 g_29_142 (.ZN (n_29_142), .A (n_33_140), .B (n_34_138), .C1 (n_30_140), .C2 (n_25_144) );
AOI211_X1 g_27_143 (.ZN (n_27_143), .A (n_31_141), .B (n_36_137), .C1 (n_32_139), .C2 (n_26_142) );
AOI211_X1 g_26_145 (.ZN (n_26_145), .A (n_29_142), .B (n_35_139), .C1 (n_34_138), .C2 (n_28_141) );
AOI211_X1 g_28_144 (.ZN (n_28_144), .A (n_27_143), .B (n_33_140), .C1 (n_36_137), .C2 (n_30_140) );
AOI211_X1 g_30_143 (.ZN (n_30_143), .A (n_26_145), .B (n_31_141), .C1 (n_35_139), .C2 (n_32_139) );
AOI211_X1 g_32_142 (.ZN (n_32_142), .A (n_28_144), .B (n_29_142), .C1 (n_33_140), .C2 (n_34_138) );
AOI211_X1 g_34_141 (.ZN (n_34_141), .A (n_30_143), .B (n_27_143), .C1 (n_31_141), .C2 (n_36_137) );
AOI211_X1 g_36_140 (.ZN (n_36_140), .A (n_32_142), .B (n_26_145), .C1 (n_29_142), .C2 (n_35_139) );
AOI211_X1 g_38_139 (.ZN (n_38_139), .A (n_34_141), .B (n_28_144), .C1 (n_27_143), .C2 (n_33_140) );
AOI211_X1 g_40_138 (.ZN (n_40_138), .A (n_36_140), .B (n_30_143), .C1 (n_26_145), .C2 (n_31_141) );
AOI211_X1 g_42_137 (.ZN (n_42_137), .A (n_38_139), .B (n_32_142), .C1 (n_28_144), .C2 (n_29_142) );
AOI211_X1 g_44_136 (.ZN (n_44_136), .A (n_40_138), .B (n_34_141), .C1 (n_30_143), .C2 (n_27_143) );
AOI211_X1 g_46_135 (.ZN (n_46_135), .A (n_42_137), .B (n_36_140), .C1 (n_32_142), .C2 (n_26_145) );
AOI211_X1 g_45_137 (.ZN (n_45_137), .A (n_44_136), .B (n_38_139), .C1 (n_34_141), .C2 (n_28_144) );
AOI211_X1 g_43_136 (.ZN (n_43_136), .A (n_46_135), .B (n_40_138), .C1 (n_36_140), .C2 (n_30_143) );
AOI211_X1 g_45_135 (.ZN (n_45_135), .A (n_45_137), .B (n_42_137), .C1 (n_38_139), .C2 (n_32_142) );
AOI211_X1 g_47_134 (.ZN (n_47_134), .A (n_43_136), .B (n_44_136), .C1 (n_40_138), .C2 (n_34_141) );
AOI211_X1 g_49_133 (.ZN (n_49_133), .A (n_45_135), .B (n_46_135), .C1 (n_42_137), .C2 (n_36_140) );
AOI211_X1 g_51_132 (.ZN (n_51_132), .A (n_47_134), .B (n_45_137), .C1 (n_44_136), .C2 (n_38_139) );
AOI211_X1 g_53_131 (.ZN (n_53_131), .A (n_49_133), .B (n_43_136), .C1 (n_46_135), .C2 (n_40_138) );
AOI211_X1 g_55_130 (.ZN (n_55_130), .A (n_51_132), .B (n_45_135), .C1 (n_45_137), .C2 (n_42_137) );
AOI211_X1 g_56_128 (.ZN (n_56_128), .A (n_53_131), .B (n_47_134), .C1 (n_43_136), .C2 (n_44_136) );
AOI211_X1 g_58_127 (.ZN (n_58_127), .A (n_55_130), .B (n_49_133), .C1 (n_45_135), .C2 (n_46_135) );
AOI211_X1 g_60_126 (.ZN (n_60_126), .A (n_56_128), .B (n_51_132), .C1 (n_47_134), .C2 (n_45_137) );
AOI211_X1 g_62_125 (.ZN (n_62_125), .A (n_58_127), .B (n_53_131), .C1 (n_49_133), .C2 (n_43_136) );
AOI211_X1 g_64_124 (.ZN (n_64_124), .A (n_60_126), .B (n_55_130), .C1 (n_51_132), .C2 (n_45_135) );
AOI211_X1 g_66_123 (.ZN (n_66_123), .A (n_62_125), .B (n_56_128), .C1 (n_53_131), .C2 (n_47_134) );
AOI211_X1 g_68_122 (.ZN (n_68_122), .A (n_64_124), .B (n_58_127), .C1 (n_55_130), .C2 (n_49_133) );
AOI211_X1 g_67_124 (.ZN (n_67_124), .A (n_66_123), .B (n_60_126), .C1 (n_56_128), .C2 (n_51_132) );
AOI211_X1 g_69_123 (.ZN (n_69_123), .A (n_68_122), .B (n_62_125), .C1 (n_58_127), .C2 (n_53_131) );
AOI211_X1 g_71_122 (.ZN (n_71_122), .A (n_67_124), .B (n_64_124), .C1 (n_60_126), .C2 (n_55_130) );
AOI211_X1 g_73_121 (.ZN (n_73_121), .A (n_69_123), .B (n_66_123), .C1 (n_62_125), .C2 (n_56_128) );
AOI211_X1 g_75_120 (.ZN (n_75_120), .A (n_71_122), .B (n_68_122), .C1 (n_64_124), .C2 (n_58_127) );
AOI211_X1 g_77_119 (.ZN (n_77_119), .A (n_73_121), .B (n_67_124), .C1 (n_66_123), .C2 (n_60_126) );
AOI211_X1 g_79_118 (.ZN (n_79_118), .A (n_75_120), .B (n_69_123), .C1 (n_68_122), .C2 (n_62_125) );
AOI211_X1 g_81_117 (.ZN (n_81_117), .A (n_77_119), .B (n_71_122), .C1 (n_67_124), .C2 (n_64_124) );
AOI211_X1 g_83_116 (.ZN (n_83_116), .A (n_79_118), .B (n_73_121), .C1 (n_69_123), .C2 (n_66_123) );
AOI211_X1 g_85_115 (.ZN (n_85_115), .A (n_81_117), .B (n_75_120), .C1 (n_71_122), .C2 (n_68_122) );
AOI211_X1 g_87_114 (.ZN (n_87_114), .A (n_83_116), .B (n_77_119), .C1 (n_73_121), .C2 (n_67_124) );
AOI211_X1 g_89_113 (.ZN (n_89_113), .A (n_85_115), .B (n_79_118), .C1 (n_75_120), .C2 (n_69_123) );
AOI211_X1 g_91_112 (.ZN (n_91_112), .A (n_87_114), .B (n_81_117), .C1 (n_77_119), .C2 (n_71_122) );
AOI211_X1 g_93_111 (.ZN (n_93_111), .A (n_89_113), .B (n_83_116), .C1 (n_79_118), .C2 (n_73_121) );
AOI211_X1 g_92_113 (.ZN (n_92_113), .A (n_91_112), .B (n_85_115), .C1 (n_81_117), .C2 (n_75_120) );
AOI211_X1 g_94_112 (.ZN (n_94_112), .A (n_93_111), .B (n_87_114), .C1 (n_83_116), .C2 (n_77_119) );
AOI211_X1 g_96_111 (.ZN (n_96_111), .A (n_92_113), .B (n_89_113), .C1 (n_85_115), .C2 (n_79_118) );
AOI211_X1 g_98_110 (.ZN (n_98_110), .A (n_94_112), .B (n_91_112), .C1 (n_87_114), .C2 (n_81_117) );
AOI211_X1 g_100_109 (.ZN (n_100_109), .A (n_96_111), .B (n_93_111), .C1 (n_89_113), .C2 (n_83_116) );
AOI211_X1 g_102_108 (.ZN (n_102_108), .A (n_98_110), .B (n_92_113), .C1 (n_91_112), .C2 (n_85_115) );
AOI211_X1 g_104_107 (.ZN (n_104_107), .A (n_100_109), .B (n_94_112), .C1 (n_93_111), .C2 (n_87_114) );
AOI211_X1 g_106_106 (.ZN (n_106_106), .A (n_102_108), .B (n_96_111), .C1 (n_92_113), .C2 (n_89_113) );
AOI211_X1 g_108_105 (.ZN (n_108_105), .A (n_104_107), .B (n_98_110), .C1 (n_94_112), .C2 (n_91_112) );
AOI211_X1 g_110_104 (.ZN (n_110_104), .A (n_106_106), .B (n_100_109), .C1 (n_96_111), .C2 (n_93_111) );
AOI211_X1 g_112_103 (.ZN (n_112_103), .A (n_108_105), .B (n_102_108), .C1 (n_98_110), .C2 (n_92_113) );
AOI211_X1 g_114_102 (.ZN (n_114_102), .A (n_110_104), .B (n_104_107), .C1 (n_100_109), .C2 (n_94_112) );
AOI211_X1 g_116_101 (.ZN (n_116_101), .A (n_112_103), .B (n_106_106), .C1 (n_102_108), .C2 (n_96_111) );
AOI211_X1 g_118_100 (.ZN (n_118_100), .A (n_114_102), .B (n_108_105), .C1 (n_104_107), .C2 (n_98_110) );
AOI211_X1 g_117_102 (.ZN (n_117_102), .A (n_116_101), .B (n_110_104), .C1 (n_106_106), .C2 (n_100_109) );
AOI211_X1 g_115_103 (.ZN (n_115_103), .A (n_118_100), .B (n_112_103), .C1 (n_108_105), .C2 (n_102_108) );
AOI211_X1 g_113_102 (.ZN (n_113_102), .A (n_117_102), .B (n_114_102), .C1 (n_110_104), .C2 (n_104_107) );
AOI211_X1 g_111_103 (.ZN (n_111_103), .A (n_115_103), .B (n_116_101), .C1 (n_112_103), .C2 (n_106_106) );
AOI211_X1 g_109_104 (.ZN (n_109_104), .A (n_113_102), .B (n_118_100), .C1 (n_114_102), .C2 (n_108_105) );
AOI211_X1 g_107_105 (.ZN (n_107_105), .A (n_111_103), .B (n_117_102), .C1 (n_116_101), .C2 (n_110_104) );
AOI211_X1 g_105_106 (.ZN (n_105_106), .A (n_109_104), .B (n_115_103), .C1 (n_118_100), .C2 (n_112_103) );
AOI211_X1 g_103_107 (.ZN (n_103_107), .A (n_107_105), .B (n_113_102), .C1 (n_117_102), .C2 (n_114_102) );
AOI211_X1 g_101_108 (.ZN (n_101_108), .A (n_105_106), .B (n_111_103), .C1 (n_115_103), .C2 (n_116_101) );
AOI211_X1 g_99_109 (.ZN (n_99_109), .A (n_103_107), .B (n_109_104), .C1 (n_113_102), .C2 (n_118_100) );
AOI211_X1 g_97_110 (.ZN (n_97_110), .A (n_101_108), .B (n_107_105), .C1 (n_111_103), .C2 (n_117_102) );
AOI211_X1 g_95_111 (.ZN (n_95_111), .A (n_99_109), .B (n_105_106), .C1 (n_109_104), .C2 (n_115_103) );
AOI211_X1 g_93_112 (.ZN (n_93_112), .A (n_97_110), .B (n_103_107), .C1 (n_107_105), .C2 (n_113_102) );
AOI211_X1 g_91_113 (.ZN (n_91_113), .A (n_95_111), .B (n_101_108), .C1 (n_105_106), .C2 (n_111_103) );
AOI211_X1 g_89_112 (.ZN (n_89_112), .A (n_93_112), .B (n_99_109), .C1 (n_103_107), .C2 (n_109_104) );
AOI211_X1 g_87_113 (.ZN (n_87_113), .A (n_91_113), .B (n_97_110), .C1 (n_101_108), .C2 (n_107_105) );
AOI211_X1 g_85_114 (.ZN (n_85_114), .A (n_89_112), .B (n_95_111), .C1 (n_99_109), .C2 (n_105_106) );
AOI211_X1 g_83_115 (.ZN (n_83_115), .A (n_87_113), .B (n_93_112), .C1 (n_97_110), .C2 (n_103_107) );
AOI211_X1 g_81_116 (.ZN (n_81_116), .A (n_85_114), .B (n_91_113), .C1 (n_95_111), .C2 (n_101_108) );
AOI211_X1 g_79_117 (.ZN (n_79_117), .A (n_83_115), .B (n_89_112), .C1 (n_93_112), .C2 (n_99_109) );
AOI211_X1 g_77_118 (.ZN (n_77_118), .A (n_81_116), .B (n_87_113), .C1 (n_91_113), .C2 (n_97_110) );
AOI211_X1 g_75_119 (.ZN (n_75_119), .A (n_79_117), .B (n_85_114), .C1 (n_89_112), .C2 (n_95_111) );
AOI211_X1 g_73_120 (.ZN (n_73_120), .A (n_77_118), .B (n_83_115), .C1 (n_87_113), .C2 (n_93_112) );
AOI211_X1 g_71_121 (.ZN (n_71_121), .A (n_75_119), .B (n_81_116), .C1 (n_85_114), .C2 (n_91_113) );
AOI211_X1 g_69_122 (.ZN (n_69_122), .A (n_73_120), .B (n_79_117), .C1 (n_83_115), .C2 (n_89_112) );
AOI211_X1 g_67_123 (.ZN (n_67_123), .A (n_71_121), .B (n_77_118), .C1 (n_81_116), .C2 (n_87_113) );
AOI211_X1 g_65_124 (.ZN (n_65_124), .A (n_69_122), .B (n_75_119), .C1 (n_79_117), .C2 (n_85_114) );
AOI211_X1 g_63_125 (.ZN (n_63_125), .A (n_67_123), .B (n_73_120), .C1 (n_77_118), .C2 (n_83_115) );
AOI211_X1 g_61_126 (.ZN (n_61_126), .A (n_65_124), .B (n_71_121), .C1 (n_75_119), .C2 (n_81_116) );
AOI211_X1 g_59_127 (.ZN (n_59_127), .A (n_63_125), .B (n_69_122), .C1 (n_73_120), .C2 (n_79_117) );
AOI211_X1 g_57_128 (.ZN (n_57_128), .A (n_61_126), .B (n_67_123), .C1 (n_71_121), .C2 (n_77_118) );
AOI211_X1 g_55_129 (.ZN (n_55_129), .A (n_59_127), .B (n_65_124), .C1 (n_69_122), .C2 (n_75_119) );
AOI211_X1 g_57_130 (.ZN (n_57_130), .A (n_57_128), .B (n_63_125), .C1 (n_67_123), .C2 (n_73_120) );
AOI211_X1 g_59_129 (.ZN (n_59_129), .A (n_55_129), .B (n_61_126), .C1 (n_65_124), .C2 (n_71_121) );
AOI211_X1 g_61_128 (.ZN (n_61_128), .A (n_57_130), .B (n_59_127), .C1 (n_63_125), .C2 (n_69_122) );
AOI211_X1 g_63_127 (.ZN (n_63_127), .A (n_59_129), .B (n_57_128), .C1 (n_61_126), .C2 (n_67_123) );
AOI211_X1 g_64_125 (.ZN (n_64_125), .A (n_61_128), .B (n_55_129), .C1 (n_59_127), .C2 (n_65_124) );
AOI211_X1 g_66_124 (.ZN (n_66_124), .A (n_63_127), .B (n_57_130), .C1 (n_57_128), .C2 (n_63_125) );
AOI211_X1 g_68_123 (.ZN (n_68_123), .A (n_64_125), .B (n_59_129), .C1 (n_55_129), .C2 (n_61_126) );
AOI211_X1 g_70_122 (.ZN (n_70_122), .A (n_66_124), .B (n_61_128), .C1 (n_57_130), .C2 (n_59_127) );
AOI211_X1 g_72_121 (.ZN (n_72_121), .A (n_68_123), .B (n_63_127), .C1 (n_59_129), .C2 (n_57_128) );
AOI211_X1 g_74_120 (.ZN (n_74_120), .A (n_70_122), .B (n_64_125), .C1 (n_61_128), .C2 (n_55_129) );
AOI211_X1 g_76_119 (.ZN (n_76_119), .A (n_72_121), .B (n_66_124), .C1 (n_63_127), .C2 (n_57_130) );
AOI211_X1 g_78_118 (.ZN (n_78_118), .A (n_74_120), .B (n_68_123), .C1 (n_64_125), .C2 (n_59_129) );
AOI211_X1 g_80_117 (.ZN (n_80_117), .A (n_76_119), .B (n_70_122), .C1 (n_66_124), .C2 (n_61_128) );
AOI211_X1 g_79_119 (.ZN (n_79_119), .A (n_78_118), .B (n_72_121), .C1 (n_68_123), .C2 (n_63_127) );
AOI211_X1 g_81_118 (.ZN (n_81_118), .A (n_80_117), .B (n_74_120), .C1 (n_70_122), .C2 (n_64_125) );
AOI211_X1 g_83_117 (.ZN (n_83_117), .A (n_79_119), .B (n_76_119), .C1 (n_72_121), .C2 (n_66_124) );
AOI211_X1 g_85_116 (.ZN (n_85_116), .A (n_81_118), .B (n_78_118), .C1 (n_74_120), .C2 (n_68_123) );
AOI211_X1 g_87_115 (.ZN (n_87_115), .A (n_83_117), .B (n_80_117), .C1 (n_76_119), .C2 (n_70_122) );
AOI211_X1 g_89_114 (.ZN (n_89_114), .A (n_85_116), .B (n_79_119), .C1 (n_78_118), .C2 (n_72_121) );
AOI211_X1 g_88_116 (.ZN (n_88_116), .A (n_87_115), .B (n_81_118), .C1 (n_80_117), .C2 (n_74_120) );
AOI211_X1 g_86_115 (.ZN (n_86_115), .A (n_89_114), .B (n_83_117), .C1 (n_79_119), .C2 (n_76_119) );
AOI211_X1 g_88_114 (.ZN (n_88_114), .A (n_88_116), .B (n_85_116), .C1 (n_81_118), .C2 (n_78_118) );
AOI211_X1 g_90_113 (.ZN (n_90_113), .A (n_86_115), .B (n_87_115), .C1 (n_83_117), .C2 (n_80_117) );
AOI211_X1 g_92_112 (.ZN (n_92_112), .A (n_88_114), .B (n_89_114), .C1 (n_85_116), .C2 (n_79_119) );
AOI211_X1 g_94_111 (.ZN (n_94_111), .A (n_90_113), .B (n_88_116), .C1 (n_87_115), .C2 (n_81_118) );
AOI211_X1 g_96_110 (.ZN (n_96_110), .A (n_92_112), .B (n_86_115), .C1 (n_89_114), .C2 (n_83_117) );
AOI211_X1 g_98_109 (.ZN (n_98_109), .A (n_94_111), .B (n_88_114), .C1 (n_88_116), .C2 (n_85_116) );
AOI211_X1 g_100_108 (.ZN (n_100_108), .A (n_96_110), .B (n_90_113), .C1 (n_86_115), .C2 (n_87_115) );
AOI211_X1 g_102_107 (.ZN (n_102_107), .A (n_98_109), .B (n_92_112), .C1 (n_88_114), .C2 (n_89_114) );
AOI211_X1 g_104_106 (.ZN (n_104_106), .A (n_100_108), .B (n_94_111), .C1 (n_90_113), .C2 (n_88_116) );
AOI211_X1 g_103_108 (.ZN (n_103_108), .A (n_102_107), .B (n_96_110), .C1 (n_92_112), .C2 (n_86_115) );
AOI211_X1 g_105_107 (.ZN (n_105_107), .A (n_104_106), .B (n_98_109), .C1 (n_94_111), .C2 (n_88_114) );
AOI211_X1 g_107_106 (.ZN (n_107_106), .A (n_103_108), .B (n_100_108), .C1 (n_96_110), .C2 (n_90_113) );
AOI211_X1 g_109_105 (.ZN (n_109_105), .A (n_105_107), .B (n_102_107), .C1 (n_98_109), .C2 (n_92_112) );
AOI211_X1 g_111_104 (.ZN (n_111_104), .A (n_107_106), .B (n_104_106), .C1 (n_100_108), .C2 (n_94_111) );
AOI211_X1 g_113_103 (.ZN (n_113_103), .A (n_109_105), .B (n_103_108), .C1 (n_102_107), .C2 (n_96_110) );
AOI211_X1 g_115_102 (.ZN (n_115_102), .A (n_111_104), .B (n_105_107), .C1 (n_104_106), .C2 (n_98_109) );
AOI211_X1 g_117_101 (.ZN (n_117_101), .A (n_113_103), .B (n_107_106), .C1 (n_103_108), .C2 (n_100_108) );
AOI211_X1 g_118_103 (.ZN (n_118_103), .A (n_115_102), .B (n_109_105), .C1 (n_105_107), .C2 (n_102_107) );
AOI211_X1 g_116_104 (.ZN (n_116_104), .A (n_117_101), .B (n_111_104), .C1 (n_107_106), .C2 (n_104_106) );
AOI211_X1 g_114_105 (.ZN (n_114_105), .A (n_118_103), .B (n_113_103), .C1 (n_109_105), .C2 (n_103_108) );
AOI211_X1 g_112_104 (.ZN (n_112_104), .A (n_116_104), .B (n_115_102), .C1 (n_111_104), .C2 (n_105_107) );
AOI211_X1 g_110_105 (.ZN (n_110_105), .A (n_114_105), .B (n_117_101), .C1 (n_113_103), .C2 (n_107_106) );
AOI211_X1 g_108_106 (.ZN (n_108_106), .A (n_112_104), .B (n_118_103), .C1 (n_115_102), .C2 (n_109_105) );
AOI211_X1 g_106_107 (.ZN (n_106_107), .A (n_110_105), .B (n_116_104), .C1 (n_117_101), .C2 (n_111_104) );
AOI211_X1 g_104_108 (.ZN (n_104_108), .A (n_108_106), .B (n_114_105), .C1 (n_118_103), .C2 (n_113_103) );
AOI211_X1 g_102_109 (.ZN (n_102_109), .A (n_106_107), .B (n_112_104), .C1 (n_116_104), .C2 (n_115_102) );
AOI211_X1 g_100_110 (.ZN (n_100_110), .A (n_104_108), .B (n_110_105), .C1 (n_114_105), .C2 (n_117_101) );
AOI211_X1 g_98_111 (.ZN (n_98_111), .A (n_102_109), .B (n_108_106), .C1 (n_112_104), .C2 (n_118_103) );
AOI211_X1 g_96_112 (.ZN (n_96_112), .A (n_100_110), .B (n_106_107), .C1 (n_110_105), .C2 (n_116_104) );
AOI211_X1 g_94_113 (.ZN (n_94_113), .A (n_98_111), .B (n_104_108), .C1 (n_108_106), .C2 (n_114_105) );
AOI211_X1 g_92_114 (.ZN (n_92_114), .A (n_96_112), .B (n_102_109), .C1 (n_106_107), .C2 (n_112_104) );
AOI211_X1 g_90_115 (.ZN (n_90_115), .A (n_94_113), .B (n_100_110), .C1 (n_104_108), .C2 (n_110_105) );
AOI211_X1 g_89_117 (.ZN (n_89_117), .A (n_92_114), .B (n_98_111), .C1 (n_102_109), .C2 (n_108_106) );
AOI211_X1 g_88_115 (.ZN (n_88_115), .A (n_90_115), .B (n_96_112), .C1 (n_100_110), .C2 (n_106_107) );
AOI211_X1 g_90_114 (.ZN (n_90_114), .A (n_89_117), .B (n_94_113), .C1 (n_98_111), .C2 (n_104_108) );
AOI211_X1 g_89_116 (.ZN (n_89_116), .A (n_88_115), .B (n_92_114), .C1 (n_96_112), .C2 (n_102_109) );
AOI211_X1 g_91_115 (.ZN (n_91_115), .A (n_90_114), .B (n_90_115), .C1 (n_94_113), .C2 (n_100_110) );
AOI211_X1 g_93_114 (.ZN (n_93_114), .A (n_89_116), .B (n_89_117), .C1 (n_92_114), .C2 (n_98_111) );
AOI211_X1 g_95_113 (.ZN (n_95_113), .A (n_91_115), .B (n_88_115), .C1 (n_90_115), .C2 (n_96_112) );
AOI211_X1 g_97_112 (.ZN (n_97_112), .A (n_93_114), .B (n_90_114), .C1 (n_89_117), .C2 (n_94_113) );
AOI211_X1 g_99_111 (.ZN (n_99_111), .A (n_95_113), .B (n_89_116), .C1 (n_88_115), .C2 (n_92_114) );
AOI211_X1 g_101_110 (.ZN (n_101_110), .A (n_97_112), .B (n_91_115), .C1 (n_90_114), .C2 (n_90_115) );
AOI211_X1 g_103_109 (.ZN (n_103_109), .A (n_99_111), .B (n_93_114), .C1 (n_89_116), .C2 (n_89_117) );
AOI211_X1 g_105_108 (.ZN (n_105_108), .A (n_101_110), .B (n_95_113), .C1 (n_91_115), .C2 (n_88_115) );
AOI211_X1 g_107_107 (.ZN (n_107_107), .A (n_103_109), .B (n_97_112), .C1 (n_93_114), .C2 (n_90_114) );
AOI211_X1 g_109_106 (.ZN (n_109_106), .A (n_105_108), .B (n_99_111), .C1 (n_95_113), .C2 (n_89_116) );
AOI211_X1 g_111_105 (.ZN (n_111_105), .A (n_107_107), .B (n_101_110), .C1 (n_97_112), .C2 (n_91_115) );
AOI211_X1 g_113_104 (.ZN (n_113_104), .A (n_109_106), .B (n_103_109), .C1 (n_99_111), .C2 (n_93_114) );
AOI211_X1 g_112_106 (.ZN (n_112_106), .A (n_111_105), .B (n_105_108), .C1 (n_101_110), .C2 (n_95_113) );
AOI211_X1 g_110_107 (.ZN (n_110_107), .A (n_113_104), .B (n_107_107), .C1 (n_103_109), .C2 (n_97_112) );
AOI211_X1 g_108_108 (.ZN (n_108_108), .A (n_112_106), .B (n_109_106), .C1 (n_105_108), .C2 (n_99_111) );
AOI211_X1 g_106_109 (.ZN (n_106_109), .A (n_110_107), .B (n_111_105), .C1 (n_107_107), .C2 (n_101_110) );
AOI211_X1 g_104_110 (.ZN (n_104_110), .A (n_108_108), .B (n_113_104), .C1 (n_109_106), .C2 (n_103_109) );
AOI211_X1 g_102_111 (.ZN (n_102_111), .A (n_106_109), .B (n_112_106), .C1 (n_111_105), .C2 (n_105_108) );
AOI211_X1 g_101_109 (.ZN (n_101_109), .A (n_104_110), .B (n_110_107), .C1 (n_113_104), .C2 (n_107_107) );
AOI211_X1 g_99_110 (.ZN (n_99_110), .A (n_102_111), .B (n_108_108), .C1 (n_112_106), .C2 (n_109_106) );
AOI211_X1 g_97_111 (.ZN (n_97_111), .A (n_101_109), .B (n_106_109), .C1 (n_110_107), .C2 (n_111_105) );
AOI211_X1 g_95_112 (.ZN (n_95_112), .A (n_99_110), .B (n_104_110), .C1 (n_108_108), .C2 (n_113_104) );
AOI211_X1 g_93_113 (.ZN (n_93_113), .A (n_97_111), .B (n_102_111), .C1 (n_106_109), .C2 (n_112_106) );
AOI211_X1 g_91_114 (.ZN (n_91_114), .A (n_95_112), .B (n_101_109), .C1 (n_104_110), .C2 (n_110_107) );
AOI211_X1 g_89_115 (.ZN (n_89_115), .A (n_93_113), .B (n_99_110), .C1 (n_102_111), .C2 (n_108_108) );
AOI211_X1 g_87_116 (.ZN (n_87_116), .A (n_91_114), .B (n_97_111), .C1 (n_101_109), .C2 (n_106_109) );
AOI211_X1 g_85_117 (.ZN (n_85_117), .A (n_89_115), .B (n_95_112), .C1 (n_99_110), .C2 (n_104_110) );
AOI211_X1 g_83_118 (.ZN (n_83_118), .A (n_87_116), .B (n_93_113), .C1 (n_97_111), .C2 (n_102_111) );
AOI211_X1 g_84_116 (.ZN (n_84_116), .A (n_85_117), .B (n_91_114), .C1 (n_95_112), .C2 (n_101_109) );
AOI211_X1 g_82_117 (.ZN (n_82_117), .A (n_83_118), .B (n_89_115), .C1 (n_93_113), .C2 (n_99_110) );
AOI211_X1 g_80_118 (.ZN (n_80_118), .A (n_84_116), .B (n_87_116), .C1 (n_91_114), .C2 (n_97_111) );
AOI211_X1 g_78_119 (.ZN (n_78_119), .A (n_82_117), .B (n_85_117), .C1 (n_89_115), .C2 (n_95_112) );
AOI211_X1 g_76_120 (.ZN (n_76_120), .A (n_80_118), .B (n_83_118), .C1 (n_87_116), .C2 (n_93_113) );
AOI211_X1 g_74_121 (.ZN (n_74_121), .A (n_78_119), .B (n_84_116), .C1 (n_85_117), .C2 (n_91_114) );
AOI211_X1 g_72_122 (.ZN (n_72_122), .A (n_76_120), .B (n_82_117), .C1 (n_83_118), .C2 (n_89_115) );
AOI211_X1 g_70_123 (.ZN (n_70_123), .A (n_74_121), .B (n_80_118), .C1 (n_84_116), .C2 (n_87_116) );
AOI211_X1 g_68_124 (.ZN (n_68_124), .A (n_72_122), .B (n_78_119), .C1 (n_82_117), .C2 (n_85_117) );
AOI211_X1 g_66_125 (.ZN (n_66_125), .A (n_70_123), .B (n_76_120), .C1 (n_80_118), .C2 (n_83_118) );
AOI211_X1 g_64_126 (.ZN (n_64_126), .A (n_68_124), .B (n_74_121), .C1 (n_78_119), .C2 (n_84_116) );
AOI211_X1 g_62_127 (.ZN (n_62_127), .A (n_66_125), .B (n_72_122), .C1 (n_76_120), .C2 (n_82_117) );
AOI211_X1 g_60_128 (.ZN (n_60_128), .A (n_64_126), .B (n_70_123), .C1 (n_74_121), .C2 (n_80_118) );
AOI211_X1 g_58_129 (.ZN (n_58_129), .A (n_62_127), .B (n_68_124), .C1 (n_72_122), .C2 (n_78_119) );
AOI211_X1 g_56_130 (.ZN (n_56_130), .A (n_60_128), .B (n_66_125), .C1 (n_70_123), .C2 (n_76_120) );
AOI211_X1 g_54_131 (.ZN (n_54_131), .A (n_58_129), .B (n_64_126), .C1 (n_68_124), .C2 (n_74_121) );
AOI211_X1 g_52_132 (.ZN (n_52_132), .A (n_56_130), .B (n_62_127), .C1 (n_66_125), .C2 (n_72_122) );
AOI211_X1 g_50_133 (.ZN (n_50_133), .A (n_54_131), .B (n_60_128), .C1 (n_64_126), .C2 (n_70_123) );
AOI211_X1 g_49_135 (.ZN (n_49_135), .A (n_52_132), .B (n_58_129), .C1 (n_62_127), .C2 (n_68_124) );
AOI211_X1 g_47_136 (.ZN (n_47_136), .A (n_50_133), .B (n_56_130), .C1 (n_60_128), .C2 (n_66_125) );
AOI211_X1 g_46_138 (.ZN (n_46_138), .A (n_49_135), .B (n_54_131), .C1 (n_58_129), .C2 (n_64_126) );
AOI211_X1 g_45_136 (.ZN (n_45_136), .A (n_47_136), .B (n_52_132), .C1 (n_56_130), .C2 (n_62_127) );
AOI211_X1 g_47_135 (.ZN (n_47_135), .A (n_46_138), .B (n_50_133), .C1 (n_54_131), .C2 (n_60_128) );
AOI211_X1 g_46_137 (.ZN (n_46_137), .A (n_45_136), .B (n_49_135), .C1 (n_52_132), .C2 (n_58_129) );
AOI211_X1 g_48_136 (.ZN (n_48_136), .A (n_47_135), .B (n_47_136), .C1 (n_50_133), .C2 (n_56_130) );
AOI211_X1 g_50_135 (.ZN (n_50_135), .A (n_46_137), .B (n_46_138), .C1 (n_49_135), .C2 (n_54_131) );
AOI211_X1 g_52_134 (.ZN (n_52_134), .A (n_48_136), .B (n_45_136), .C1 (n_47_136), .C2 (n_52_132) );
AOI211_X1 g_54_133 (.ZN (n_54_133), .A (n_50_135), .B (n_47_135), .C1 (n_46_138), .C2 (n_50_133) );
AOI211_X1 g_56_132 (.ZN (n_56_132), .A (n_52_134), .B (n_46_137), .C1 (n_45_136), .C2 (n_49_135) );
AOI211_X1 g_58_131 (.ZN (n_58_131), .A (n_54_133), .B (n_48_136), .C1 (n_47_135), .C2 (n_47_136) );
AOI211_X1 g_57_129 (.ZN (n_57_129), .A (n_56_132), .B (n_50_135), .C1 (n_46_137), .C2 (n_46_138) );
AOI211_X1 g_59_128 (.ZN (n_59_128), .A (n_58_131), .B (n_52_134), .C1 (n_48_136), .C2 (n_45_136) );
AOI211_X1 g_61_127 (.ZN (n_61_127), .A (n_57_129), .B (n_54_133), .C1 (n_50_135), .C2 (n_47_135) );
AOI211_X1 g_63_126 (.ZN (n_63_126), .A (n_59_128), .B (n_56_132), .C1 (n_52_134), .C2 (n_46_137) );
AOI211_X1 g_65_125 (.ZN (n_65_125), .A (n_61_127), .B (n_58_131), .C1 (n_54_133), .C2 (n_48_136) );
AOI211_X1 g_64_127 (.ZN (n_64_127), .A (n_63_126), .B (n_57_129), .C1 (n_56_132), .C2 (n_50_135) );
AOI211_X1 g_66_126 (.ZN (n_66_126), .A (n_65_125), .B (n_59_128), .C1 (n_58_131), .C2 (n_52_134) );
AOI211_X1 g_68_125 (.ZN (n_68_125), .A (n_64_127), .B (n_61_127), .C1 (n_57_129), .C2 (n_54_133) );
AOI211_X1 g_70_124 (.ZN (n_70_124), .A (n_66_126), .B (n_63_126), .C1 (n_59_128), .C2 (n_56_132) );
AOI211_X1 g_72_123 (.ZN (n_72_123), .A (n_68_125), .B (n_65_125), .C1 (n_61_127), .C2 (n_58_131) );
AOI211_X1 g_74_122 (.ZN (n_74_122), .A (n_70_124), .B (n_64_127), .C1 (n_63_126), .C2 (n_57_129) );
AOI211_X1 g_76_121 (.ZN (n_76_121), .A (n_72_123), .B (n_66_126), .C1 (n_65_125), .C2 (n_59_128) );
AOI211_X1 g_78_120 (.ZN (n_78_120), .A (n_74_122), .B (n_68_125), .C1 (n_64_127), .C2 (n_61_127) );
AOI211_X1 g_80_119 (.ZN (n_80_119), .A (n_76_121), .B (n_70_124), .C1 (n_66_126), .C2 (n_63_126) );
AOI211_X1 g_82_118 (.ZN (n_82_118), .A (n_78_120), .B (n_72_123), .C1 (n_68_125), .C2 (n_65_125) );
AOI211_X1 g_84_117 (.ZN (n_84_117), .A (n_80_119), .B (n_74_122), .C1 (n_70_124), .C2 (n_64_127) );
AOI211_X1 g_86_116 (.ZN (n_86_116), .A (n_82_118), .B (n_76_121), .C1 (n_72_123), .C2 (n_66_126) );
AOI211_X1 g_87_118 (.ZN (n_87_118), .A (n_84_117), .B (n_78_120), .C1 (n_74_122), .C2 (n_68_125) );
AOI211_X1 g_85_119 (.ZN (n_85_119), .A (n_86_116), .B (n_80_119), .C1 (n_76_121), .C2 (n_70_124) );
AOI211_X1 g_86_117 (.ZN (n_86_117), .A (n_87_118), .B (n_82_118), .C1 (n_78_120), .C2 (n_72_123) );
AOI211_X1 g_84_118 (.ZN (n_84_118), .A (n_85_119), .B (n_84_117), .C1 (n_80_119), .C2 (n_74_122) );
AOI211_X1 g_82_119 (.ZN (n_82_119), .A (n_86_117), .B (n_86_116), .C1 (n_82_118), .C2 (n_76_121) );
AOI211_X1 g_80_120 (.ZN (n_80_120), .A (n_84_118), .B (n_87_118), .C1 (n_84_117), .C2 (n_78_120) );
AOI211_X1 g_78_121 (.ZN (n_78_121), .A (n_82_119), .B (n_85_119), .C1 (n_86_116), .C2 (n_80_119) );
AOI211_X1 g_76_122 (.ZN (n_76_122), .A (n_80_120), .B (n_86_117), .C1 (n_87_118), .C2 (n_82_118) );
AOI211_X1 g_77_120 (.ZN (n_77_120), .A (n_78_121), .B (n_84_118), .C1 (n_85_119), .C2 (n_84_117) );
AOI211_X1 g_75_121 (.ZN (n_75_121), .A (n_76_122), .B (n_82_119), .C1 (n_86_117), .C2 (n_86_116) );
AOI211_X1 g_73_122 (.ZN (n_73_122), .A (n_77_120), .B (n_80_120), .C1 (n_84_118), .C2 (n_87_118) );
AOI211_X1 g_71_123 (.ZN (n_71_123), .A (n_75_121), .B (n_78_121), .C1 (n_82_119), .C2 (n_85_119) );
AOI211_X1 g_69_124 (.ZN (n_69_124), .A (n_73_122), .B (n_76_122), .C1 (n_80_120), .C2 (n_86_117) );
AOI211_X1 g_67_125 (.ZN (n_67_125), .A (n_71_123), .B (n_77_120), .C1 (n_78_121), .C2 (n_84_118) );
AOI211_X1 g_65_126 (.ZN (n_65_126), .A (n_69_124), .B (n_75_121), .C1 (n_76_122), .C2 (n_82_119) );
AOI211_X1 g_64_128 (.ZN (n_64_128), .A (n_67_125), .B (n_73_122), .C1 (n_77_120), .C2 (n_80_120) );
AOI211_X1 g_66_127 (.ZN (n_66_127), .A (n_65_126), .B (n_71_123), .C1 (n_75_121), .C2 (n_78_121) );
AOI211_X1 g_68_126 (.ZN (n_68_126), .A (n_64_128), .B (n_69_124), .C1 (n_73_122), .C2 (n_76_122) );
AOI211_X1 g_70_125 (.ZN (n_70_125), .A (n_66_127), .B (n_67_125), .C1 (n_71_123), .C2 (n_77_120) );
AOI211_X1 g_72_124 (.ZN (n_72_124), .A (n_68_126), .B (n_65_126), .C1 (n_69_124), .C2 (n_75_121) );
AOI211_X1 g_74_123 (.ZN (n_74_123), .A (n_70_125), .B (n_64_128), .C1 (n_67_125), .C2 (n_73_122) );
AOI211_X1 g_73_125 (.ZN (n_73_125), .A (n_72_124), .B (n_66_127), .C1 (n_65_126), .C2 (n_71_123) );
AOI211_X1 g_71_124 (.ZN (n_71_124), .A (n_74_123), .B (n_68_126), .C1 (n_64_128), .C2 (n_69_124) );
AOI211_X1 g_73_123 (.ZN (n_73_123), .A (n_73_125), .B (n_70_125), .C1 (n_66_127), .C2 (n_67_125) );
AOI211_X1 g_75_122 (.ZN (n_75_122), .A (n_71_124), .B (n_72_124), .C1 (n_68_126), .C2 (n_65_126) );
AOI211_X1 g_77_121 (.ZN (n_77_121), .A (n_73_123), .B (n_74_123), .C1 (n_70_125), .C2 (n_64_128) );
AOI211_X1 g_79_120 (.ZN (n_79_120), .A (n_75_122), .B (n_73_125), .C1 (n_72_124), .C2 (n_66_127) );
AOI211_X1 g_81_119 (.ZN (n_81_119), .A (n_77_121), .B (n_71_124), .C1 (n_74_123), .C2 (n_68_126) );
AOI211_X1 g_83_120 (.ZN (n_83_120), .A (n_79_120), .B (n_73_123), .C1 (n_73_125), .C2 (n_70_125) );
AOI211_X1 g_81_121 (.ZN (n_81_121), .A (n_81_119), .B (n_75_122), .C1 (n_71_124), .C2 (n_72_124) );
AOI211_X1 g_79_122 (.ZN (n_79_122), .A (n_83_120), .B (n_77_121), .C1 (n_73_123), .C2 (n_74_123) );
AOI211_X1 g_77_123 (.ZN (n_77_123), .A (n_81_121), .B (n_79_120), .C1 (n_75_122), .C2 (n_73_125) );
AOI211_X1 g_75_124 (.ZN (n_75_124), .A (n_79_122), .B (n_81_119), .C1 (n_77_121), .C2 (n_71_124) );
AOI211_X1 g_74_126 (.ZN (n_74_126), .A (n_77_123), .B (n_83_120), .C1 (n_79_120), .C2 (n_73_123) );
AOI211_X1 g_73_124 (.ZN (n_73_124), .A (n_75_124), .B (n_81_121), .C1 (n_81_119), .C2 (n_75_122) );
AOI211_X1 g_75_123 (.ZN (n_75_123), .A (n_74_126), .B (n_79_122), .C1 (n_83_120), .C2 (n_77_121) );
AOI211_X1 g_77_122 (.ZN (n_77_122), .A (n_73_124), .B (n_77_123), .C1 (n_81_121), .C2 (n_79_120) );
AOI211_X1 g_79_121 (.ZN (n_79_121), .A (n_75_123), .B (n_75_124), .C1 (n_79_122), .C2 (n_81_119) );
AOI211_X1 g_81_120 (.ZN (n_81_120), .A (n_77_122), .B (n_74_126), .C1 (n_77_123), .C2 (n_83_120) );
AOI211_X1 g_83_119 (.ZN (n_83_119), .A (n_79_121), .B (n_73_124), .C1 (n_75_124), .C2 (n_81_121) );
AOI211_X1 g_85_118 (.ZN (n_85_118), .A (n_81_120), .B (n_75_123), .C1 (n_74_126), .C2 (n_79_122) );
AOI211_X1 g_87_117 (.ZN (n_87_117), .A (n_83_119), .B (n_77_122), .C1 (n_73_124), .C2 (n_77_123) );
AOI211_X1 g_86_119 (.ZN (n_86_119), .A (n_85_118), .B (n_79_121), .C1 (n_75_123), .C2 (n_75_124) );
AOI211_X1 g_88_118 (.ZN (n_88_118), .A (n_87_117), .B (n_81_120), .C1 (n_77_122), .C2 (n_74_126) );
AOI211_X1 g_90_117 (.ZN (n_90_117), .A (n_86_119), .B (n_83_119), .C1 (n_79_121), .C2 (n_73_124) );
AOI211_X1 g_92_116 (.ZN (n_92_116), .A (n_88_118), .B (n_85_118), .C1 (n_81_120), .C2 (n_75_123) );
AOI211_X1 g_94_115 (.ZN (n_94_115), .A (n_90_117), .B (n_87_117), .C1 (n_83_119), .C2 (n_77_122) );
AOI211_X1 g_96_114 (.ZN (n_96_114), .A (n_92_116), .B (n_86_119), .C1 (n_85_118), .C2 (n_79_121) );
AOI211_X1 g_98_113 (.ZN (n_98_113), .A (n_94_115), .B (n_88_118), .C1 (n_87_117), .C2 (n_81_120) );
AOI211_X1 g_100_112 (.ZN (n_100_112), .A (n_96_114), .B (n_90_117), .C1 (n_86_119), .C2 (n_83_119) );
AOI211_X1 g_99_114 (.ZN (n_99_114), .A (n_98_113), .B (n_92_116), .C1 (n_88_118), .C2 (n_85_118) );
AOI211_X1 g_98_112 (.ZN (n_98_112), .A (n_100_112), .B (n_94_115), .C1 (n_90_117), .C2 (n_87_117) );
AOI211_X1 g_100_111 (.ZN (n_100_111), .A (n_99_114), .B (n_96_114), .C1 (n_92_116), .C2 (n_86_119) );
AOI211_X1 g_102_110 (.ZN (n_102_110), .A (n_98_112), .B (n_98_113), .C1 (n_94_115), .C2 (n_88_118) );
AOI211_X1 g_104_109 (.ZN (n_104_109), .A (n_100_111), .B (n_100_112), .C1 (n_96_114), .C2 (n_90_117) );
AOI211_X1 g_106_108 (.ZN (n_106_108), .A (n_102_110), .B (n_99_114), .C1 (n_98_113), .C2 (n_92_116) );
AOI211_X1 g_108_107 (.ZN (n_108_107), .A (n_104_109), .B (n_98_112), .C1 (n_100_112), .C2 (n_94_115) );
AOI211_X1 g_110_106 (.ZN (n_110_106), .A (n_106_108), .B (n_100_111), .C1 (n_99_114), .C2 (n_96_114) );
AOI211_X1 g_112_105 (.ZN (n_112_105), .A (n_108_107), .B (n_102_110), .C1 (n_98_112), .C2 (n_98_113) );
AOI211_X1 g_114_104 (.ZN (n_114_104), .A (n_110_106), .B (n_104_109), .C1 (n_100_111), .C2 (n_100_112) );
AOI211_X1 g_116_103 (.ZN (n_116_103), .A (n_112_105), .B (n_106_108), .C1 (n_102_110), .C2 (n_99_114) );
AOI211_X1 g_118_102 (.ZN (n_118_102), .A (n_114_104), .B (n_108_107), .C1 (n_104_109), .C2 (n_98_112) );
AOI211_X1 g_120_101 (.ZN (n_120_101), .A (n_116_103), .B (n_110_106), .C1 (n_106_108), .C2 (n_100_111) );
AOI211_X1 g_119_103 (.ZN (n_119_103), .A (n_118_102), .B (n_112_105), .C1 (n_108_107), .C2 (n_102_110) );
AOI211_X1 g_117_104 (.ZN (n_117_104), .A (n_120_101), .B (n_114_104), .C1 (n_110_106), .C2 (n_104_109) );
AOI211_X1 g_115_105 (.ZN (n_115_105), .A (n_119_103), .B (n_116_103), .C1 (n_112_105), .C2 (n_106_108) );
AOI211_X1 g_113_106 (.ZN (n_113_106), .A (n_117_104), .B (n_118_102), .C1 (n_114_104), .C2 (n_108_107) );
AOI211_X1 g_111_107 (.ZN (n_111_107), .A (n_115_105), .B (n_120_101), .C1 (n_116_103), .C2 (n_110_106) );
AOI211_X1 g_109_108 (.ZN (n_109_108), .A (n_113_106), .B (n_119_103), .C1 (n_118_102), .C2 (n_112_105) );
AOI211_X1 g_107_109 (.ZN (n_107_109), .A (n_111_107), .B (n_117_104), .C1 (n_120_101), .C2 (n_114_104) );
AOI211_X1 g_105_110 (.ZN (n_105_110), .A (n_109_108), .B (n_115_105), .C1 (n_119_103), .C2 (n_116_103) );
AOI211_X1 g_103_111 (.ZN (n_103_111), .A (n_107_109), .B (n_113_106), .C1 (n_117_104), .C2 (n_118_102) );
AOI211_X1 g_101_112 (.ZN (n_101_112), .A (n_105_110), .B (n_111_107), .C1 (n_115_105), .C2 (n_120_101) );
AOI211_X1 g_99_113 (.ZN (n_99_113), .A (n_103_111), .B (n_109_108), .C1 (n_113_106), .C2 (n_119_103) );
AOI211_X1 g_97_114 (.ZN (n_97_114), .A (n_101_112), .B (n_107_109), .C1 (n_111_107), .C2 (n_117_104) );
AOI211_X1 g_95_115 (.ZN (n_95_115), .A (n_99_113), .B (n_105_110), .C1 (n_109_108), .C2 (n_115_105) );
AOI211_X1 g_96_113 (.ZN (n_96_113), .A (n_97_114), .B (n_103_111), .C1 (n_107_109), .C2 (n_113_106) );
AOI211_X1 g_94_114 (.ZN (n_94_114), .A (n_95_115), .B (n_101_112), .C1 (n_105_110), .C2 (n_111_107) );
AOI211_X1 g_92_115 (.ZN (n_92_115), .A (n_96_113), .B (n_99_113), .C1 (n_103_111), .C2 (n_109_108) );
AOI211_X1 g_90_116 (.ZN (n_90_116), .A (n_94_114), .B (n_97_114), .C1 (n_101_112), .C2 (n_107_109) );
AOI211_X1 g_88_117 (.ZN (n_88_117), .A (n_92_115), .B (n_95_115), .C1 (n_99_113), .C2 (n_105_110) );
AOI211_X1 g_86_118 (.ZN (n_86_118), .A (n_90_116), .B (n_96_113), .C1 (n_97_114), .C2 (n_103_111) );
AOI211_X1 g_84_119 (.ZN (n_84_119), .A (n_88_117), .B (n_94_114), .C1 (n_95_115), .C2 (n_101_112) );
AOI211_X1 g_82_120 (.ZN (n_82_120), .A (n_86_118), .B (n_92_115), .C1 (n_96_113), .C2 (n_99_113) );
AOI211_X1 g_80_121 (.ZN (n_80_121), .A (n_84_119), .B (n_90_116), .C1 (n_94_114), .C2 (n_97_114) );
AOI211_X1 g_78_122 (.ZN (n_78_122), .A (n_82_120), .B (n_88_117), .C1 (n_92_115), .C2 (n_95_115) );
AOI211_X1 g_76_123 (.ZN (n_76_123), .A (n_80_121), .B (n_86_118), .C1 (n_90_116), .C2 (n_96_113) );
AOI211_X1 g_74_124 (.ZN (n_74_124), .A (n_78_122), .B (n_84_119), .C1 (n_88_117), .C2 (n_94_114) );
AOI211_X1 g_72_125 (.ZN (n_72_125), .A (n_76_123), .B (n_82_120), .C1 (n_86_118), .C2 (n_92_115) );
AOI211_X1 g_70_126 (.ZN (n_70_126), .A (n_74_124), .B (n_80_121), .C1 (n_84_119), .C2 (n_90_116) );
AOI211_X1 g_68_127 (.ZN (n_68_127), .A (n_72_125), .B (n_78_122), .C1 (n_82_120), .C2 (n_88_117) );
AOI211_X1 g_69_125 (.ZN (n_69_125), .A (n_70_126), .B (n_76_123), .C1 (n_80_121), .C2 (n_86_118) );
AOI211_X1 g_67_126 (.ZN (n_67_126), .A (n_68_127), .B (n_74_124), .C1 (n_78_122), .C2 (n_84_119) );
AOI211_X1 g_65_127 (.ZN (n_65_127), .A (n_69_125), .B (n_72_125), .C1 (n_76_123), .C2 (n_82_120) );
AOI211_X1 g_63_128 (.ZN (n_63_128), .A (n_67_126), .B (n_70_126), .C1 (n_74_124), .C2 (n_80_121) );
AOI211_X1 g_61_129 (.ZN (n_61_129), .A (n_65_127), .B (n_68_127), .C1 (n_72_125), .C2 (n_78_122) );
AOI211_X1 g_59_130 (.ZN (n_59_130), .A (n_63_128), .B (n_69_125), .C1 (n_70_126), .C2 (n_76_123) );
AOI211_X1 g_57_131 (.ZN (n_57_131), .A (n_61_129), .B (n_67_126), .C1 (n_68_127), .C2 (n_74_124) );
AOI211_X1 g_55_132 (.ZN (n_55_132), .A (n_59_130), .B (n_65_127), .C1 (n_69_125), .C2 (n_72_125) );
AOI211_X1 g_53_133 (.ZN (n_53_133), .A (n_57_131), .B (n_63_128), .C1 (n_67_126), .C2 (n_70_126) );
AOI211_X1 g_51_134 (.ZN (n_51_134), .A (n_55_132), .B (n_61_129), .C1 (n_65_127), .C2 (n_68_127) );
AOI211_X1 g_50_136 (.ZN (n_50_136), .A (n_53_133), .B (n_59_130), .C1 (n_63_128), .C2 (n_69_125) );
AOI211_X1 g_48_135 (.ZN (n_48_135), .A (n_51_134), .B (n_57_131), .C1 (n_61_129), .C2 (n_67_126) );
AOI211_X1 g_50_134 (.ZN (n_50_134), .A (n_50_136), .B (n_55_132), .C1 (n_59_130), .C2 (n_65_127) );
AOI211_X1 g_52_133 (.ZN (n_52_133), .A (n_48_135), .B (n_53_133), .C1 (n_57_131), .C2 (n_63_128) );
AOI211_X1 g_54_132 (.ZN (n_54_132), .A (n_50_134), .B (n_51_134), .C1 (n_55_132), .C2 (n_61_129) );
AOI211_X1 g_56_131 (.ZN (n_56_131), .A (n_52_133), .B (n_50_136), .C1 (n_53_133), .C2 (n_59_130) );
AOI211_X1 g_58_130 (.ZN (n_58_130), .A (n_54_132), .B (n_48_135), .C1 (n_51_134), .C2 (n_57_131) );
AOI211_X1 g_60_129 (.ZN (n_60_129), .A (n_56_131), .B (n_50_134), .C1 (n_50_136), .C2 (n_55_132) );
AOI211_X1 g_62_128 (.ZN (n_62_128), .A (n_58_130), .B (n_52_133), .C1 (n_48_135), .C2 (n_53_133) );
AOI211_X1 g_61_130 (.ZN (n_61_130), .A (n_60_129), .B (n_54_132), .C1 (n_50_134), .C2 (n_51_134) );
AOI211_X1 g_63_129 (.ZN (n_63_129), .A (n_62_128), .B (n_56_131), .C1 (n_52_133), .C2 (n_50_136) );
AOI211_X1 g_65_128 (.ZN (n_65_128), .A (n_61_130), .B (n_58_130), .C1 (n_54_132), .C2 (n_48_135) );
AOI211_X1 g_67_127 (.ZN (n_67_127), .A (n_63_129), .B (n_60_129), .C1 (n_56_131), .C2 (n_50_134) );
AOI211_X1 g_69_126 (.ZN (n_69_126), .A (n_65_128), .B (n_62_128), .C1 (n_58_130), .C2 (n_52_133) );
AOI211_X1 g_71_125 (.ZN (n_71_125), .A (n_67_127), .B (n_61_130), .C1 (n_60_129), .C2 (n_54_132) );
AOI211_X1 g_72_127 (.ZN (n_72_127), .A (n_69_126), .B (n_63_129), .C1 (n_62_128), .C2 (n_56_131) );
AOI211_X1 g_70_128 (.ZN (n_70_128), .A (n_71_125), .B (n_65_128), .C1 (n_61_130), .C2 (n_58_130) );
AOI211_X1 g_71_126 (.ZN (n_71_126), .A (n_72_127), .B (n_67_127), .C1 (n_63_129), .C2 (n_60_129) );
AOI211_X1 g_69_127 (.ZN (n_69_127), .A (n_70_128), .B (n_69_126), .C1 (n_65_128), .C2 (n_62_128) );
AOI211_X1 g_67_128 (.ZN (n_67_128), .A (n_71_126), .B (n_71_125), .C1 (n_67_127), .C2 (n_61_130) );
AOI211_X1 g_65_129 (.ZN (n_65_129), .A (n_69_127), .B (n_72_127), .C1 (n_69_126), .C2 (n_63_129) );
AOI211_X1 g_63_130 (.ZN (n_63_130), .A (n_67_128), .B (n_70_128), .C1 (n_71_125), .C2 (n_65_128) );
AOI211_X1 g_61_131 (.ZN (n_61_131), .A (n_65_129), .B (n_71_126), .C1 (n_72_127), .C2 (n_67_127) );
AOI211_X1 g_62_129 (.ZN (n_62_129), .A (n_63_130), .B (n_69_127), .C1 (n_70_128), .C2 (n_69_126) );
AOI211_X1 g_60_130 (.ZN (n_60_130), .A (n_61_131), .B (n_67_128), .C1 (n_71_126), .C2 (n_71_125) );
AOI211_X1 g_59_132 (.ZN (n_59_132), .A (n_62_129), .B (n_65_129), .C1 (n_69_127), .C2 (n_72_127) );
AOI211_X1 g_57_133 (.ZN (n_57_133), .A (n_60_130), .B (n_63_130), .C1 (n_67_128), .C2 (n_70_128) );
AOI211_X1 g_55_134 (.ZN (n_55_134), .A (n_59_132), .B (n_61_131), .C1 (n_65_129), .C2 (n_71_126) );
AOI211_X1 g_53_135 (.ZN (n_53_135), .A (n_57_133), .B (n_62_129), .C1 (n_63_130), .C2 (n_69_127) );
AOI211_X1 g_51_136 (.ZN (n_51_136), .A (n_55_134), .B (n_60_130), .C1 (n_61_131), .C2 (n_67_128) );
AOI211_X1 g_49_137 (.ZN (n_49_137), .A (n_53_135), .B (n_59_132), .C1 (n_62_129), .C2 (n_65_129) );
AOI211_X1 g_47_138 (.ZN (n_47_138), .A (n_51_136), .B (n_57_133), .C1 (n_60_130), .C2 (n_63_130) );
AOI211_X1 g_46_136 (.ZN (n_46_136), .A (n_49_137), .B (n_55_134), .C1 (n_59_132), .C2 (n_61_131) );
AOI211_X1 g_48_137 (.ZN (n_48_137), .A (n_47_138), .B (n_53_135), .C1 (n_57_133), .C2 (n_62_129) );
AOI211_X1 g_47_139 (.ZN (n_47_139), .A (n_46_136), .B (n_51_136), .C1 (n_55_134), .C2 (n_60_130) );
AOI211_X1 g_49_138 (.ZN (n_49_138), .A (n_48_137), .B (n_49_137), .C1 (n_53_135), .C2 (n_59_132) );
AOI211_X1 g_47_137 (.ZN (n_47_137), .A (n_47_139), .B (n_47_138), .C1 (n_51_136), .C2 (n_57_133) );
AOI211_X1 g_49_136 (.ZN (n_49_136), .A (n_49_138), .B (n_46_136), .C1 (n_49_137), .C2 (n_55_134) );
AOI211_X1 g_51_135 (.ZN (n_51_135), .A (n_47_137), .B (n_48_137), .C1 (n_47_138), .C2 (n_53_135) );
AOI211_X1 g_53_134 (.ZN (n_53_134), .A (n_49_136), .B (n_47_139), .C1 (n_46_136), .C2 (n_51_136) );
AOI211_X1 g_55_133 (.ZN (n_55_133), .A (n_51_135), .B (n_49_138), .C1 (n_48_137), .C2 (n_49_137) );
AOI211_X1 g_57_132 (.ZN (n_57_132), .A (n_53_134), .B (n_47_137), .C1 (n_47_139), .C2 (n_47_138) );
AOI211_X1 g_59_131 (.ZN (n_59_131), .A (n_55_133), .B (n_49_136), .C1 (n_49_138), .C2 (n_46_136) );
AOI211_X1 g_58_133 (.ZN (n_58_133), .A (n_57_132), .B (n_51_135), .C1 (n_47_137), .C2 (n_48_137) );
AOI211_X1 g_60_132 (.ZN (n_60_132), .A (n_59_131), .B (n_53_134), .C1 (n_49_136), .C2 (n_47_139) );
AOI211_X1 g_62_131 (.ZN (n_62_131), .A (n_58_133), .B (n_55_133), .C1 (n_51_135), .C2 (n_49_138) );
AOI211_X1 g_64_130 (.ZN (n_64_130), .A (n_60_132), .B (n_57_132), .C1 (n_53_134), .C2 (n_47_137) );
AOI211_X1 g_66_129 (.ZN (n_66_129), .A (n_62_131), .B (n_59_131), .C1 (n_55_133), .C2 (n_49_136) );
AOI211_X1 g_68_128 (.ZN (n_68_128), .A (n_64_130), .B (n_58_133), .C1 (n_57_132), .C2 (n_51_135) );
AOI211_X1 g_70_127 (.ZN (n_70_127), .A (n_66_129), .B (n_60_132), .C1 (n_59_131), .C2 (n_53_134) );
AOI211_X1 g_72_126 (.ZN (n_72_126), .A (n_68_128), .B (n_62_131), .C1 (n_58_133), .C2 (n_55_133) );
AOI211_X1 g_74_125 (.ZN (n_74_125), .A (n_70_127), .B (n_64_130), .C1 (n_60_132), .C2 (n_57_132) );
AOI211_X1 g_76_124 (.ZN (n_76_124), .A (n_72_126), .B (n_66_129), .C1 (n_62_131), .C2 (n_59_131) );
AOI211_X1 g_78_123 (.ZN (n_78_123), .A (n_74_125), .B (n_68_128), .C1 (n_64_130), .C2 (n_58_133) );
AOI211_X1 g_80_122 (.ZN (n_80_122), .A (n_76_124), .B (n_70_127), .C1 (n_66_129), .C2 (n_60_132) );
AOI211_X1 g_82_121 (.ZN (n_82_121), .A (n_78_123), .B (n_72_126), .C1 (n_68_128), .C2 (n_62_131) );
AOI211_X1 g_84_120 (.ZN (n_84_120), .A (n_80_122), .B (n_74_125), .C1 (n_70_127), .C2 (n_64_130) );
AOI211_X1 g_83_122 (.ZN (n_83_122), .A (n_82_121), .B (n_76_124), .C1 (n_72_126), .C2 (n_66_129) );
AOI211_X1 g_85_121 (.ZN (n_85_121), .A (n_84_120), .B (n_78_123), .C1 (n_74_125), .C2 (n_68_128) );
AOI211_X1 g_87_120 (.ZN (n_87_120), .A (n_83_122), .B (n_80_122), .C1 (n_76_124), .C2 (n_70_127) );
AOI211_X1 g_89_119 (.ZN (n_89_119), .A (n_85_121), .B (n_82_121), .C1 (n_78_123), .C2 (n_72_126) );
AOI211_X1 g_91_118 (.ZN (n_91_118), .A (n_87_120), .B (n_84_120), .C1 (n_80_122), .C2 (n_74_125) );
AOI211_X1 g_93_117 (.ZN (n_93_117), .A (n_89_119), .B (n_83_122), .C1 (n_82_121), .C2 (n_76_124) );
AOI211_X1 g_91_116 (.ZN (n_91_116), .A (n_91_118), .B (n_85_121), .C1 (n_84_120), .C2 (n_78_123) );
AOI211_X1 g_93_115 (.ZN (n_93_115), .A (n_93_117), .B (n_87_120), .C1 (n_83_122), .C2 (n_80_122) );
AOI211_X1 g_95_114 (.ZN (n_95_114), .A (n_91_116), .B (n_89_119), .C1 (n_85_121), .C2 (n_82_121) );
AOI211_X1 g_97_113 (.ZN (n_97_113), .A (n_93_115), .B (n_91_118), .C1 (n_87_120), .C2 (n_84_120) );
AOI211_X1 g_99_112 (.ZN (n_99_112), .A (n_95_114), .B (n_93_117), .C1 (n_89_119), .C2 (n_83_122) );
AOI211_X1 g_101_111 (.ZN (n_101_111), .A (n_97_113), .B (n_91_116), .C1 (n_91_118), .C2 (n_85_121) );
AOI211_X1 g_103_110 (.ZN (n_103_110), .A (n_99_112), .B (n_93_115), .C1 (n_93_117), .C2 (n_87_120) );
AOI211_X1 g_105_109 (.ZN (n_105_109), .A (n_101_111), .B (n_95_114), .C1 (n_91_116), .C2 (n_89_119) );
AOI211_X1 g_107_108 (.ZN (n_107_108), .A (n_103_110), .B (n_97_113), .C1 (n_93_115), .C2 (n_91_118) );
AOI211_X1 g_109_107 (.ZN (n_109_107), .A (n_105_109), .B (n_99_112), .C1 (n_95_114), .C2 (n_93_117) );
AOI211_X1 g_111_106 (.ZN (n_111_106), .A (n_107_108), .B (n_101_111), .C1 (n_97_113), .C2 (n_91_116) );
AOI211_X1 g_113_105 (.ZN (n_113_105), .A (n_109_107), .B (n_103_110), .C1 (n_99_112), .C2 (n_93_115) );
AOI211_X1 g_115_104 (.ZN (n_115_104), .A (n_111_106), .B (n_105_109), .C1 (n_101_111), .C2 (n_95_114) );
AOI211_X1 g_117_103 (.ZN (n_117_103), .A (n_113_105), .B (n_107_108), .C1 (n_103_110), .C2 (n_97_113) );
AOI211_X1 g_119_102 (.ZN (n_119_102), .A (n_115_104), .B (n_109_107), .C1 (n_105_109), .C2 (n_99_112) );
AOI211_X1 g_120_104 (.ZN (n_120_104), .A (n_117_103), .B (n_111_106), .C1 (n_107_108), .C2 (n_101_111) );
AOI211_X1 g_118_105 (.ZN (n_118_105), .A (n_119_102), .B (n_113_105), .C1 (n_109_107), .C2 (n_103_110) );
AOI211_X1 g_116_106 (.ZN (n_116_106), .A (n_120_104), .B (n_115_104), .C1 (n_111_106), .C2 (n_105_109) );
AOI211_X1 g_114_107 (.ZN (n_114_107), .A (n_118_105), .B (n_117_103), .C1 (n_113_105), .C2 (n_107_108) );
AOI211_X1 g_112_108 (.ZN (n_112_108), .A (n_116_106), .B (n_119_102), .C1 (n_115_104), .C2 (n_109_107) );
AOI211_X1 g_110_109 (.ZN (n_110_109), .A (n_114_107), .B (n_120_104), .C1 (n_117_103), .C2 (n_111_106) );
AOI211_X1 g_108_110 (.ZN (n_108_110), .A (n_112_108), .B (n_118_105), .C1 (n_119_102), .C2 (n_113_105) );
AOI211_X1 g_106_111 (.ZN (n_106_111), .A (n_110_109), .B (n_116_106), .C1 (n_120_104), .C2 (n_115_104) );
AOI211_X1 g_104_112 (.ZN (n_104_112), .A (n_108_110), .B (n_114_107), .C1 (n_118_105), .C2 (n_117_103) );
AOI211_X1 g_102_113 (.ZN (n_102_113), .A (n_106_111), .B (n_112_108), .C1 (n_116_106), .C2 (n_119_102) );
AOI211_X1 g_100_114 (.ZN (n_100_114), .A (n_104_112), .B (n_110_109), .C1 (n_114_107), .C2 (n_120_104) );
AOI211_X1 g_98_115 (.ZN (n_98_115), .A (n_102_113), .B (n_108_110), .C1 (n_112_108), .C2 (n_118_105) );
AOI211_X1 g_96_116 (.ZN (n_96_116), .A (n_100_114), .B (n_106_111), .C1 (n_110_109), .C2 (n_116_106) );
AOI211_X1 g_94_117 (.ZN (n_94_117), .A (n_98_115), .B (n_104_112), .C1 (n_108_110), .C2 (n_114_107) );
AOI211_X1 g_92_118 (.ZN (n_92_118), .A (n_96_116), .B (n_102_113), .C1 (n_106_111), .C2 (n_112_108) );
AOI211_X1 g_93_116 (.ZN (n_93_116), .A (n_94_117), .B (n_100_114), .C1 (n_104_112), .C2 (n_110_109) );
AOI211_X1 g_91_117 (.ZN (n_91_117), .A (n_92_118), .B (n_98_115), .C1 (n_102_113), .C2 (n_108_110) );
AOI211_X1 g_89_118 (.ZN (n_89_118), .A (n_93_116), .B (n_96_116), .C1 (n_100_114), .C2 (n_106_111) );
AOI211_X1 g_87_119 (.ZN (n_87_119), .A (n_91_117), .B (n_94_117), .C1 (n_98_115), .C2 (n_104_112) );
AOI211_X1 g_85_120 (.ZN (n_85_120), .A (n_89_118), .B (n_92_118), .C1 (n_96_116), .C2 (n_102_113) );
AOI211_X1 g_83_121 (.ZN (n_83_121), .A (n_87_119), .B (n_93_116), .C1 (n_94_117), .C2 (n_100_114) );
AOI211_X1 g_81_122 (.ZN (n_81_122), .A (n_85_120), .B (n_91_117), .C1 (n_92_118), .C2 (n_98_115) );
AOI211_X1 g_79_123 (.ZN (n_79_123), .A (n_83_121), .B (n_89_118), .C1 (n_93_116), .C2 (n_96_116) );
AOI211_X1 g_77_124 (.ZN (n_77_124), .A (n_81_122), .B (n_87_119), .C1 (n_91_117), .C2 (n_94_117) );
AOI211_X1 g_75_125 (.ZN (n_75_125), .A (n_79_123), .B (n_85_120), .C1 (n_89_118), .C2 (n_92_118) );
AOI211_X1 g_73_126 (.ZN (n_73_126), .A (n_77_124), .B (n_83_121), .C1 (n_87_119), .C2 (n_93_116) );
AOI211_X1 g_71_127 (.ZN (n_71_127), .A (n_75_125), .B (n_81_122), .C1 (n_85_120), .C2 (n_91_117) );
AOI211_X1 g_69_128 (.ZN (n_69_128), .A (n_73_126), .B (n_79_123), .C1 (n_83_121), .C2 (n_89_118) );
AOI211_X1 g_67_129 (.ZN (n_67_129), .A (n_71_127), .B (n_77_124), .C1 (n_81_122), .C2 (n_87_119) );
AOI211_X1 g_65_130 (.ZN (n_65_130), .A (n_69_128), .B (n_75_125), .C1 (n_79_123), .C2 (n_85_120) );
AOI211_X1 g_66_128 (.ZN (n_66_128), .A (n_67_129), .B (n_73_126), .C1 (n_77_124), .C2 (n_83_121) );
AOI211_X1 g_64_129 (.ZN (n_64_129), .A (n_65_130), .B (n_71_127), .C1 (n_75_125), .C2 (n_81_122) );
AOI211_X1 g_62_130 (.ZN (n_62_130), .A (n_66_128), .B (n_69_128), .C1 (n_73_126), .C2 (n_79_123) );
AOI211_X1 g_60_131 (.ZN (n_60_131), .A (n_64_129), .B (n_67_129), .C1 (n_71_127), .C2 (n_77_124) );
AOI211_X1 g_58_132 (.ZN (n_58_132), .A (n_62_130), .B (n_65_130), .C1 (n_69_128), .C2 (n_75_125) );
AOI211_X1 g_56_133 (.ZN (n_56_133), .A (n_60_131), .B (n_66_128), .C1 (n_67_129), .C2 (n_73_126) );
AOI211_X1 g_54_134 (.ZN (n_54_134), .A (n_58_132), .B (n_64_129), .C1 (n_65_130), .C2 (n_71_127) );
AOI211_X1 g_52_135 (.ZN (n_52_135), .A (n_56_133), .B (n_62_130), .C1 (n_66_128), .C2 (n_69_128) );
AOI211_X1 g_51_137 (.ZN (n_51_137), .A (n_54_134), .B (n_60_131), .C1 (n_64_129), .C2 (n_67_129) );
AOI211_X1 g_53_136 (.ZN (n_53_136), .A (n_52_135), .B (n_58_132), .C1 (n_62_130), .C2 (n_65_130) );
AOI211_X1 g_55_135 (.ZN (n_55_135), .A (n_51_137), .B (n_56_133), .C1 (n_60_131), .C2 (n_66_128) );
AOI211_X1 g_57_134 (.ZN (n_57_134), .A (n_53_136), .B (n_54_134), .C1 (n_58_132), .C2 (n_64_129) );
AOI211_X1 g_59_133 (.ZN (n_59_133), .A (n_55_135), .B (n_52_135), .C1 (n_56_133), .C2 (n_62_130) );
AOI211_X1 g_61_132 (.ZN (n_61_132), .A (n_57_134), .B (n_51_137), .C1 (n_54_134), .C2 (n_60_131) );
AOI211_X1 g_63_131 (.ZN (n_63_131), .A (n_59_133), .B (n_53_136), .C1 (n_52_135), .C2 (n_58_132) );
AOI211_X1 g_62_133 (.ZN (n_62_133), .A (n_61_132), .B (n_55_135), .C1 (n_51_137), .C2 (n_56_133) );
AOI211_X1 g_64_132 (.ZN (n_64_132), .A (n_63_131), .B (n_57_134), .C1 (n_53_136), .C2 (n_54_134) );
AOI211_X1 g_66_131 (.ZN (n_66_131), .A (n_62_133), .B (n_59_133), .C1 (n_55_135), .C2 (n_52_135) );
AOI211_X1 g_68_130 (.ZN (n_68_130), .A (n_64_132), .B (n_61_132), .C1 (n_57_134), .C2 (n_51_137) );
AOI211_X1 g_70_129 (.ZN (n_70_129), .A (n_66_131), .B (n_63_131), .C1 (n_59_133), .C2 (n_53_136) );
AOI211_X1 g_72_128 (.ZN (n_72_128), .A (n_68_130), .B (n_62_133), .C1 (n_61_132), .C2 (n_55_135) );
AOI211_X1 g_74_127 (.ZN (n_74_127), .A (n_70_129), .B (n_64_132), .C1 (n_63_131), .C2 (n_57_134) );
AOI211_X1 g_76_126 (.ZN (n_76_126), .A (n_72_128), .B (n_66_131), .C1 (n_62_133), .C2 (n_59_133) );
AOI211_X1 g_78_125 (.ZN (n_78_125), .A (n_74_127), .B (n_68_130), .C1 (n_64_132), .C2 (n_61_132) );
AOI211_X1 g_80_124 (.ZN (n_80_124), .A (n_76_126), .B (n_70_129), .C1 (n_66_131), .C2 (n_63_131) );
AOI211_X1 g_82_123 (.ZN (n_82_123), .A (n_78_125), .B (n_72_128), .C1 (n_68_130), .C2 (n_62_133) );
AOI211_X1 g_84_122 (.ZN (n_84_122), .A (n_80_124), .B (n_74_127), .C1 (n_70_129), .C2 (n_64_132) );
AOI211_X1 g_86_121 (.ZN (n_86_121), .A (n_82_123), .B (n_76_126), .C1 (n_72_128), .C2 (n_66_131) );
AOI211_X1 g_88_120 (.ZN (n_88_120), .A (n_84_122), .B (n_78_125), .C1 (n_74_127), .C2 (n_68_130) );
AOI211_X1 g_90_119 (.ZN (n_90_119), .A (n_86_121), .B (n_80_124), .C1 (n_76_126), .C2 (n_70_129) );
AOI211_X1 g_89_121 (.ZN (n_89_121), .A (n_88_120), .B (n_82_123), .C1 (n_78_125), .C2 (n_72_128) );
AOI211_X1 g_88_119 (.ZN (n_88_119), .A (n_90_119), .B (n_84_122), .C1 (n_80_124), .C2 (n_74_127) );
AOI211_X1 g_90_118 (.ZN (n_90_118), .A (n_89_121), .B (n_86_121), .C1 (n_82_123), .C2 (n_76_126) );
AOI211_X1 g_92_117 (.ZN (n_92_117), .A (n_88_119), .B (n_88_120), .C1 (n_84_122), .C2 (n_78_125) );
AOI211_X1 g_94_116 (.ZN (n_94_116), .A (n_90_118), .B (n_90_119), .C1 (n_86_121), .C2 (n_80_124) );
AOI211_X1 g_96_115 (.ZN (n_96_115), .A (n_92_117), .B (n_89_121), .C1 (n_88_120), .C2 (n_82_123) );
AOI211_X1 g_98_114 (.ZN (n_98_114), .A (n_94_116), .B (n_88_119), .C1 (n_90_119), .C2 (n_84_122) );
AOI211_X1 g_100_113 (.ZN (n_100_113), .A (n_96_115), .B (n_90_118), .C1 (n_89_121), .C2 (n_86_121) );
AOI211_X1 g_102_112 (.ZN (n_102_112), .A (n_98_114), .B (n_92_117), .C1 (n_88_119), .C2 (n_88_120) );
AOI211_X1 g_104_111 (.ZN (n_104_111), .A (n_100_113), .B (n_94_116), .C1 (n_90_118), .C2 (n_90_119) );
AOI211_X1 g_106_110 (.ZN (n_106_110), .A (n_102_112), .B (n_96_115), .C1 (n_92_117), .C2 (n_89_121) );
AOI211_X1 g_108_109 (.ZN (n_108_109), .A (n_104_111), .B (n_98_114), .C1 (n_94_116), .C2 (n_88_119) );
AOI211_X1 g_110_108 (.ZN (n_110_108), .A (n_106_110), .B (n_100_113), .C1 (n_96_115), .C2 (n_90_118) );
AOI211_X1 g_112_107 (.ZN (n_112_107), .A (n_108_109), .B (n_102_112), .C1 (n_98_114), .C2 (n_92_117) );
AOI211_X1 g_114_106 (.ZN (n_114_106), .A (n_110_108), .B (n_104_111), .C1 (n_100_113), .C2 (n_94_116) );
AOI211_X1 g_116_105 (.ZN (n_116_105), .A (n_112_107), .B (n_106_110), .C1 (n_102_112), .C2 (n_96_115) );
AOI211_X1 g_118_104 (.ZN (n_118_104), .A (n_114_106), .B (n_108_109), .C1 (n_104_111), .C2 (n_98_114) );
AOI211_X1 g_120_103 (.ZN (n_120_103), .A (n_116_105), .B (n_110_108), .C1 (n_106_110), .C2 (n_100_113) );
AOI211_X1 g_122_102 (.ZN (n_122_102), .A (n_118_104), .B (n_112_107), .C1 (n_108_109), .C2 (n_102_112) );
AOI211_X1 g_121_104 (.ZN (n_121_104), .A (n_120_103), .B (n_114_106), .C1 (n_110_108), .C2 (n_104_111) );
AOI211_X1 g_119_105 (.ZN (n_119_105), .A (n_122_102), .B (n_116_105), .C1 (n_112_107), .C2 (n_106_110) );
AOI211_X1 g_117_106 (.ZN (n_117_106), .A (n_121_104), .B (n_118_104), .C1 (n_114_106), .C2 (n_108_109) );
AOI211_X1 g_115_107 (.ZN (n_115_107), .A (n_119_105), .B (n_120_103), .C1 (n_116_105), .C2 (n_110_108) );
AOI211_X1 g_113_108 (.ZN (n_113_108), .A (n_117_106), .B (n_122_102), .C1 (n_118_104), .C2 (n_112_107) );
AOI211_X1 g_111_109 (.ZN (n_111_109), .A (n_115_107), .B (n_121_104), .C1 (n_120_103), .C2 (n_114_106) );
AOI211_X1 g_109_110 (.ZN (n_109_110), .A (n_113_108), .B (n_119_105), .C1 (n_122_102), .C2 (n_116_105) );
AOI211_X1 g_107_111 (.ZN (n_107_111), .A (n_111_109), .B (n_117_106), .C1 (n_121_104), .C2 (n_118_104) );
AOI211_X1 g_105_112 (.ZN (n_105_112), .A (n_109_110), .B (n_115_107), .C1 (n_119_105), .C2 (n_120_103) );
AOI211_X1 g_103_113 (.ZN (n_103_113), .A (n_107_111), .B (n_113_108), .C1 (n_117_106), .C2 (n_122_102) );
AOI211_X1 g_101_114 (.ZN (n_101_114), .A (n_105_112), .B (n_111_109), .C1 (n_115_107), .C2 (n_121_104) );
AOI211_X1 g_99_115 (.ZN (n_99_115), .A (n_103_113), .B (n_109_110), .C1 (n_113_108), .C2 (n_119_105) );
AOI211_X1 g_97_116 (.ZN (n_97_116), .A (n_101_114), .B (n_107_111), .C1 (n_111_109), .C2 (n_117_106) );
AOI211_X1 g_95_117 (.ZN (n_95_117), .A (n_99_115), .B (n_105_112), .C1 (n_109_110), .C2 (n_115_107) );
AOI211_X1 g_93_118 (.ZN (n_93_118), .A (n_97_116), .B (n_103_113), .C1 (n_107_111), .C2 (n_113_108) );
AOI211_X1 g_91_119 (.ZN (n_91_119), .A (n_95_117), .B (n_101_114), .C1 (n_105_112), .C2 (n_111_109) );
AOI211_X1 g_89_120 (.ZN (n_89_120), .A (n_93_118), .B (n_99_115), .C1 (n_103_113), .C2 (n_109_110) );
AOI211_X1 g_87_121 (.ZN (n_87_121), .A (n_91_119), .B (n_97_116), .C1 (n_101_114), .C2 (n_107_111) );
AOI211_X1 g_85_122 (.ZN (n_85_122), .A (n_89_120), .B (n_95_117), .C1 (n_99_115), .C2 (n_105_112) );
AOI211_X1 g_86_120 (.ZN (n_86_120), .A (n_87_121), .B (n_93_118), .C1 (n_97_116), .C2 (n_103_113) );
AOI211_X1 g_84_121 (.ZN (n_84_121), .A (n_85_122), .B (n_91_119), .C1 (n_95_117), .C2 (n_101_114) );
AOI211_X1 g_82_122 (.ZN (n_82_122), .A (n_86_120), .B (n_89_120), .C1 (n_93_118), .C2 (n_99_115) );
AOI211_X1 g_80_123 (.ZN (n_80_123), .A (n_84_121), .B (n_87_121), .C1 (n_91_119), .C2 (n_97_116) );
AOI211_X1 g_78_124 (.ZN (n_78_124), .A (n_82_122), .B (n_85_122), .C1 (n_89_120), .C2 (n_95_117) );
AOI211_X1 g_76_125 (.ZN (n_76_125), .A (n_80_123), .B (n_86_120), .C1 (n_87_121), .C2 (n_93_118) );
AOI211_X1 g_75_127 (.ZN (n_75_127), .A (n_78_124), .B (n_84_121), .C1 (n_85_122), .C2 (n_91_119) );
AOI211_X1 g_77_126 (.ZN (n_77_126), .A (n_76_125), .B (n_82_122), .C1 (n_86_120), .C2 (n_89_120) );
AOI211_X1 g_79_125 (.ZN (n_79_125), .A (n_75_127), .B (n_80_123), .C1 (n_84_121), .C2 (n_87_121) );
AOI211_X1 g_81_124 (.ZN (n_81_124), .A (n_77_126), .B (n_78_124), .C1 (n_82_122), .C2 (n_85_122) );
AOI211_X1 g_83_123 (.ZN (n_83_123), .A (n_79_125), .B (n_76_125), .C1 (n_80_123), .C2 (n_86_120) );
AOI211_X1 g_82_125 (.ZN (n_82_125), .A (n_81_124), .B (n_75_127), .C1 (n_78_124), .C2 (n_84_121) );
AOI211_X1 g_81_123 (.ZN (n_81_123), .A (n_83_123), .B (n_77_126), .C1 (n_76_125), .C2 (n_82_122) );
AOI211_X1 g_79_124 (.ZN (n_79_124), .A (n_82_125), .B (n_79_125), .C1 (n_75_127), .C2 (n_80_123) );
AOI211_X1 g_77_125 (.ZN (n_77_125), .A (n_81_123), .B (n_81_124), .C1 (n_77_126), .C2 (n_78_124) );
AOI211_X1 g_75_126 (.ZN (n_75_126), .A (n_79_124), .B (n_83_123), .C1 (n_79_125), .C2 (n_76_125) );
AOI211_X1 g_73_127 (.ZN (n_73_127), .A (n_77_125), .B (n_82_125), .C1 (n_81_124), .C2 (n_75_127) );
AOI211_X1 g_71_128 (.ZN (n_71_128), .A (n_75_126), .B (n_81_123), .C1 (n_83_123), .C2 (n_77_126) );
AOI211_X1 g_69_129 (.ZN (n_69_129), .A (n_73_127), .B (n_79_124), .C1 (n_82_125), .C2 (n_79_125) );
AOI211_X1 g_67_130 (.ZN (n_67_130), .A (n_71_128), .B (n_77_125), .C1 (n_81_123), .C2 (n_81_124) );
AOI211_X1 g_65_131 (.ZN (n_65_131), .A (n_69_129), .B (n_75_126), .C1 (n_79_124), .C2 (n_83_123) );
AOI211_X1 g_63_132 (.ZN (n_63_132), .A (n_67_130), .B (n_73_127), .C1 (n_77_125), .C2 (n_82_125) );
AOI211_X1 g_61_133 (.ZN (n_61_133), .A (n_65_131), .B (n_71_128), .C1 (n_75_126), .C2 (n_81_123) );
AOI211_X1 g_59_134 (.ZN (n_59_134), .A (n_63_132), .B (n_69_129), .C1 (n_73_127), .C2 (n_79_124) );
AOI211_X1 g_57_135 (.ZN (n_57_135), .A (n_61_133), .B (n_67_130), .C1 (n_71_128), .C2 (n_77_125) );
AOI211_X1 g_55_136 (.ZN (n_55_136), .A (n_59_134), .B (n_65_131), .C1 (n_69_129), .C2 (n_75_126) );
AOI211_X1 g_56_134 (.ZN (n_56_134), .A (n_57_135), .B (n_63_132), .C1 (n_67_130), .C2 (n_73_127) );
AOI211_X1 g_54_135 (.ZN (n_54_135), .A (n_55_136), .B (n_61_133), .C1 (n_65_131), .C2 (n_71_128) );
AOI211_X1 g_52_136 (.ZN (n_52_136), .A (n_56_134), .B (n_59_134), .C1 (n_63_132), .C2 (n_69_129) );
AOI211_X1 g_50_137 (.ZN (n_50_137), .A (n_54_135), .B (n_57_135), .C1 (n_61_133), .C2 (n_67_130) );
AOI211_X1 g_48_138 (.ZN (n_48_138), .A (n_52_136), .B (n_55_136), .C1 (n_59_134), .C2 (n_65_131) );
AOI211_X1 g_46_139 (.ZN (n_46_139), .A (n_50_137), .B (n_56_134), .C1 (n_57_135), .C2 (n_63_132) );
AOI211_X1 g_44_138 (.ZN (n_44_138), .A (n_48_138), .B (n_54_135), .C1 (n_55_136), .C2 (n_61_133) );
AOI211_X1 g_45_140 (.ZN (n_45_140), .A (n_46_139), .B (n_52_136), .C1 (n_56_134), .C2 (n_59_134) );
AOI211_X1 g_43_139 (.ZN (n_43_139), .A (n_44_138), .B (n_50_137), .C1 (n_54_135), .C2 (n_57_135) );
AOI211_X1 g_45_138 (.ZN (n_45_138), .A (n_45_140), .B (n_48_138), .C1 (n_52_136), .C2 (n_55_136) );
AOI211_X1 g_43_137 (.ZN (n_43_137), .A (n_43_139), .B (n_46_139), .C1 (n_50_137), .C2 (n_56_134) );
AOI211_X1 g_41_138 (.ZN (n_41_138), .A (n_45_138), .B (n_44_138), .C1 (n_48_138), .C2 (n_54_135) );
AOI211_X1 g_42_136 (.ZN (n_42_136), .A (n_43_137), .B (n_45_140), .C1 (n_46_139), .C2 (n_52_136) );
AOI211_X1 g_44_137 (.ZN (n_44_137), .A (n_41_138), .B (n_43_139), .C1 (n_44_138), .C2 (n_50_137) );
AOI211_X1 g_42_138 (.ZN (n_42_138), .A (n_42_136), .B (n_45_138), .C1 (n_45_140), .C2 (n_48_138) );
AOI211_X1 g_40_137 (.ZN (n_40_137), .A (n_44_137), .B (n_43_137), .C1 (n_43_139), .C2 (n_46_139) );
AOI211_X1 g_38_138 (.ZN (n_38_138), .A (n_42_138), .B (n_41_138), .C1 (n_45_138), .C2 (n_44_138) );
AOI211_X1 g_36_139 (.ZN (n_36_139), .A (n_40_137), .B (n_42_136), .C1 (n_43_137), .C2 (n_45_140) );
AOI211_X1 g_34_140 (.ZN (n_34_140), .A (n_38_138), .B (n_44_137), .C1 (n_41_138), .C2 (n_43_139) );
AOI211_X1 g_32_141 (.ZN (n_32_141), .A (n_36_139), .B (n_42_138), .C1 (n_42_136), .C2 (n_45_138) );
AOI211_X1 g_30_142 (.ZN (n_30_142), .A (n_34_140), .B (n_40_137), .C1 (n_44_137), .C2 (n_43_137) );
AOI211_X1 g_28_143 (.ZN (n_28_143), .A (n_32_141), .B (n_38_138), .C1 (n_42_138), .C2 (n_41_138) );
AOI211_X1 g_27_145 (.ZN (n_27_145), .A (n_30_142), .B (n_36_139), .C1 (n_40_137), .C2 (n_42_136) );
AOI211_X1 g_25_146 (.ZN (n_25_146), .A (n_28_143), .B (n_34_140), .C1 (n_38_138), .C2 (n_44_137) );
AOI211_X1 g_23_147 (.ZN (n_23_147), .A (n_27_145), .B (n_32_141), .C1 (n_36_139), .C2 (n_42_138) );
AOI211_X1 g_24_145 (.ZN (n_24_145), .A (n_25_146), .B (n_30_142), .C1 (n_34_140), .C2 (n_40_137) );
AOI211_X1 g_25_147 (.ZN (n_25_147), .A (n_23_147), .B (n_28_143), .C1 (n_32_141), .C2 (n_38_138) );
AOI211_X1 g_23_146 (.ZN (n_23_146), .A (n_24_145), .B (n_27_145), .C1 (n_30_142), .C2 (n_36_139) );
AOI211_X1 g_22_148 (.ZN (n_22_148), .A (n_25_147), .B (n_25_146), .C1 (n_28_143), .C2 (n_34_140) );
AOI211_X1 g_24_149 (.ZN (n_24_149), .A (n_23_146), .B (n_23_147), .C1 (n_27_145), .C2 (n_32_141) );
AOI211_X1 g_26_150 (.ZN (n_26_150), .A (n_22_148), .B (n_24_145), .C1 (n_25_146), .C2 (n_30_142) );
AOI211_X1 g_25_148 (.ZN (n_25_148), .A (n_24_149), .B (n_25_147), .C1 (n_23_147), .C2 (n_28_143) );
AOI211_X1 g_27_147 (.ZN (n_27_147), .A (n_26_150), .B (n_23_146), .C1 (n_24_145), .C2 (n_27_145) );
AOI211_X1 g_29_146 (.ZN (n_29_146), .A (n_25_148), .B (n_22_148), .C1 (n_25_147), .C2 (n_25_146) );
AOI211_X1 g_31_145 (.ZN (n_31_145), .A (n_27_147), .B (n_24_149), .C1 (n_23_146), .C2 (n_23_147) );
AOI211_X1 g_29_144 (.ZN (n_29_144), .A (n_29_146), .B (n_26_150), .C1 (n_22_148), .C2 (n_24_145) );
AOI211_X1 g_31_143 (.ZN (n_31_143), .A (n_31_145), .B (n_25_148), .C1 (n_24_149), .C2 (n_25_147) );
AOI211_X1 g_33_142 (.ZN (n_33_142), .A (n_29_144), .B (n_27_147), .C1 (n_26_150), .C2 (n_23_146) );
AOI211_X1 g_35_141 (.ZN (n_35_141), .A (n_31_143), .B (n_29_146), .C1 (n_25_148), .C2 (n_22_148) );
AOI211_X1 g_37_140 (.ZN (n_37_140), .A (n_33_142), .B (n_31_145), .C1 (n_27_147), .C2 (n_24_149) );
AOI211_X1 g_39_139 (.ZN (n_39_139), .A (n_35_141), .B (n_29_144), .C1 (n_29_146), .C2 (n_26_150) );
AOI211_X1 g_41_140 (.ZN (n_41_140), .A (n_37_140), .B (n_31_143), .C1 (n_31_145), .C2 (n_25_148) );
AOI211_X1 g_39_141 (.ZN (n_39_141), .A (n_39_139), .B (n_33_142), .C1 (n_29_144), .C2 (n_27_147) );
AOI211_X1 g_40_139 (.ZN (n_40_139), .A (n_41_140), .B (n_35_141), .C1 (n_31_143), .C2 (n_29_146) );
AOI211_X1 g_41_137 (.ZN (n_41_137), .A (n_39_141), .B (n_37_140), .C1 (n_33_142), .C2 (n_31_145) );
AOI211_X1 g_39_138 (.ZN (n_39_138), .A (n_40_139), .B (n_39_139), .C1 (n_35_141), .C2 (n_29_144) );
AOI211_X1 g_37_139 (.ZN (n_37_139), .A (n_41_137), .B (n_41_140), .C1 (n_37_140), .C2 (n_31_143) );
AOI211_X1 g_35_140 (.ZN (n_35_140), .A (n_39_138), .B (n_39_141), .C1 (n_39_139), .C2 (n_33_142) );
AOI211_X1 g_33_141 (.ZN (n_33_141), .A (n_37_139), .B (n_40_139), .C1 (n_41_140), .C2 (n_35_141) );
AOI211_X1 g_31_142 (.ZN (n_31_142), .A (n_35_140), .B (n_41_137), .C1 (n_39_141), .C2 (n_37_140) );
AOI211_X1 g_29_143 (.ZN (n_29_143), .A (n_33_141), .B (n_39_138), .C1 (n_40_139), .C2 (n_39_139) );
AOI211_X1 g_27_144 (.ZN (n_27_144), .A (n_31_142), .B (n_37_139), .C1 (n_41_137), .C2 (n_41_140) );
AOI211_X1 g_25_145 (.ZN (n_25_145), .A (n_29_143), .B (n_35_140), .C1 (n_39_138), .C2 (n_39_141) );
AOI211_X1 g_24_147 (.ZN (n_24_147), .A (n_27_144), .B (n_33_141), .C1 (n_37_139), .C2 (n_40_139) );
AOI211_X1 g_26_146 (.ZN (n_26_146), .A (n_25_145), .B (n_31_142), .C1 (n_35_140), .C2 (n_41_137) );
AOI211_X1 g_27_148 (.ZN (n_27_148), .A (n_24_147), .B (n_29_143), .C1 (n_33_141), .C2 (n_39_138) );
AOI211_X1 g_28_146 (.ZN (n_28_146), .A (n_26_146), .B (n_27_144), .C1 (n_31_142), .C2 (n_37_139) );
AOI211_X1 g_29_148 (.ZN (n_29_148), .A (n_27_148), .B (n_25_145), .C1 (n_29_143), .C2 (n_35_140) );
AOI211_X1 g_30_150 (.ZN (n_30_150), .A (n_28_146), .B (n_24_147), .C1 (n_27_144), .C2 (n_33_141) );
AOI211_X1 g_28_149 (.ZN (n_28_149), .A (n_29_148), .B (n_26_146), .C1 (n_25_145), .C2 (n_31_142) );
AOI211_X1 g_26_148 (.ZN (n_26_148), .A (n_30_150), .B (n_27_148), .C1 (n_24_147), .C2 (n_29_143) );
AOI211_X1 g_27_146 (.ZN (n_27_146), .A (n_28_149), .B (n_28_146), .C1 (n_26_146), .C2 (n_27_144) );
AOI211_X1 g_29_145 (.ZN (n_29_145), .A (n_26_148), .B (n_29_148), .C1 (n_27_148), .C2 (n_25_145) );
AOI211_X1 g_28_147 (.ZN (n_28_147), .A (n_27_146), .B (n_30_150), .C1 (n_28_146), .C2 (n_24_147) );
AOI211_X1 g_30_148 (.ZN (n_30_148), .A (n_29_145), .B (n_28_149), .C1 (n_29_148), .C2 (n_26_146) );
AOI211_X1 g_32_147 (.ZN (n_32_147), .A (n_28_147), .B (n_26_148), .C1 (n_30_150), .C2 (n_27_148) );
AOI211_X1 g_30_146 (.ZN (n_30_146), .A (n_30_148), .B (n_27_146), .C1 (n_28_149), .C2 (n_28_146) );
AOI211_X1 g_28_145 (.ZN (n_28_145), .A (n_32_147), .B (n_29_145), .C1 (n_26_148), .C2 (n_29_148) );
AOI211_X1 g_30_144 (.ZN (n_30_144), .A (n_30_146), .B (n_28_147), .C1 (n_27_146), .C2 (n_30_150) );
AOI211_X1 g_32_143 (.ZN (n_32_143), .A (n_28_145), .B (n_30_148), .C1 (n_29_145), .C2 (n_28_149) );
AOI211_X1 g_34_142 (.ZN (n_34_142), .A (n_30_144), .B (n_32_147), .C1 (n_28_147), .C2 (n_26_148) );
AOI211_X1 g_36_141 (.ZN (n_36_141), .A (n_32_143), .B (n_30_146), .C1 (n_30_148), .C2 (n_27_146) );
AOI211_X1 g_38_140 (.ZN (n_38_140), .A (n_34_142), .B (n_28_145), .C1 (n_32_147), .C2 (n_29_145) );
AOI211_X1 g_37_142 (.ZN (n_37_142), .A (n_36_141), .B (n_30_144), .C1 (n_30_146), .C2 (n_28_147) );
AOI211_X1 g_35_143 (.ZN (n_35_143), .A (n_38_140), .B (n_32_143), .C1 (n_28_145), .C2 (n_30_148) );
AOI211_X1 g_33_144 (.ZN (n_33_144), .A (n_37_142), .B (n_34_142), .C1 (n_30_144), .C2 (n_32_147) );
AOI211_X1 g_32_146 (.ZN (n_32_146), .A (n_35_143), .B (n_36_141), .C1 (n_32_143), .C2 (n_30_146) );
AOI211_X1 g_31_144 (.ZN (n_31_144), .A (n_33_144), .B (n_38_140), .C1 (n_34_142), .C2 (n_28_145) );
AOI211_X1 g_33_143 (.ZN (n_33_143), .A (n_32_146), .B (n_37_142), .C1 (n_36_141), .C2 (n_30_144) );
AOI211_X1 g_35_142 (.ZN (n_35_142), .A (n_31_144), .B (n_35_143), .C1 (n_38_140), .C2 (n_32_143) );
AOI211_X1 g_37_141 (.ZN (n_37_141), .A (n_33_143), .B (n_33_144), .C1 (n_37_142), .C2 (n_34_142) );
AOI211_X1 g_39_140 (.ZN (n_39_140), .A (n_35_142), .B (n_32_146), .C1 (n_35_143), .C2 (n_36_141) );
AOI211_X1 g_41_139 (.ZN (n_41_139), .A (n_37_141), .B (n_31_144), .C1 (n_33_144), .C2 (n_38_140) );
AOI211_X1 g_43_138 (.ZN (n_43_138), .A (n_39_140), .B (n_33_143), .C1 (n_32_146), .C2 (n_37_142) );
AOI211_X1 g_45_139 (.ZN (n_45_139), .A (n_41_139), .B (n_35_142), .C1 (n_31_144), .C2 (n_35_143) );
AOI211_X1 g_43_140 (.ZN (n_43_140), .A (n_43_138), .B (n_37_141), .C1 (n_33_143), .C2 (n_33_144) );
AOI211_X1 g_41_141 (.ZN (n_41_141), .A (n_45_139), .B (n_39_140), .C1 (n_35_142), .C2 (n_32_146) );
AOI211_X1 g_42_139 (.ZN (n_42_139), .A (n_43_140), .B (n_41_139), .C1 (n_37_141), .C2 (n_31_144) );
AOI211_X1 g_40_140 (.ZN (n_40_140), .A (n_41_141), .B (n_43_138), .C1 (n_39_140), .C2 (n_33_143) );
AOI211_X1 g_38_141 (.ZN (n_38_141), .A (n_42_139), .B (n_45_139), .C1 (n_41_139), .C2 (n_35_142) );
AOI211_X1 g_36_142 (.ZN (n_36_142), .A (n_40_140), .B (n_43_140), .C1 (n_43_138), .C2 (n_37_141) );
AOI211_X1 g_34_143 (.ZN (n_34_143), .A (n_38_141), .B (n_41_141), .C1 (n_45_139), .C2 (n_39_140) );
AOI211_X1 g_33_145 (.ZN (n_33_145), .A (n_36_142), .B (n_42_139), .C1 (n_43_140), .C2 (n_41_139) );
AOI211_X1 g_31_146 (.ZN (n_31_146), .A (n_34_143), .B (n_40_140), .C1 (n_41_141), .C2 (n_43_138) );
AOI211_X1 g_29_147 (.ZN (n_29_147), .A (n_33_145), .B (n_38_141), .C1 (n_42_139), .C2 (n_45_139) );
AOI211_X1 g_31_148 (.ZN (n_31_148), .A (n_31_146), .B (n_36_142), .C1 (n_40_140), .C2 (n_43_140) );
AOI211_X1 g_33_147 (.ZN (n_33_147), .A (n_29_147), .B (n_34_143), .C1 (n_38_141), .C2 (n_41_141) );
AOI211_X1 g_32_145 (.ZN (n_32_145), .A (n_31_148), .B (n_33_145), .C1 (n_36_142), .C2 (n_42_139) );
AOI211_X1 g_34_144 (.ZN (n_34_144), .A (n_33_147), .B (n_31_146), .C1 (n_34_143), .C2 (n_40_140) );
AOI211_X1 g_36_143 (.ZN (n_36_143), .A (n_32_145), .B (n_29_147), .C1 (n_33_145), .C2 (n_38_141) );
AOI211_X1 g_38_142 (.ZN (n_38_142), .A (n_34_144), .B (n_31_148), .C1 (n_31_146), .C2 (n_36_142) );
AOI211_X1 g_40_141 (.ZN (n_40_141), .A (n_36_143), .B (n_33_147), .C1 (n_29_147), .C2 (n_34_143) );
AOI211_X1 g_42_140 (.ZN (n_42_140), .A (n_38_142), .B (n_32_145), .C1 (n_31_148), .C2 (n_33_145) );
AOI211_X1 g_44_139 (.ZN (n_44_139), .A (n_40_141), .B (n_34_144), .C1 (n_33_147), .C2 (n_31_146) );
AOI211_X1 g_43_141 (.ZN (n_43_141), .A (n_42_140), .B (n_36_143), .C1 (n_32_145), .C2 (n_29_147) );
AOI211_X1 g_41_142 (.ZN (n_41_142), .A (n_44_139), .B (n_38_142), .C1 (n_34_144), .C2 (n_31_148) );
AOI211_X1 g_39_143 (.ZN (n_39_143), .A (n_43_141), .B (n_40_141), .C1 (n_36_143), .C2 (n_33_147) );
AOI211_X1 g_37_144 (.ZN (n_37_144), .A (n_41_142), .B (n_42_140), .C1 (n_38_142), .C2 (n_32_145) );
AOI211_X1 g_35_145 (.ZN (n_35_145), .A (n_39_143), .B (n_44_139), .C1 (n_40_141), .C2 (n_34_144) );
AOI211_X1 g_33_146 (.ZN (n_33_146), .A (n_37_144), .B (n_43_141), .C1 (n_42_140), .C2 (n_36_143) );
AOI211_X1 g_32_144 (.ZN (n_32_144), .A (n_35_145), .B (n_41_142), .C1 (n_44_139), .C2 (n_38_142) );
AOI211_X1 g_30_145 (.ZN (n_30_145), .A (n_33_146), .B (n_39_143), .C1 (n_43_141), .C2 (n_40_141) );
AOI211_X1 g_31_147 (.ZN (n_31_147), .A (n_32_144), .B (n_37_144), .C1 (n_41_142), .C2 (n_42_140) );
AOI211_X1 g_32_149 (.ZN (n_32_149), .A (n_30_145), .B (n_35_145), .C1 (n_39_143), .C2 (n_44_139) );
AOI211_X1 g_34_148 (.ZN (n_34_148), .A (n_31_147), .B (n_33_146), .C1 (n_37_144), .C2 (n_43_141) );
AOI211_X1 g_35_146 (.ZN (n_35_146), .A (n_32_149), .B (n_32_144), .C1 (n_35_145), .C2 (n_41_142) );
AOI211_X1 g_36_144 (.ZN (n_36_144), .A (n_34_148), .B (n_30_145), .C1 (n_33_146), .C2 (n_39_143) );
AOI211_X1 g_34_145 (.ZN (n_34_145), .A (n_35_146), .B (n_31_147), .C1 (n_32_144), .C2 (n_37_144) );
AOI211_X1 g_36_146 (.ZN (n_36_146), .A (n_36_144), .B (n_32_149), .C1 (n_30_145), .C2 (n_35_145) );
AOI211_X1 g_35_144 (.ZN (n_35_144), .A (n_34_145), .B (n_34_148), .C1 (n_31_147), .C2 (n_33_146) );
AOI211_X1 g_37_143 (.ZN (n_37_143), .A (n_36_146), .B (n_35_146), .C1 (n_32_149), .C2 (n_32_144) );
AOI211_X1 g_39_142 (.ZN (n_39_142), .A (n_35_144), .B (n_36_144), .C1 (n_34_148), .C2 (n_30_145) );
AOI211_X1 g_38_144 (.ZN (n_38_144), .A (n_37_143), .B (n_34_145), .C1 (n_35_146), .C2 (n_31_147) );
AOI211_X1 g_40_143 (.ZN (n_40_143), .A (n_39_142), .B (n_36_146), .C1 (n_36_144), .C2 (n_32_149) );
AOI211_X1 g_42_142 (.ZN (n_42_142), .A (n_38_144), .B (n_35_144), .C1 (n_34_145), .C2 (n_34_148) );
AOI211_X1 g_44_141 (.ZN (n_44_141), .A (n_40_143), .B (n_37_143), .C1 (n_36_146), .C2 (n_35_146) );
AOI211_X1 g_46_140 (.ZN (n_46_140), .A (n_42_142), .B (n_39_142), .C1 (n_35_144), .C2 (n_36_144) );
AOI211_X1 g_48_139 (.ZN (n_48_139), .A (n_44_141), .B (n_38_144), .C1 (n_37_143), .C2 (n_34_145) );
AOI211_X1 g_50_138 (.ZN (n_50_138), .A (n_46_140), .B (n_40_143), .C1 (n_39_142), .C2 (n_36_146) );
AOI211_X1 g_52_137 (.ZN (n_52_137), .A (n_48_139), .B (n_42_142), .C1 (n_38_144), .C2 (n_35_144) );
AOI211_X1 g_54_136 (.ZN (n_54_136), .A (n_50_138), .B (n_44_141), .C1 (n_40_143), .C2 (n_37_143) );
AOI211_X1 g_56_135 (.ZN (n_56_135), .A (n_52_137), .B (n_46_140), .C1 (n_42_142), .C2 (n_39_142) );
AOI211_X1 g_58_134 (.ZN (n_58_134), .A (n_54_136), .B (n_48_139), .C1 (n_44_141), .C2 (n_38_144) );
AOI211_X1 g_60_133 (.ZN (n_60_133), .A (n_56_135), .B (n_50_138), .C1 (n_46_140), .C2 (n_40_143) );
AOI211_X1 g_62_132 (.ZN (n_62_132), .A (n_58_134), .B (n_52_137), .C1 (n_48_139), .C2 (n_42_142) );
AOI211_X1 g_64_131 (.ZN (n_64_131), .A (n_60_133), .B (n_54_136), .C1 (n_50_138), .C2 (n_44_141) );
AOI211_X1 g_66_130 (.ZN (n_66_130), .A (n_62_132), .B (n_56_135), .C1 (n_52_137), .C2 (n_46_140) );
AOI211_X1 g_68_129 (.ZN (n_68_129), .A (n_64_131), .B (n_58_134), .C1 (n_54_136), .C2 (n_48_139) );
AOI211_X1 g_67_131 (.ZN (n_67_131), .A (n_66_130), .B (n_60_133), .C1 (n_56_135), .C2 (n_50_138) );
AOI211_X1 g_69_130 (.ZN (n_69_130), .A (n_68_129), .B (n_62_132), .C1 (n_58_134), .C2 (n_52_137) );
AOI211_X1 g_71_129 (.ZN (n_71_129), .A (n_67_131), .B (n_64_131), .C1 (n_60_133), .C2 (n_54_136) );
AOI211_X1 g_73_128 (.ZN (n_73_128), .A (n_69_130), .B (n_66_130), .C1 (n_62_132), .C2 (n_56_135) );
AOI211_X1 g_72_130 (.ZN (n_72_130), .A (n_71_129), .B (n_68_129), .C1 (n_64_131), .C2 (n_58_134) );
AOI211_X1 g_74_129 (.ZN (n_74_129), .A (n_73_128), .B (n_67_131), .C1 (n_66_130), .C2 (n_60_133) );
AOI211_X1 g_76_128 (.ZN (n_76_128), .A (n_72_130), .B (n_69_130), .C1 (n_68_129), .C2 (n_62_132) );
AOI211_X1 g_78_127 (.ZN (n_78_127), .A (n_74_129), .B (n_71_129), .C1 (n_67_131), .C2 (n_64_131) );
AOI211_X1 g_80_126 (.ZN (n_80_126), .A (n_76_128), .B (n_73_128), .C1 (n_69_130), .C2 (n_66_130) );
AOI211_X1 g_79_128 (.ZN (n_79_128), .A (n_78_127), .B (n_72_130), .C1 (n_71_129), .C2 (n_68_129) );
AOI211_X1 g_78_126 (.ZN (n_78_126), .A (n_80_126), .B (n_74_129), .C1 (n_73_128), .C2 (n_67_131) );
AOI211_X1 g_80_125 (.ZN (n_80_125), .A (n_79_128), .B (n_76_128), .C1 (n_72_130), .C2 (n_69_130) );
AOI211_X1 g_82_124 (.ZN (n_82_124), .A (n_78_126), .B (n_78_127), .C1 (n_74_129), .C2 (n_71_129) );
AOI211_X1 g_84_123 (.ZN (n_84_123), .A (n_80_125), .B (n_80_126), .C1 (n_76_128), .C2 (n_73_128) );
AOI211_X1 g_86_122 (.ZN (n_86_122), .A (n_82_124), .B (n_79_128), .C1 (n_78_127), .C2 (n_72_130) );
AOI211_X1 g_88_121 (.ZN (n_88_121), .A (n_84_123), .B (n_78_126), .C1 (n_80_126), .C2 (n_74_129) );
AOI211_X1 g_90_120 (.ZN (n_90_120), .A (n_86_122), .B (n_80_125), .C1 (n_79_128), .C2 (n_76_128) );
AOI211_X1 g_92_119 (.ZN (n_92_119), .A (n_88_121), .B (n_82_124), .C1 (n_78_126), .C2 (n_78_127) );
AOI211_X1 g_94_118 (.ZN (n_94_118), .A (n_90_120), .B (n_84_123), .C1 (n_80_125), .C2 (n_80_126) );
AOI211_X1 g_95_116 (.ZN (n_95_116), .A (n_92_119), .B (n_86_122), .C1 (n_82_124), .C2 (n_79_128) );
AOI211_X1 g_97_115 (.ZN (n_97_115), .A (n_94_118), .B (n_88_121), .C1 (n_84_123), .C2 (n_78_126) );
AOI211_X1 g_96_117 (.ZN (n_96_117), .A (n_95_116), .B (n_90_120), .C1 (n_86_122), .C2 (n_80_125) );
AOI211_X1 g_98_116 (.ZN (n_98_116), .A (n_97_115), .B (n_92_119), .C1 (n_88_121), .C2 (n_82_124) );
AOI211_X1 g_100_115 (.ZN (n_100_115), .A (n_96_117), .B (n_94_118), .C1 (n_90_120), .C2 (n_84_123) );
AOI211_X1 g_101_113 (.ZN (n_101_113), .A (n_98_116), .B (n_95_116), .C1 (n_92_119), .C2 (n_86_122) );
AOI211_X1 g_103_112 (.ZN (n_103_112), .A (n_100_115), .B (n_97_115), .C1 (n_94_118), .C2 (n_88_121) );
AOI211_X1 g_105_111 (.ZN (n_105_111), .A (n_101_113), .B (n_96_117), .C1 (n_95_116), .C2 (n_90_120) );
AOI211_X1 g_107_110 (.ZN (n_107_110), .A (n_103_112), .B (n_98_116), .C1 (n_97_115), .C2 (n_92_119) );
AOI211_X1 g_109_109 (.ZN (n_109_109), .A (n_105_111), .B (n_100_115), .C1 (n_96_117), .C2 (n_94_118) );
AOI211_X1 g_111_108 (.ZN (n_111_108), .A (n_107_110), .B (n_101_113), .C1 (n_98_116), .C2 (n_95_116) );
AOI211_X1 g_113_107 (.ZN (n_113_107), .A (n_109_109), .B (n_103_112), .C1 (n_100_115), .C2 (n_97_115) );
AOI211_X1 g_115_106 (.ZN (n_115_106), .A (n_111_108), .B (n_105_111), .C1 (n_101_113), .C2 (n_96_117) );
AOI211_X1 g_117_105 (.ZN (n_117_105), .A (n_113_107), .B (n_107_110), .C1 (n_103_112), .C2 (n_98_116) );
AOI211_X1 g_119_104 (.ZN (n_119_104), .A (n_115_106), .B (n_109_109), .C1 (n_105_111), .C2 (n_100_115) );
AOI211_X1 g_121_103 (.ZN (n_121_103), .A (n_117_105), .B (n_111_108), .C1 (n_107_110), .C2 (n_101_113) );
AOI211_X1 g_120_105 (.ZN (n_120_105), .A (n_119_104), .B (n_113_107), .C1 (n_109_109), .C2 (n_103_112) );
AOI211_X1 g_122_104 (.ZN (n_122_104), .A (n_121_103), .B (n_115_106), .C1 (n_111_108), .C2 (n_105_111) );
AOI211_X1 g_124_103 (.ZN (n_124_103), .A (n_120_105), .B (n_117_105), .C1 (n_113_107), .C2 (n_107_110) );
AOI211_X1 g_126_102 (.ZN (n_126_102), .A (n_122_104), .B (n_119_104), .C1 (n_115_106), .C2 (n_109_109) );
AOI211_X1 g_128_101 (.ZN (n_128_101), .A (n_124_103), .B (n_121_103), .C1 (n_117_105), .C2 (n_111_108) );
AOI211_X1 g_130_100 (.ZN (n_130_100), .A (n_126_102), .B (n_120_105), .C1 (n_119_104), .C2 (n_113_107) );
AOI211_X1 g_132_99 (.ZN (n_132_99), .A (n_128_101), .B (n_122_104), .C1 (n_121_103), .C2 (n_115_106) );
AOI211_X1 g_134_98 (.ZN (n_134_98), .A (n_130_100), .B (n_124_103), .C1 (n_120_105), .C2 (n_117_105) );
AOI211_X1 g_136_97 (.ZN (n_136_97), .A (n_132_99), .B (n_126_102), .C1 (n_122_104), .C2 (n_119_104) );
AOI211_X1 g_138_98 (.ZN (n_138_98), .A (n_134_98), .B (n_128_101), .C1 (n_124_103), .C2 (n_121_103) );
AOI211_X1 g_139_96 (.ZN (n_139_96), .A (n_136_97), .B (n_130_100), .C1 (n_126_102), .C2 (n_120_105) );
AOI211_X1 g_141_95 (.ZN (n_141_95), .A (n_138_98), .B (n_132_99), .C1 (n_128_101), .C2 (n_122_104) );
AOI211_X1 g_142_93 (.ZN (n_142_93), .A (n_139_96), .B (n_134_98), .C1 (n_130_100), .C2 (n_124_103) );
AOI211_X1 g_140_94 (.ZN (n_140_94), .A (n_141_95), .B (n_136_97), .C1 (n_132_99), .C2 (n_126_102) );
AOI211_X1 g_138_95 (.ZN (n_138_95), .A (n_142_93), .B (n_138_98), .C1 (n_134_98), .C2 (n_128_101) );
AOI211_X1 g_136_96 (.ZN (n_136_96), .A (n_140_94), .B (n_139_96), .C1 (n_136_97), .C2 (n_130_100) );
AOI211_X1 g_134_97 (.ZN (n_134_97), .A (n_138_95), .B (n_141_95), .C1 (n_138_98), .C2 (n_132_99) );
AOI211_X1 g_132_98 (.ZN (n_132_98), .A (n_136_96), .B (n_142_93), .C1 (n_139_96), .C2 (n_134_98) );
AOI211_X1 g_130_99 (.ZN (n_130_99), .A (n_134_97), .B (n_140_94), .C1 (n_141_95), .C2 (n_136_97) );
AOI211_X1 g_128_100 (.ZN (n_128_100), .A (n_132_98), .B (n_138_95), .C1 (n_142_93), .C2 (n_138_98) );
AOI211_X1 g_126_101 (.ZN (n_126_101), .A (n_130_99), .B (n_136_96), .C1 (n_140_94), .C2 (n_139_96) );
AOI211_X1 g_124_102 (.ZN (n_124_102), .A (n_128_100), .B (n_134_97), .C1 (n_138_95), .C2 (n_141_95) );
AOI211_X1 g_123_104 (.ZN (n_123_104), .A (n_126_101), .B (n_132_98), .C1 (n_136_96), .C2 (n_142_93) );
AOI211_X1 g_125_103 (.ZN (n_125_103), .A (n_124_102), .B (n_130_99), .C1 (n_134_97), .C2 (n_140_94) );
AOI211_X1 g_127_102 (.ZN (n_127_102), .A (n_123_104), .B (n_128_100), .C1 (n_132_98), .C2 (n_138_95) );
AOI211_X1 g_129_101 (.ZN (n_129_101), .A (n_125_103), .B (n_126_101), .C1 (n_130_99), .C2 (n_136_96) );
AOI211_X1 g_131_100 (.ZN (n_131_100), .A (n_127_102), .B (n_124_102), .C1 (n_128_100), .C2 (n_134_97) );
AOI211_X1 g_133_99 (.ZN (n_133_99), .A (n_129_101), .B (n_123_104), .C1 (n_126_101), .C2 (n_132_98) );
AOI211_X1 g_135_98 (.ZN (n_135_98), .A (n_131_100), .B (n_125_103), .C1 (n_124_102), .C2 (n_130_99) );
AOI211_X1 g_137_97 (.ZN (n_137_97), .A (n_133_99), .B (n_127_102), .C1 (n_123_104), .C2 (n_128_100) );
AOI211_X1 g_136_99 (.ZN (n_136_99), .A (n_135_98), .B (n_129_101), .C1 (n_125_103), .C2 (n_126_101) );
AOI211_X1 g_134_100 (.ZN (n_134_100), .A (n_137_97), .B (n_131_100), .C1 (n_127_102), .C2 (n_124_102) );
AOI211_X1 g_132_101 (.ZN (n_132_101), .A (n_136_99), .B (n_133_99), .C1 (n_129_101), .C2 (n_123_104) );
AOI211_X1 g_130_102 (.ZN (n_130_102), .A (n_134_100), .B (n_135_98), .C1 (n_131_100), .C2 (n_125_103) );
AOI211_X1 g_128_103 (.ZN (n_128_103), .A (n_132_101), .B (n_137_97), .C1 (n_133_99), .C2 (n_127_102) );
AOI211_X1 g_126_104 (.ZN (n_126_104), .A (n_130_102), .B (n_136_99), .C1 (n_135_98), .C2 (n_129_101) );
AOI211_X1 g_124_105 (.ZN (n_124_105), .A (n_128_103), .B (n_134_100), .C1 (n_137_97), .C2 (n_131_100) );
AOI211_X1 g_122_106 (.ZN (n_122_106), .A (n_126_104), .B (n_132_101), .C1 (n_136_99), .C2 (n_133_99) );
AOI211_X1 g_120_107 (.ZN (n_120_107), .A (n_124_105), .B (n_130_102), .C1 (n_134_100), .C2 (n_135_98) );
AOI211_X1 g_121_105 (.ZN (n_121_105), .A (n_122_106), .B (n_128_103), .C1 (n_132_101), .C2 (n_137_97) );
AOI211_X1 g_119_106 (.ZN (n_119_106), .A (n_120_107), .B (n_126_104), .C1 (n_130_102), .C2 (n_136_99) );
AOI211_X1 g_117_107 (.ZN (n_117_107), .A (n_121_105), .B (n_124_105), .C1 (n_128_103), .C2 (n_134_100) );
AOI211_X1 g_115_108 (.ZN (n_115_108), .A (n_119_106), .B (n_122_106), .C1 (n_126_104), .C2 (n_132_101) );
AOI211_X1 g_113_109 (.ZN (n_113_109), .A (n_117_107), .B (n_120_107), .C1 (n_124_105), .C2 (n_130_102) );
AOI211_X1 g_111_110 (.ZN (n_111_110), .A (n_115_108), .B (n_121_105), .C1 (n_122_106), .C2 (n_128_103) );
AOI211_X1 g_109_111 (.ZN (n_109_111), .A (n_113_109), .B (n_119_106), .C1 (n_120_107), .C2 (n_126_104) );
AOI211_X1 g_107_112 (.ZN (n_107_112), .A (n_111_110), .B (n_117_107), .C1 (n_121_105), .C2 (n_124_105) );
AOI211_X1 g_105_113 (.ZN (n_105_113), .A (n_109_111), .B (n_115_108), .C1 (n_119_106), .C2 (n_122_106) );
AOI211_X1 g_103_114 (.ZN (n_103_114), .A (n_107_112), .B (n_113_109), .C1 (n_117_107), .C2 (n_120_107) );
AOI211_X1 g_101_115 (.ZN (n_101_115), .A (n_105_113), .B (n_111_110), .C1 (n_115_108), .C2 (n_121_105) );
AOI211_X1 g_99_116 (.ZN (n_99_116), .A (n_103_114), .B (n_109_111), .C1 (n_113_109), .C2 (n_119_106) );
AOI211_X1 g_97_117 (.ZN (n_97_117), .A (n_101_115), .B (n_107_112), .C1 (n_111_110), .C2 (n_117_107) );
AOI211_X1 g_95_118 (.ZN (n_95_118), .A (n_99_116), .B (n_105_113), .C1 (n_109_111), .C2 (n_115_108) );
AOI211_X1 g_93_119 (.ZN (n_93_119), .A (n_97_117), .B (n_103_114), .C1 (n_107_112), .C2 (n_113_109) );
AOI211_X1 g_91_120 (.ZN (n_91_120), .A (n_95_118), .B (n_101_115), .C1 (n_105_113), .C2 (n_111_110) );
AOI211_X1 g_90_122 (.ZN (n_90_122), .A (n_93_119), .B (n_99_116), .C1 (n_103_114), .C2 (n_109_111) );
AOI211_X1 g_92_121 (.ZN (n_92_121), .A (n_91_120), .B (n_97_117), .C1 (n_101_115), .C2 (n_107_112) );
AOI211_X1 g_94_120 (.ZN (n_94_120), .A (n_90_122), .B (n_95_118), .C1 (n_99_116), .C2 (n_105_113) );
AOI211_X1 g_96_119 (.ZN (n_96_119), .A (n_92_121), .B (n_93_119), .C1 (n_97_117), .C2 (n_103_114) );
AOI211_X1 g_98_118 (.ZN (n_98_118), .A (n_94_120), .B (n_91_120), .C1 (n_95_118), .C2 (n_101_115) );
AOI211_X1 g_100_117 (.ZN (n_100_117), .A (n_96_119), .B (n_90_122), .C1 (n_93_119), .C2 (n_99_116) );
AOI211_X1 g_102_116 (.ZN (n_102_116), .A (n_98_118), .B (n_92_121), .C1 (n_91_120), .C2 (n_97_117) );
AOI211_X1 g_104_115 (.ZN (n_104_115), .A (n_100_117), .B (n_94_120), .C1 (n_90_122), .C2 (n_95_118) );
AOI211_X1 g_102_114 (.ZN (n_102_114), .A (n_102_116), .B (n_96_119), .C1 (n_92_121), .C2 (n_93_119) );
AOI211_X1 g_104_113 (.ZN (n_104_113), .A (n_104_115), .B (n_98_118), .C1 (n_94_120), .C2 (n_91_120) );
AOI211_X1 g_106_112 (.ZN (n_106_112), .A (n_102_114), .B (n_100_117), .C1 (n_96_119), .C2 (n_90_122) );
AOI211_X1 g_108_111 (.ZN (n_108_111), .A (n_104_113), .B (n_102_116), .C1 (n_98_118), .C2 (n_92_121) );
AOI211_X1 g_110_110 (.ZN (n_110_110), .A (n_106_112), .B (n_104_115), .C1 (n_100_117), .C2 (n_94_120) );
AOI211_X1 g_112_109 (.ZN (n_112_109), .A (n_108_111), .B (n_102_114), .C1 (n_102_116), .C2 (n_96_119) );
AOI211_X1 g_114_108 (.ZN (n_114_108), .A (n_110_110), .B (n_104_113), .C1 (n_104_115), .C2 (n_98_118) );
AOI211_X1 g_116_107 (.ZN (n_116_107), .A (n_112_109), .B (n_106_112), .C1 (n_102_114), .C2 (n_100_117) );
AOI211_X1 g_118_106 (.ZN (n_118_106), .A (n_114_108), .B (n_108_111), .C1 (n_104_113), .C2 (n_102_116) );
AOI211_X1 g_117_108 (.ZN (n_117_108), .A (n_116_107), .B (n_110_110), .C1 (n_106_112), .C2 (n_104_115) );
AOI211_X1 g_119_107 (.ZN (n_119_107), .A (n_118_106), .B (n_112_109), .C1 (n_108_111), .C2 (n_102_114) );
AOI211_X1 g_121_106 (.ZN (n_121_106), .A (n_117_108), .B (n_114_108), .C1 (n_110_110), .C2 (n_104_113) );
AOI211_X1 g_123_105 (.ZN (n_123_105), .A (n_119_107), .B (n_116_107), .C1 (n_112_109), .C2 (n_106_112) );
AOI211_X1 g_125_104 (.ZN (n_125_104), .A (n_121_106), .B (n_118_106), .C1 (n_114_108), .C2 (n_108_111) );
AOI211_X1 g_127_103 (.ZN (n_127_103), .A (n_123_105), .B (n_117_108), .C1 (n_116_107), .C2 (n_110_110) );
AOI211_X1 g_129_102 (.ZN (n_129_102), .A (n_125_104), .B (n_119_107), .C1 (n_118_106), .C2 (n_112_109) );
AOI211_X1 g_131_101 (.ZN (n_131_101), .A (n_127_103), .B (n_121_106), .C1 (n_117_108), .C2 (n_114_108) );
AOI211_X1 g_133_100 (.ZN (n_133_100), .A (n_129_102), .B (n_123_105), .C1 (n_119_107), .C2 (n_116_107) );
AOI211_X1 g_135_99 (.ZN (n_135_99), .A (n_131_101), .B (n_125_104), .C1 (n_121_106), .C2 (n_118_106) );
AOI211_X1 g_137_98 (.ZN (n_137_98), .A (n_133_100), .B (n_127_103), .C1 (n_123_105), .C2 (n_117_108) );
AOI211_X1 g_139_97 (.ZN (n_139_97), .A (n_135_99), .B (n_129_102), .C1 (n_125_104), .C2 (n_119_107) );
AOI211_X1 g_141_96 (.ZN (n_141_96), .A (n_137_98), .B (n_131_101), .C1 (n_127_103), .C2 (n_121_106) );
AOI211_X1 g_143_95 (.ZN (n_143_95), .A (n_139_97), .B (n_133_100), .C1 (n_129_102), .C2 (n_123_105) );
AOI211_X1 g_144_97 (.ZN (n_144_97), .A (n_141_96), .B (n_135_99), .C1 (n_131_101), .C2 (n_125_104) );
AOI211_X1 g_146_98 (.ZN (n_146_98), .A (n_143_95), .B (n_137_98), .C1 (n_133_100), .C2 (n_127_103) );
AOI211_X1 g_148_99 (.ZN (n_148_99), .A (n_144_97), .B (n_139_97), .C1 (n_135_99), .C2 (n_129_102) );
AOI211_X1 g_147_97 (.ZN (n_147_97), .A (n_146_98), .B (n_141_96), .C1 (n_137_98), .C2 (n_131_101) );
AOI211_X1 g_146_95 (.ZN (n_146_95), .A (n_148_99), .B (n_143_95), .C1 (n_139_97), .C2 (n_133_100) );
AOI211_X1 g_144_94 (.ZN (n_144_94), .A (n_147_97), .B (n_144_97), .C1 (n_141_96), .C2 (n_135_99) );
AOI211_X1 g_145_96 (.ZN (n_145_96), .A (n_146_95), .B (n_146_98), .C1 (n_143_95), .C2 (n_137_98) );
AOI211_X1 g_143_97 (.ZN (n_143_97), .A (n_144_94), .B (n_148_99), .C1 (n_144_97), .C2 (n_139_97) );
AOI211_X1 g_142_95 (.ZN (n_142_95), .A (n_145_96), .B (n_147_97), .C1 (n_146_98), .C2 (n_141_96) );
AOI211_X1 g_144_96 (.ZN (n_144_96), .A (n_143_97), .B (n_146_95), .C1 (n_148_99), .C2 (n_143_95) );
AOI211_X1 g_145_98 (.ZN (n_145_98), .A (n_142_95), .B (n_144_94), .C1 (n_147_97), .C2 (n_144_97) );
AOI211_X1 g_146_100 (.ZN (n_146_100), .A (n_144_96), .B (n_145_96), .C1 (n_146_95), .C2 (n_146_98) );
AOI211_X1 g_144_99 (.ZN (n_144_99), .A (n_145_98), .B (n_143_97), .C1 (n_144_94), .C2 (n_148_99) );
AOI211_X1 g_145_97 (.ZN (n_145_97), .A (n_146_100), .B (n_142_95), .C1 (n_145_96), .C2 (n_147_97) );
AOI211_X1 g_143_96 (.ZN (n_143_96), .A (n_144_99), .B (n_144_96), .C1 (n_143_97), .C2 (n_146_95) );
AOI211_X1 g_142_98 (.ZN (n_142_98), .A (n_145_97), .B (n_145_98), .C1 (n_142_95), .C2 (n_144_94) );
AOI211_X1 g_140_99 (.ZN (n_140_99), .A (n_143_96), .B (n_146_100), .C1 (n_144_96), .C2 (n_145_96) );
AOI211_X1 g_141_97 (.ZN (n_141_97), .A (n_142_98), .B (n_144_99), .C1 (n_145_98), .C2 (n_143_97) );
AOI211_X1 g_143_98 (.ZN (n_143_98), .A (n_140_99), .B (n_145_97), .C1 (n_146_100), .C2 (n_142_95) );
AOI211_X1 g_142_100 (.ZN (n_142_100), .A (n_141_97), .B (n_143_96), .C1 (n_144_99), .C2 (n_144_96) );
AOI211_X1 g_141_98 (.ZN (n_141_98), .A (n_143_98), .B (n_142_98), .C1 (n_145_97), .C2 (n_145_98) );
AOI211_X1 g_140_96 (.ZN (n_140_96), .A (n_142_100), .B (n_140_99), .C1 (n_143_96), .C2 (n_146_100) );
AOI211_X1 g_138_97 (.ZN (n_138_97), .A (n_141_98), .B (n_141_97), .C1 (n_142_98), .C2 (n_144_99) );
AOI211_X1 g_136_98 (.ZN (n_136_98), .A (n_140_96), .B (n_143_98), .C1 (n_140_99), .C2 (n_145_97) );
AOI211_X1 g_134_99 (.ZN (n_134_99), .A (n_138_97), .B (n_142_100), .C1 (n_141_97), .C2 (n_143_96) );
AOI211_X1 g_133_101 (.ZN (n_133_101), .A (n_136_98), .B (n_141_98), .C1 (n_143_98), .C2 (n_142_98) );
AOI211_X1 g_135_100 (.ZN (n_135_100), .A (n_134_99), .B (n_140_96), .C1 (n_142_100), .C2 (n_140_99) );
AOI211_X1 g_137_99 (.ZN (n_137_99), .A (n_133_101), .B (n_138_97), .C1 (n_141_98), .C2 (n_141_97) );
AOI211_X1 g_139_98 (.ZN (n_139_98), .A (n_135_100), .B (n_136_98), .C1 (n_140_96), .C2 (n_143_98) );
AOI211_X1 g_138_100 (.ZN (n_138_100), .A (n_137_99), .B (n_134_99), .C1 (n_138_97), .C2 (n_142_100) );
AOI211_X1 g_136_101 (.ZN (n_136_101), .A (n_139_98), .B (n_133_101), .C1 (n_136_98), .C2 (n_141_98) );
AOI211_X1 g_134_102 (.ZN (n_134_102), .A (n_138_100), .B (n_135_100), .C1 (n_134_99), .C2 (n_140_96) );
AOI211_X1 g_132_103 (.ZN (n_132_103), .A (n_136_101), .B (n_137_99), .C1 (n_133_101), .C2 (n_138_97) );
AOI211_X1 g_130_104 (.ZN (n_130_104), .A (n_134_102), .B (n_139_98), .C1 (n_135_100), .C2 (n_136_98) );
AOI211_X1 g_131_102 (.ZN (n_131_102), .A (n_132_103), .B (n_138_100), .C1 (n_137_99), .C2 (n_134_99) );
AOI211_X1 g_129_103 (.ZN (n_129_103), .A (n_130_104), .B (n_136_101), .C1 (n_139_98), .C2 (n_133_101) );
AOI211_X1 g_130_101 (.ZN (n_130_101), .A (n_131_102), .B (n_134_102), .C1 (n_138_100), .C2 (n_135_100) );
AOI211_X1 g_128_102 (.ZN (n_128_102), .A (n_129_103), .B (n_132_103), .C1 (n_136_101), .C2 (n_137_99) );
AOI211_X1 g_126_103 (.ZN (n_126_103), .A (n_130_101), .B (n_130_104), .C1 (n_134_102), .C2 (n_139_98) );
AOI211_X1 g_124_104 (.ZN (n_124_104), .A (n_128_102), .B (n_131_102), .C1 (n_132_103), .C2 (n_138_100) );
AOI211_X1 g_122_105 (.ZN (n_122_105), .A (n_126_103), .B (n_129_103), .C1 (n_130_104), .C2 (n_136_101) );
AOI211_X1 g_120_106 (.ZN (n_120_106), .A (n_124_104), .B (n_130_101), .C1 (n_131_102), .C2 (n_134_102) );
AOI211_X1 g_118_107 (.ZN (n_118_107), .A (n_122_105), .B (n_128_102), .C1 (n_129_103), .C2 (n_132_103) );
AOI211_X1 g_116_108 (.ZN (n_116_108), .A (n_120_106), .B (n_126_103), .C1 (n_130_101), .C2 (n_130_104) );
AOI211_X1 g_114_109 (.ZN (n_114_109), .A (n_118_107), .B (n_124_104), .C1 (n_128_102), .C2 (n_131_102) );
AOI211_X1 g_112_110 (.ZN (n_112_110), .A (n_116_108), .B (n_122_105), .C1 (n_126_103), .C2 (n_129_103) );
AOI211_X1 g_110_111 (.ZN (n_110_111), .A (n_114_109), .B (n_120_106), .C1 (n_124_104), .C2 (n_130_101) );
AOI211_X1 g_108_112 (.ZN (n_108_112), .A (n_112_110), .B (n_118_107), .C1 (n_122_105), .C2 (n_128_102) );
AOI211_X1 g_106_113 (.ZN (n_106_113), .A (n_110_111), .B (n_116_108), .C1 (n_120_106), .C2 (n_126_103) );
AOI211_X1 g_104_114 (.ZN (n_104_114), .A (n_108_112), .B (n_114_109), .C1 (n_118_107), .C2 (n_124_104) );
AOI211_X1 g_102_115 (.ZN (n_102_115), .A (n_106_113), .B (n_112_110), .C1 (n_116_108), .C2 (n_122_105) );
AOI211_X1 g_100_116 (.ZN (n_100_116), .A (n_104_114), .B (n_110_111), .C1 (n_114_109), .C2 (n_120_106) );
AOI211_X1 g_98_117 (.ZN (n_98_117), .A (n_102_115), .B (n_108_112), .C1 (n_112_110), .C2 (n_118_107) );
AOI211_X1 g_96_118 (.ZN (n_96_118), .A (n_100_116), .B (n_106_113), .C1 (n_110_111), .C2 (n_116_108) );
AOI211_X1 g_94_119 (.ZN (n_94_119), .A (n_98_117), .B (n_104_114), .C1 (n_108_112), .C2 (n_114_109) );
AOI211_X1 g_92_120 (.ZN (n_92_120), .A (n_96_118), .B (n_102_115), .C1 (n_106_113), .C2 (n_112_110) );
AOI211_X1 g_90_121 (.ZN (n_90_121), .A (n_94_119), .B (n_100_116), .C1 (n_104_114), .C2 (n_110_111) );
AOI211_X1 g_88_122 (.ZN (n_88_122), .A (n_92_120), .B (n_98_117), .C1 (n_102_115), .C2 (n_108_112) );
AOI211_X1 g_86_123 (.ZN (n_86_123), .A (n_90_121), .B (n_96_118), .C1 (n_100_116), .C2 (n_106_113) );
AOI211_X1 g_84_124 (.ZN (n_84_124), .A (n_88_122), .B (n_94_119), .C1 (n_98_117), .C2 (n_104_114) );
AOI211_X1 g_83_126 (.ZN (n_83_126), .A (n_86_123), .B (n_92_120), .C1 (n_96_118), .C2 (n_102_115) );
AOI211_X1 g_81_125 (.ZN (n_81_125), .A (n_84_124), .B (n_90_121), .C1 (n_94_119), .C2 (n_100_116) );
AOI211_X1 g_83_124 (.ZN (n_83_124), .A (n_83_126), .B (n_88_122), .C1 (n_92_120), .C2 (n_98_117) );
AOI211_X1 g_85_123 (.ZN (n_85_123), .A (n_81_125), .B (n_86_123), .C1 (n_90_121), .C2 (n_96_118) );
AOI211_X1 g_87_122 (.ZN (n_87_122), .A (n_83_124), .B (n_84_124), .C1 (n_88_122), .C2 (n_94_119) );
AOI211_X1 g_86_124 (.ZN (n_86_124), .A (n_85_123), .B (n_83_126), .C1 (n_86_123), .C2 (n_92_120) );
AOI211_X1 g_88_123 (.ZN (n_88_123), .A (n_87_122), .B (n_81_125), .C1 (n_84_124), .C2 (n_90_121) );
AOI211_X1 g_87_125 (.ZN (n_87_125), .A (n_86_124), .B (n_83_124), .C1 (n_83_126), .C2 (n_88_122) );
AOI211_X1 g_85_124 (.ZN (n_85_124), .A (n_88_123), .B (n_85_123), .C1 (n_81_125), .C2 (n_86_123) );
AOI211_X1 g_87_123 (.ZN (n_87_123), .A (n_87_125), .B (n_87_122), .C1 (n_83_124), .C2 (n_84_124) );
AOI211_X1 g_89_122 (.ZN (n_89_122), .A (n_85_124), .B (n_86_124), .C1 (n_85_123), .C2 (n_83_126) );
AOI211_X1 g_91_121 (.ZN (n_91_121), .A (n_87_123), .B (n_88_123), .C1 (n_87_122), .C2 (n_81_125) );
AOI211_X1 g_93_120 (.ZN (n_93_120), .A (n_89_122), .B (n_87_125), .C1 (n_86_124), .C2 (n_83_124) );
AOI211_X1 g_95_119 (.ZN (n_95_119), .A (n_91_121), .B (n_85_124), .C1 (n_88_123), .C2 (n_85_123) );
AOI211_X1 g_97_118 (.ZN (n_97_118), .A (n_93_120), .B (n_87_123), .C1 (n_87_125), .C2 (n_87_122) );
AOI211_X1 g_99_117 (.ZN (n_99_117), .A (n_95_119), .B (n_89_122), .C1 (n_85_124), .C2 (n_86_124) );
AOI211_X1 g_101_116 (.ZN (n_101_116), .A (n_97_118), .B (n_91_121), .C1 (n_87_123), .C2 (n_88_123) );
AOI211_X1 g_103_115 (.ZN (n_103_115), .A (n_99_117), .B (n_93_120), .C1 (n_89_122), .C2 (n_87_125) );
AOI211_X1 g_105_114 (.ZN (n_105_114), .A (n_101_116), .B (n_95_119), .C1 (n_91_121), .C2 (n_85_124) );
AOI211_X1 g_107_113 (.ZN (n_107_113), .A (n_103_115), .B (n_97_118), .C1 (n_93_120), .C2 (n_87_123) );
AOI211_X1 g_109_112 (.ZN (n_109_112), .A (n_105_114), .B (n_99_117), .C1 (n_95_119), .C2 (n_89_122) );
AOI211_X1 g_111_111 (.ZN (n_111_111), .A (n_107_113), .B (n_101_116), .C1 (n_97_118), .C2 (n_91_121) );
AOI211_X1 g_113_110 (.ZN (n_113_110), .A (n_109_112), .B (n_103_115), .C1 (n_99_117), .C2 (n_93_120) );
AOI211_X1 g_115_109 (.ZN (n_115_109), .A (n_111_111), .B (n_105_114), .C1 (n_101_116), .C2 (n_95_119) );
AOI211_X1 g_114_111 (.ZN (n_114_111), .A (n_113_110), .B (n_107_113), .C1 (n_103_115), .C2 (n_97_118) );
AOI211_X1 g_116_110 (.ZN (n_116_110), .A (n_115_109), .B (n_109_112), .C1 (n_105_114), .C2 (n_99_117) );
AOI211_X1 g_118_109 (.ZN (n_118_109), .A (n_114_111), .B (n_111_111), .C1 (n_107_113), .C2 (n_101_116) );
AOI211_X1 g_120_108 (.ZN (n_120_108), .A (n_116_110), .B (n_113_110), .C1 (n_109_112), .C2 (n_103_115) );
AOI211_X1 g_122_107 (.ZN (n_122_107), .A (n_118_109), .B (n_115_109), .C1 (n_111_111), .C2 (n_105_114) );
AOI211_X1 g_124_106 (.ZN (n_124_106), .A (n_120_108), .B (n_114_111), .C1 (n_113_110), .C2 (n_107_113) );
AOI211_X1 g_126_105 (.ZN (n_126_105), .A (n_122_107), .B (n_116_110), .C1 (n_115_109), .C2 (n_109_112) );
AOI211_X1 g_128_104 (.ZN (n_128_104), .A (n_124_106), .B (n_118_109), .C1 (n_114_111), .C2 (n_111_111) );
AOI211_X1 g_130_103 (.ZN (n_130_103), .A (n_126_105), .B (n_120_108), .C1 (n_116_110), .C2 (n_113_110) );
AOI211_X1 g_132_102 (.ZN (n_132_102), .A (n_128_104), .B (n_122_107), .C1 (n_118_109), .C2 (n_115_109) );
AOI211_X1 g_134_101 (.ZN (n_134_101), .A (n_130_103), .B (n_124_106), .C1 (n_120_108), .C2 (n_114_111) );
AOI211_X1 g_136_100 (.ZN (n_136_100), .A (n_132_102), .B (n_126_105), .C1 (n_122_107), .C2 (n_116_110) );
AOI211_X1 g_138_99 (.ZN (n_138_99), .A (n_134_101), .B (n_128_104), .C1 (n_124_106), .C2 (n_118_109) );
AOI211_X1 g_140_98 (.ZN (n_140_98), .A (n_136_100), .B (n_130_103), .C1 (n_126_105), .C2 (n_120_108) );
AOI211_X1 g_142_97 (.ZN (n_142_97), .A (n_138_99), .B (n_132_102), .C1 (n_128_104), .C2 (n_122_107) );
AOI211_X1 g_141_99 (.ZN (n_141_99), .A (n_140_98), .B (n_134_101), .C1 (n_130_103), .C2 (n_124_106) );
AOI211_X1 g_139_100 (.ZN (n_139_100), .A (n_142_97), .B (n_136_100), .C1 (n_132_102), .C2 (n_126_105) );
AOI211_X1 g_137_101 (.ZN (n_137_101), .A (n_141_99), .B (n_138_99), .C1 (n_134_101), .C2 (n_128_104) );
AOI211_X1 g_135_102 (.ZN (n_135_102), .A (n_139_100), .B (n_140_98), .C1 (n_136_100), .C2 (n_130_103) );
AOI211_X1 g_133_103 (.ZN (n_133_103), .A (n_137_101), .B (n_142_97), .C1 (n_138_99), .C2 (n_132_102) );
AOI211_X1 g_131_104 (.ZN (n_131_104), .A (n_135_102), .B (n_141_99), .C1 (n_140_98), .C2 (n_134_101) );
AOI211_X1 g_129_105 (.ZN (n_129_105), .A (n_133_103), .B (n_139_100), .C1 (n_142_97), .C2 (n_136_100) );
AOI211_X1 g_127_104 (.ZN (n_127_104), .A (n_131_104), .B (n_137_101), .C1 (n_141_99), .C2 (n_138_99) );
AOI211_X1 g_125_105 (.ZN (n_125_105), .A (n_129_105), .B (n_135_102), .C1 (n_139_100), .C2 (n_140_98) );
AOI211_X1 g_123_106 (.ZN (n_123_106), .A (n_127_104), .B (n_133_103), .C1 (n_137_101), .C2 (n_142_97) );
AOI211_X1 g_121_107 (.ZN (n_121_107), .A (n_125_105), .B (n_131_104), .C1 (n_135_102), .C2 (n_141_99) );
AOI211_X1 g_119_108 (.ZN (n_119_108), .A (n_123_106), .B (n_129_105), .C1 (n_133_103), .C2 (n_139_100) );
AOI211_X1 g_117_109 (.ZN (n_117_109), .A (n_121_107), .B (n_127_104), .C1 (n_131_104), .C2 (n_137_101) );
AOI211_X1 g_115_110 (.ZN (n_115_110), .A (n_119_108), .B (n_125_105), .C1 (n_129_105), .C2 (n_135_102) );
AOI211_X1 g_113_111 (.ZN (n_113_111), .A (n_117_109), .B (n_123_106), .C1 (n_127_104), .C2 (n_133_103) );
AOI211_X1 g_111_112 (.ZN (n_111_112), .A (n_115_110), .B (n_121_107), .C1 (n_125_105), .C2 (n_131_104) );
AOI211_X1 g_109_113 (.ZN (n_109_113), .A (n_113_111), .B (n_119_108), .C1 (n_123_106), .C2 (n_129_105) );
AOI211_X1 g_107_114 (.ZN (n_107_114), .A (n_111_112), .B (n_117_109), .C1 (n_121_107), .C2 (n_127_104) );
AOI211_X1 g_105_115 (.ZN (n_105_115), .A (n_109_113), .B (n_115_110), .C1 (n_119_108), .C2 (n_125_105) );
AOI211_X1 g_103_116 (.ZN (n_103_116), .A (n_107_114), .B (n_113_111), .C1 (n_117_109), .C2 (n_123_106) );
AOI211_X1 g_101_117 (.ZN (n_101_117), .A (n_105_115), .B (n_111_112), .C1 (n_115_110), .C2 (n_121_107) );
AOI211_X1 g_99_118 (.ZN (n_99_118), .A (n_103_116), .B (n_109_113), .C1 (n_113_111), .C2 (n_119_108) );
AOI211_X1 g_97_119 (.ZN (n_97_119), .A (n_101_117), .B (n_107_114), .C1 (n_111_112), .C2 (n_117_109) );
AOI211_X1 g_95_120 (.ZN (n_95_120), .A (n_99_118), .B (n_105_115), .C1 (n_109_113), .C2 (n_115_110) );
AOI211_X1 g_93_121 (.ZN (n_93_121), .A (n_97_119), .B (n_103_116), .C1 (n_107_114), .C2 (n_113_111) );
AOI211_X1 g_91_122 (.ZN (n_91_122), .A (n_95_120), .B (n_101_117), .C1 (n_105_115), .C2 (n_111_112) );
AOI211_X1 g_89_123 (.ZN (n_89_123), .A (n_93_121), .B (n_99_118), .C1 (n_103_116), .C2 (n_109_113) );
AOI211_X1 g_87_124 (.ZN (n_87_124), .A (n_91_122), .B (n_97_119), .C1 (n_101_117), .C2 (n_107_114) );
AOI211_X1 g_85_125 (.ZN (n_85_125), .A (n_89_123), .B (n_95_120), .C1 (n_99_118), .C2 (n_105_115) );
AOI211_X1 g_86_127 (.ZN (n_86_127), .A (n_87_124), .B (n_93_121), .C1 (n_97_119), .C2 (n_103_116) );
AOI211_X1 g_84_126 (.ZN (n_84_126), .A (n_85_125), .B (n_91_122), .C1 (n_95_120), .C2 (n_101_117) );
AOI211_X1 g_86_125 (.ZN (n_86_125), .A (n_86_127), .B (n_89_123), .C1 (n_93_121), .C2 (n_99_118) );
AOI211_X1 g_88_124 (.ZN (n_88_124), .A (n_84_126), .B (n_87_124), .C1 (n_91_122), .C2 (n_97_119) );
AOI211_X1 g_90_123 (.ZN (n_90_123), .A (n_86_125), .B (n_85_125), .C1 (n_89_123), .C2 (n_95_120) );
AOI211_X1 g_92_122 (.ZN (n_92_122), .A (n_88_124), .B (n_86_127), .C1 (n_87_124), .C2 (n_93_121) );
AOI211_X1 g_94_121 (.ZN (n_94_121), .A (n_90_123), .B (n_84_126), .C1 (n_85_125), .C2 (n_91_122) );
AOI211_X1 g_96_120 (.ZN (n_96_120), .A (n_92_122), .B (n_86_125), .C1 (n_86_127), .C2 (n_89_123) );
AOI211_X1 g_98_119 (.ZN (n_98_119), .A (n_94_121), .B (n_88_124), .C1 (n_84_126), .C2 (n_87_124) );
AOI211_X1 g_100_118 (.ZN (n_100_118), .A (n_96_120), .B (n_90_123), .C1 (n_86_125), .C2 (n_85_125) );
AOI211_X1 g_102_117 (.ZN (n_102_117), .A (n_98_119), .B (n_92_122), .C1 (n_88_124), .C2 (n_86_127) );
AOI211_X1 g_104_116 (.ZN (n_104_116), .A (n_100_118), .B (n_94_121), .C1 (n_90_123), .C2 (n_84_126) );
AOI211_X1 g_106_115 (.ZN (n_106_115), .A (n_102_117), .B (n_96_120), .C1 (n_92_122), .C2 (n_86_125) );
AOI211_X1 g_108_114 (.ZN (n_108_114), .A (n_104_116), .B (n_98_119), .C1 (n_94_121), .C2 (n_88_124) );
AOI211_X1 g_110_113 (.ZN (n_110_113), .A (n_106_115), .B (n_100_118), .C1 (n_96_120), .C2 (n_90_123) );
AOI211_X1 g_112_112 (.ZN (n_112_112), .A (n_108_114), .B (n_102_117), .C1 (n_98_119), .C2 (n_92_122) );
AOI211_X1 g_111_114 (.ZN (n_111_114), .A (n_110_113), .B (n_104_116), .C1 (n_100_118), .C2 (n_94_121) );
AOI211_X1 g_110_112 (.ZN (n_110_112), .A (n_112_112), .B (n_106_115), .C1 (n_102_117), .C2 (n_96_120) );
AOI211_X1 g_112_111 (.ZN (n_112_111), .A (n_111_114), .B (n_108_114), .C1 (n_104_116), .C2 (n_98_119) );
AOI211_X1 g_114_110 (.ZN (n_114_110), .A (n_110_112), .B (n_110_113), .C1 (n_106_115), .C2 (n_100_118) );
AOI211_X1 g_116_109 (.ZN (n_116_109), .A (n_112_111), .B (n_112_112), .C1 (n_108_114), .C2 (n_102_117) );
AOI211_X1 g_118_108 (.ZN (n_118_108), .A (n_114_110), .B (n_111_114), .C1 (n_110_113), .C2 (n_104_116) );
AOI211_X1 g_117_110 (.ZN (n_117_110), .A (n_116_109), .B (n_110_112), .C1 (n_112_112), .C2 (n_106_115) );
AOI211_X1 g_119_109 (.ZN (n_119_109), .A (n_118_108), .B (n_112_111), .C1 (n_111_114), .C2 (n_108_114) );
AOI211_X1 g_121_108 (.ZN (n_121_108), .A (n_117_110), .B (n_114_110), .C1 (n_110_112), .C2 (n_110_113) );
AOI211_X1 g_123_107 (.ZN (n_123_107), .A (n_119_109), .B (n_116_109), .C1 (n_112_111), .C2 (n_112_112) );
AOI211_X1 g_125_106 (.ZN (n_125_106), .A (n_121_108), .B (n_118_108), .C1 (n_114_110), .C2 (n_111_114) );
AOI211_X1 g_127_105 (.ZN (n_127_105), .A (n_123_107), .B (n_117_110), .C1 (n_116_109), .C2 (n_110_112) );
AOI211_X1 g_129_104 (.ZN (n_129_104), .A (n_125_106), .B (n_119_109), .C1 (n_118_108), .C2 (n_112_111) );
AOI211_X1 g_131_103 (.ZN (n_131_103), .A (n_127_105), .B (n_121_108), .C1 (n_117_110), .C2 (n_114_110) );
AOI211_X1 g_133_102 (.ZN (n_133_102), .A (n_129_104), .B (n_123_107), .C1 (n_119_109), .C2 (n_116_109) );
AOI211_X1 g_135_101 (.ZN (n_135_101), .A (n_131_103), .B (n_125_106), .C1 (n_121_108), .C2 (n_118_108) );
AOI211_X1 g_137_100 (.ZN (n_137_100), .A (n_133_102), .B (n_127_105), .C1 (n_123_107), .C2 (n_117_110) );
AOI211_X1 g_139_99 (.ZN (n_139_99), .A (n_135_101), .B (n_129_104), .C1 (n_125_106), .C2 (n_119_109) );
AOI211_X1 g_140_101 (.ZN (n_140_101), .A (n_137_100), .B (n_131_103), .C1 (n_127_105), .C2 (n_121_108) );
AOI211_X1 g_138_102 (.ZN (n_138_102), .A (n_139_99), .B (n_133_102), .C1 (n_129_104), .C2 (n_123_107) );
AOI211_X1 g_136_103 (.ZN (n_136_103), .A (n_140_101), .B (n_135_101), .C1 (n_131_103), .C2 (n_125_106) );
AOI211_X1 g_134_104 (.ZN (n_134_104), .A (n_138_102), .B (n_137_100), .C1 (n_133_102), .C2 (n_127_105) );
AOI211_X1 g_132_105 (.ZN (n_132_105), .A (n_136_103), .B (n_139_99), .C1 (n_135_101), .C2 (n_129_104) );
AOI211_X1 g_130_106 (.ZN (n_130_106), .A (n_134_104), .B (n_140_101), .C1 (n_137_100), .C2 (n_131_103) );
AOI211_X1 g_128_105 (.ZN (n_128_105), .A (n_132_105), .B (n_138_102), .C1 (n_139_99), .C2 (n_133_102) );
AOI211_X1 g_126_106 (.ZN (n_126_106), .A (n_130_106), .B (n_136_103), .C1 (n_140_101), .C2 (n_135_101) );
AOI211_X1 g_124_107 (.ZN (n_124_107), .A (n_128_105), .B (n_134_104), .C1 (n_138_102), .C2 (n_137_100) );
AOI211_X1 g_122_108 (.ZN (n_122_108), .A (n_126_106), .B (n_132_105), .C1 (n_136_103), .C2 (n_139_99) );
AOI211_X1 g_120_109 (.ZN (n_120_109), .A (n_124_107), .B (n_130_106), .C1 (n_134_104), .C2 (n_140_101) );
AOI211_X1 g_118_110 (.ZN (n_118_110), .A (n_122_108), .B (n_128_105), .C1 (n_132_105), .C2 (n_138_102) );
AOI211_X1 g_116_111 (.ZN (n_116_111), .A (n_120_109), .B (n_126_106), .C1 (n_130_106), .C2 (n_136_103) );
AOI211_X1 g_114_112 (.ZN (n_114_112), .A (n_118_110), .B (n_124_107), .C1 (n_128_105), .C2 (n_134_104) );
AOI211_X1 g_112_113 (.ZN (n_112_113), .A (n_116_111), .B (n_122_108), .C1 (n_126_106), .C2 (n_132_105) );
AOI211_X1 g_110_114 (.ZN (n_110_114), .A (n_114_112), .B (n_120_109), .C1 (n_124_107), .C2 (n_130_106) );
AOI211_X1 g_108_113 (.ZN (n_108_113), .A (n_112_113), .B (n_118_110), .C1 (n_122_108), .C2 (n_128_105) );
AOI211_X1 g_106_114 (.ZN (n_106_114), .A (n_110_114), .B (n_116_111), .C1 (n_120_109), .C2 (n_126_106) );
AOI211_X1 g_108_115 (.ZN (n_108_115), .A (n_108_113), .B (n_114_112), .C1 (n_118_110), .C2 (n_124_107) );
AOI211_X1 g_106_116 (.ZN (n_106_116), .A (n_106_114), .B (n_112_113), .C1 (n_116_111), .C2 (n_122_108) );
AOI211_X1 g_104_117 (.ZN (n_104_117), .A (n_108_115), .B (n_110_114), .C1 (n_114_112), .C2 (n_120_109) );
AOI211_X1 g_102_118 (.ZN (n_102_118), .A (n_106_116), .B (n_108_113), .C1 (n_112_113), .C2 (n_118_110) );
AOI211_X1 g_100_119 (.ZN (n_100_119), .A (n_104_117), .B (n_106_114), .C1 (n_110_114), .C2 (n_116_111) );
AOI211_X1 g_98_120 (.ZN (n_98_120), .A (n_102_118), .B (n_108_115), .C1 (n_108_113), .C2 (n_114_112) );
AOI211_X1 g_96_121 (.ZN (n_96_121), .A (n_100_119), .B (n_106_116), .C1 (n_106_114), .C2 (n_112_113) );
AOI211_X1 g_94_122 (.ZN (n_94_122), .A (n_98_120), .B (n_104_117), .C1 (n_108_115), .C2 (n_110_114) );
AOI211_X1 g_92_123 (.ZN (n_92_123), .A (n_96_121), .B (n_102_118), .C1 (n_106_116), .C2 (n_108_113) );
AOI211_X1 g_90_124 (.ZN (n_90_124), .A (n_94_122), .B (n_100_119), .C1 (n_104_117), .C2 (n_106_114) );
AOI211_X1 g_88_125 (.ZN (n_88_125), .A (n_92_123), .B (n_98_120), .C1 (n_102_118), .C2 (n_108_115) );
AOI211_X1 g_86_126 (.ZN (n_86_126), .A (n_90_124), .B (n_96_121), .C1 (n_100_119), .C2 (n_106_116) );
AOI211_X1 g_84_125 (.ZN (n_84_125), .A (n_88_125), .B (n_94_122), .C1 (n_98_120), .C2 (n_104_117) );
AOI211_X1 g_82_126 (.ZN (n_82_126), .A (n_86_126), .B (n_92_123), .C1 (n_96_121), .C2 (n_102_118) );
AOI211_X1 g_80_127 (.ZN (n_80_127), .A (n_84_125), .B (n_90_124), .C1 (n_94_122), .C2 (n_100_119) );
AOI211_X1 g_78_128 (.ZN (n_78_128), .A (n_82_126), .B (n_88_125), .C1 (n_92_123), .C2 (n_98_120) );
AOI211_X1 g_79_126 (.ZN (n_79_126), .A (n_80_127), .B (n_86_126), .C1 (n_90_124), .C2 (n_96_121) );
AOI211_X1 g_77_127 (.ZN (n_77_127), .A (n_78_128), .B (n_84_125), .C1 (n_88_125), .C2 (n_94_122) );
AOI211_X1 g_75_128 (.ZN (n_75_128), .A (n_79_126), .B (n_82_126), .C1 (n_86_126), .C2 (n_92_123) );
AOI211_X1 g_73_129 (.ZN (n_73_129), .A (n_77_127), .B (n_80_127), .C1 (n_84_125), .C2 (n_90_124) );
AOI211_X1 g_71_130 (.ZN (n_71_130), .A (n_75_128), .B (n_78_128), .C1 (n_82_126), .C2 (n_88_125) );
AOI211_X1 g_69_131 (.ZN (n_69_131), .A (n_73_129), .B (n_79_126), .C1 (n_80_127), .C2 (n_86_126) );
AOI211_X1 g_67_132 (.ZN (n_67_132), .A (n_71_130), .B (n_77_127), .C1 (n_78_128), .C2 (n_84_125) );
AOI211_X1 g_65_133 (.ZN (n_65_133), .A (n_69_131), .B (n_75_128), .C1 (n_79_126), .C2 (n_82_126) );
AOI211_X1 g_63_134 (.ZN (n_63_134), .A (n_67_132), .B (n_73_129), .C1 (n_77_127), .C2 (n_80_127) );
AOI211_X1 g_61_135 (.ZN (n_61_135), .A (n_65_133), .B (n_71_130), .C1 (n_75_128), .C2 (n_78_128) );
AOI211_X1 g_59_136 (.ZN (n_59_136), .A (n_63_134), .B (n_69_131), .C1 (n_73_129), .C2 (n_79_126) );
AOI211_X1 g_60_134 (.ZN (n_60_134), .A (n_61_135), .B (n_67_132), .C1 (n_71_130), .C2 (n_77_127) );
AOI211_X1 g_58_135 (.ZN (n_58_135), .A (n_59_136), .B (n_65_133), .C1 (n_69_131), .C2 (n_75_128) );
AOI211_X1 g_56_136 (.ZN (n_56_136), .A (n_60_134), .B (n_63_134), .C1 (n_67_132), .C2 (n_73_129) );
AOI211_X1 g_54_137 (.ZN (n_54_137), .A (n_58_135), .B (n_61_135), .C1 (n_65_133), .C2 (n_71_130) );
AOI211_X1 g_52_138 (.ZN (n_52_138), .A (n_56_136), .B (n_59_136), .C1 (n_63_134), .C2 (n_69_131) );
AOI211_X1 g_50_139 (.ZN (n_50_139), .A (n_54_137), .B (n_60_134), .C1 (n_61_135), .C2 (n_67_132) );
AOI211_X1 g_48_140 (.ZN (n_48_140), .A (n_52_138), .B (n_58_135), .C1 (n_59_136), .C2 (n_65_133) );
AOI211_X1 g_46_141 (.ZN (n_46_141), .A (n_50_139), .B (n_56_136), .C1 (n_60_134), .C2 (n_63_134) );
AOI211_X1 g_44_140 (.ZN (n_44_140), .A (n_48_140), .B (n_54_137), .C1 (n_58_135), .C2 (n_61_135) );
AOI211_X1 g_42_141 (.ZN (n_42_141), .A (n_46_141), .B (n_52_138), .C1 (n_56_136), .C2 (n_59_136) );
AOI211_X1 g_40_142 (.ZN (n_40_142), .A (n_44_140), .B (n_50_139), .C1 (n_54_137), .C2 (n_60_134) );
AOI211_X1 g_38_143 (.ZN (n_38_143), .A (n_42_141), .B (n_48_140), .C1 (n_52_138), .C2 (n_58_135) );
AOI211_X1 g_37_145 (.ZN (n_37_145), .A (n_40_142), .B (n_46_141), .C1 (n_50_139), .C2 (n_56_136) );
AOI211_X1 g_36_147 (.ZN (n_36_147), .A (n_38_143), .B (n_44_140), .C1 (n_48_140), .C2 (n_54_137) );
AOI211_X1 g_34_146 (.ZN (n_34_146), .A (n_37_145), .B (n_42_141), .C1 (n_46_141), .C2 (n_52_138) );
AOI211_X1 g_33_148 (.ZN (n_33_148), .A (n_36_147), .B (n_40_142), .C1 (n_44_140), .C2 (n_50_139) );
AOI211_X1 g_34_150 (.ZN (n_34_150), .A (n_34_146), .B (n_38_143), .C1 (n_42_141), .C2 (n_48_140) );
AOI211_X1 g_35_148 (.ZN (n_35_148), .A (n_33_148), .B (n_37_145), .C1 (n_40_142), .C2 (n_46_141) );
AOI211_X1 g_37_147 (.ZN (n_37_147), .A (n_34_150), .B (n_36_147), .C1 (n_38_143), .C2 (n_44_140) );
AOI211_X1 g_36_145 (.ZN (n_36_145), .A (n_35_148), .B (n_34_146), .C1 (n_37_145), .C2 (n_42_141) );
AOI211_X1 g_35_147 (.ZN (n_35_147), .A (n_37_147), .B (n_33_148), .C1 (n_36_147), .C2 (n_40_142) );
AOI211_X1 g_36_149 (.ZN (n_36_149), .A (n_36_145), .B (n_34_150), .C1 (n_34_146), .C2 (n_38_143) );
AOI211_X1 g_38_150 (.ZN (n_38_150), .A (n_35_147), .B (n_35_148), .C1 (n_33_148), .C2 (n_37_145) );
AOI211_X1 g_37_148 (.ZN (n_37_148), .A (n_36_149), .B (n_37_147), .C1 (n_34_150), .C2 (n_36_147) );
AOI211_X1 g_38_146 (.ZN (n_38_146), .A (n_38_150), .B (n_36_145), .C1 (n_35_148), .C2 (n_34_146) );
AOI211_X1 g_39_148 (.ZN (n_39_148), .A (n_37_148), .B (n_35_147), .C1 (n_37_147), .C2 (n_33_148) );
AOI211_X1 g_40_146 (.ZN (n_40_146), .A (n_38_146), .B (n_36_149), .C1 (n_36_145), .C2 (n_34_150) );
AOI211_X1 g_39_144 (.ZN (n_39_144), .A (n_39_148), .B (n_38_150), .C1 (n_35_147), .C2 (n_35_148) );
AOI211_X1 g_41_143 (.ZN (n_41_143), .A (n_40_146), .B (n_37_148), .C1 (n_36_149), .C2 (n_37_147) );
AOI211_X1 g_43_142 (.ZN (n_43_142), .A (n_39_144), .B (n_38_146), .C1 (n_38_150), .C2 (n_36_145) );
AOI211_X1 g_45_141 (.ZN (n_45_141), .A (n_41_143), .B (n_39_148), .C1 (n_37_148), .C2 (n_35_147) );
AOI211_X1 g_47_140 (.ZN (n_47_140), .A (n_43_142), .B (n_40_146), .C1 (n_38_146), .C2 (n_36_149) );
AOI211_X1 g_49_139 (.ZN (n_49_139), .A (n_45_141), .B (n_39_144), .C1 (n_39_148), .C2 (n_38_150) );
AOI211_X1 g_51_138 (.ZN (n_51_138), .A (n_47_140), .B (n_41_143), .C1 (n_40_146), .C2 (n_37_148) );
AOI211_X1 g_53_137 (.ZN (n_53_137), .A (n_49_139), .B (n_43_142), .C1 (n_39_144), .C2 (n_38_146) );
AOI211_X1 g_52_139 (.ZN (n_52_139), .A (n_51_138), .B (n_45_141), .C1 (n_41_143), .C2 (n_39_148) );
AOI211_X1 g_54_138 (.ZN (n_54_138), .A (n_53_137), .B (n_47_140), .C1 (n_43_142), .C2 (n_40_146) );
AOI211_X1 g_56_137 (.ZN (n_56_137), .A (n_52_139), .B (n_49_139), .C1 (n_45_141), .C2 (n_39_144) );
AOI211_X1 g_58_136 (.ZN (n_58_136), .A (n_54_138), .B (n_51_138), .C1 (n_47_140), .C2 (n_41_143) );
AOI211_X1 g_60_135 (.ZN (n_60_135), .A (n_56_137), .B (n_53_137), .C1 (n_49_139), .C2 (n_43_142) );
AOI211_X1 g_62_134 (.ZN (n_62_134), .A (n_58_136), .B (n_52_139), .C1 (n_51_138), .C2 (n_45_141) );
AOI211_X1 g_64_133 (.ZN (n_64_133), .A (n_60_135), .B (n_54_138), .C1 (n_53_137), .C2 (n_47_140) );
AOI211_X1 g_66_132 (.ZN (n_66_132), .A (n_62_134), .B (n_56_137), .C1 (n_52_139), .C2 (n_49_139) );
AOI211_X1 g_68_131 (.ZN (n_68_131), .A (n_64_133), .B (n_58_136), .C1 (n_54_138), .C2 (n_51_138) );
AOI211_X1 g_70_130 (.ZN (n_70_130), .A (n_66_132), .B (n_60_135), .C1 (n_56_137), .C2 (n_53_137) );
AOI211_X1 g_72_129 (.ZN (n_72_129), .A (n_68_131), .B (n_62_134), .C1 (n_58_136), .C2 (n_52_139) );
AOI211_X1 g_74_128 (.ZN (n_74_128), .A (n_70_130), .B (n_64_133), .C1 (n_60_135), .C2 (n_54_138) );
AOI211_X1 g_76_127 (.ZN (n_76_127), .A (n_72_129), .B (n_66_132), .C1 (n_62_134), .C2 (n_56_137) );
AOI211_X1 g_77_129 (.ZN (n_77_129), .A (n_74_128), .B (n_68_131), .C1 (n_64_133), .C2 (n_58_136) );
AOI211_X1 g_75_130 (.ZN (n_75_130), .A (n_76_127), .B (n_70_130), .C1 (n_66_132), .C2 (n_60_135) );
AOI211_X1 g_73_131 (.ZN (n_73_131), .A (n_77_129), .B (n_72_129), .C1 (n_68_131), .C2 (n_62_134) );
AOI211_X1 g_71_132 (.ZN (n_71_132), .A (n_75_130), .B (n_74_128), .C1 (n_70_130), .C2 (n_64_133) );
AOI211_X1 g_69_133 (.ZN (n_69_133), .A (n_73_131), .B (n_76_127), .C1 (n_72_129), .C2 (n_66_132) );
AOI211_X1 g_70_131 (.ZN (n_70_131), .A (n_71_132), .B (n_77_129), .C1 (n_74_128), .C2 (n_68_131) );
AOI211_X1 g_68_132 (.ZN (n_68_132), .A (n_69_133), .B (n_75_130), .C1 (n_76_127), .C2 (n_70_130) );
AOI211_X1 g_66_133 (.ZN (n_66_133), .A (n_70_131), .B (n_73_131), .C1 (n_77_129), .C2 (n_72_129) );
AOI211_X1 g_64_134 (.ZN (n_64_134), .A (n_68_132), .B (n_71_132), .C1 (n_75_130), .C2 (n_74_128) );
AOI211_X1 g_65_132 (.ZN (n_65_132), .A (n_66_133), .B (n_69_133), .C1 (n_73_131), .C2 (n_76_127) );
AOI211_X1 g_63_133 (.ZN (n_63_133), .A (n_64_134), .B (n_70_131), .C1 (n_71_132), .C2 (n_77_129) );
AOI211_X1 g_61_134 (.ZN (n_61_134), .A (n_65_132), .B (n_68_132), .C1 (n_69_133), .C2 (n_75_130) );
AOI211_X1 g_59_135 (.ZN (n_59_135), .A (n_63_133), .B (n_66_133), .C1 (n_70_131), .C2 (n_73_131) );
AOI211_X1 g_57_136 (.ZN (n_57_136), .A (n_61_134), .B (n_64_134), .C1 (n_68_132), .C2 (n_71_132) );
AOI211_X1 g_55_137 (.ZN (n_55_137), .A (n_59_135), .B (n_65_132), .C1 (n_66_133), .C2 (n_69_133) );
AOI211_X1 g_53_138 (.ZN (n_53_138), .A (n_57_136), .B (n_63_133), .C1 (n_64_134), .C2 (n_70_131) );
AOI211_X1 g_51_139 (.ZN (n_51_139), .A (n_55_137), .B (n_61_134), .C1 (n_65_132), .C2 (n_68_132) );
AOI211_X1 g_49_140 (.ZN (n_49_140), .A (n_53_138), .B (n_59_135), .C1 (n_63_133), .C2 (n_66_133) );
AOI211_X1 g_47_141 (.ZN (n_47_141), .A (n_51_139), .B (n_57_136), .C1 (n_61_134), .C2 (n_64_134) );
AOI211_X1 g_45_142 (.ZN (n_45_142), .A (n_49_140), .B (n_55_137), .C1 (n_59_135), .C2 (n_65_132) );
AOI211_X1 g_43_143 (.ZN (n_43_143), .A (n_47_141), .B (n_53_138), .C1 (n_57_136), .C2 (n_63_133) );
AOI211_X1 g_41_144 (.ZN (n_41_144), .A (n_45_142), .B (n_51_139), .C1 (n_55_137), .C2 (n_61_134) );
AOI211_X1 g_39_145 (.ZN (n_39_145), .A (n_43_143), .B (n_49_140), .C1 (n_53_138), .C2 (n_59_135) );
AOI211_X1 g_37_146 (.ZN (n_37_146), .A (n_41_144), .B (n_47_141), .C1 (n_51_139), .C2 (n_57_136) );
AOI211_X1 g_38_148 (.ZN (n_38_148), .A (n_39_145), .B (n_45_142), .C1 (n_49_140), .C2 (n_55_137) );
AOI211_X1 g_40_147 (.ZN (n_40_147), .A (n_37_146), .B (n_43_143), .C1 (n_47_141), .C2 (n_53_138) );
AOI211_X1 g_41_145 (.ZN (n_41_145), .A (n_38_148), .B (n_41_144), .C1 (n_45_142), .C2 (n_51_139) );
AOI211_X1 g_39_146 (.ZN (n_39_146), .A (n_40_147), .B (n_39_145), .C1 (n_43_143), .C2 (n_49_140) );
AOI211_X1 g_40_144 (.ZN (n_40_144), .A (n_41_145), .B (n_37_146), .C1 (n_41_144), .C2 (n_47_141) );
AOI211_X1 g_38_145 (.ZN (n_38_145), .A (n_39_146), .B (n_38_148), .C1 (n_39_145), .C2 (n_45_142) );
AOI211_X1 g_39_147 (.ZN (n_39_147), .A (n_40_144), .B (n_40_147), .C1 (n_37_146), .C2 (n_43_143) );
AOI211_X1 g_40_145 (.ZN (n_40_145), .A (n_38_145), .B (n_41_145), .C1 (n_38_148), .C2 (n_41_144) );
AOI211_X1 g_42_144 (.ZN (n_42_144), .A (n_39_147), .B (n_39_146), .C1 (n_40_147), .C2 (n_39_145) );
AOI211_X1 g_41_146 (.ZN (n_41_146), .A (n_40_145), .B (n_40_144), .C1 (n_41_145), .C2 (n_37_146) );
AOI211_X1 g_42_148 (.ZN (n_42_148), .A (n_42_144), .B (n_38_145), .C1 (n_39_146), .C2 (n_38_148) );
AOI211_X1 g_40_149 (.ZN (n_40_149), .A (n_41_146), .B (n_39_147), .C1 (n_40_144), .C2 (n_40_147) );
AOI211_X1 g_41_147 (.ZN (n_41_147), .A (n_42_148), .B (n_40_145), .C1 (n_38_145), .C2 (n_41_145) );
AOI211_X1 g_43_146 (.ZN (n_43_146), .A (n_40_149), .B (n_42_144), .C1 (n_39_147), .C2 (n_39_146) );
AOI211_X1 g_44_144 (.ZN (n_44_144), .A (n_41_147), .B (n_41_146), .C1 (n_40_145), .C2 (n_40_144) );
AOI211_X1 g_42_143 (.ZN (n_42_143), .A (n_43_146), .B (n_42_148), .C1 (n_42_144), .C2 (n_38_145) );
AOI211_X1 g_44_142 (.ZN (n_44_142), .A (n_44_144), .B (n_40_149), .C1 (n_41_146), .C2 (n_39_147) );
AOI211_X1 g_43_144 (.ZN (n_43_144), .A (n_42_143), .B (n_41_147), .C1 (n_42_148), .C2 (n_40_145) );
AOI211_X1 g_45_143 (.ZN (n_45_143), .A (n_44_142), .B (n_43_146), .C1 (n_40_149), .C2 (n_42_144) );
AOI211_X1 g_47_142 (.ZN (n_47_142), .A (n_43_144), .B (n_44_144), .C1 (n_41_147), .C2 (n_41_146) );
AOI211_X1 g_49_141 (.ZN (n_49_141), .A (n_45_143), .B (n_42_143), .C1 (n_43_146), .C2 (n_42_148) );
AOI211_X1 g_51_140 (.ZN (n_51_140), .A (n_47_142), .B (n_44_142), .C1 (n_44_144), .C2 (n_40_149) );
AOI211_X1 g_53_139 (.ZN (n_53_139), .A (n_49_141), .B (n_43_144), .C1 (n_42_143), .C2 (n_41_147) );
AOI211_X1 g_55_138 (.ZN (n_55_138), .A (n_51_140), .B (n_45_143), .C1 (n_44_142), .C2 (n_43_146) );
AOI211_X1 g_57_137 (.ZN (n_57_137), .A (n_53_139), .B (n_47_142), .C1 (n_43_144), .C2 (n_44_144) );
AOI211_X1 g_56_139 (.ZN (n_56_139), .A (n_55_138), .B (n_49_141), .C1 (n_45_143), .C2 (n_42_143) );
AOI211_X1 g_58_138 (.ZN (n_58_138), .A (n_57_137), .B (n_51_140), .C1 (n_47_142), .C2 (n_44_142) );
AOI211_X1 g_60_137 (.ZN (n_60_137), .A (n_56_139), .B (n_53_139), .C1 (n_49_141), .C2 (n_43_144) );
AOI211_X1 g_62_136 (.ZN (n_62_136), .A (n_58_138), .B (n_55_138), .C1 (n_51_140), .C2 (n_45_143) );
AOI211_X1 g_64_135 (.ZN (n_64_135), .A (n_60_137), .B (n_57_137), .C1 (n_53_139), .C2 (n_47_142) );
AOI211_X1 g_66_134 (.ZN (n_66_134), .A (n_62_136), .B (n_56_139), .C1 (n_55_138), .C2 (n_49_141) );
AOI211_X1 g_68_133 (.ZN (n_68_133), .A (n_64_135), .B (n_58_138), .C1 (n_57_137), .C2 (n_51_140) );
AOI211_X1 g_70_132 (.ZN (n_70_132), .A (n_66_134), .B (n_60_137), .C1 (n_56_139), .C2 (n_53_139) );
AOI211_X1 g_72_131 (.ZN (n_72_131), .A (n_68_133), .B (n_62_136), .C1 (n_58_138), .C2 (n_55_138) );
AOI211_X1 g_74_130 (.ZN (n_74_130), .A (n_70_132), .B (n_64_135), .C1 (n_60_137), .C2 (n_57_137) );
AOI211_X1 g_76_129 (.ZN (n_76_129), .A (n_72_131), .B (n_66_134), .C1 (n_62_136), .C2 (n_56_139) );
AOI211_X1 g_75_131 (.ZN (n_75_131), .A (n_74_130), .B (n_68_133), .C1 (n_64_135), .C2 (n_58_138) );
AOI211_X1 g_73_130 (.ZN (n_73_130), .A (n_76_129), .B (n_70_132), .C1 (n_66_134), .C2 (n_60_137) );
AOI211_X1 g_75_129 (.ZN (n_75_129), .A (n_75_131), .B (n_72_131), .C1 (n_68_133), .C2 (n_62_136) );
AOI211_X1 g_77_128 (.ZN (n_77_128), .A (n_73_130), .B (n_74_130), .C1 (n_70_132), .C2 (n_64_135) );
AOI211_X1 g_79_127 (.ZN (n_79_127), .A (n_75_129), .B (n_76_129), .C1 (n_72_131), .C2 (n_66_134) );
AOI211_X1 g_81_126 (.ZN (n_81_126), .A (n_77_128), .B (n_75_131), .C1 (n_74_130), .C2 (n_68_133) );
AOI211_X1 g_83_125 (.ZN (n_83_125), .A (n_79_127), .B (n_73_130), .C1 (n_76_129), .C2 (n_70_132) );
AOI211_X1 g_82_127 (.ZN (n_82_127), .A (n_81_126), .B (n_75_129), .C1 (n_75_131), .C2 (n_72_131) );
AOI211_X1 g_80_128 (.ZN (n_80_128), .A (n_83_125), .B (n_77_128), .C1 (n_73_130), .C2 (n_74_130) );
AOI211_X1 g_78_129 (.ZN (n_78_129), .A (n_82_127), .B (n_79_127), .C1 (n_75_129), .C2 (n_76_129) );
AOI211_X1 g_76_130 (.ZN (n_76_130), .A (n_80_128), .B (n_81_126), .C1 (n_77_128), .C2 (n_75_131) );
AOI211_X1 g_74_131 (.ZN (n_74_131), .A (n_78_129), .B (n_83_125), .C1 (n_79_127), .C2 (n_73_130) );
AOI211_X1 g_72_132 (.ZN (n_72_132), .A (n_76_130), .B (n_82_127), .C1 (n_81_126), .C2 (n_75_129) );
AOI211_X1 g_70_133 (.ZN (n_70_133), .A (n_74_131), .B (n_80_128), .C1 (n_83_125), .C2 (n_77_128) );
AOI211_X1 g_71_131 (.ZN (n_71_131), .A (n_72_132), .B (n_78_129), .C1 (n_82_127), .C2 (n_79_127) );
AOI211_X1 g_69_132 (.ZN (n_69_132), .A (n_70_133), .B (n_76_130), .C1 (n_80_128), .C2 (n_81_126) );
AOI211_X1 g_67_133 (.ZN (n_67_133), .A (n_71_131), .B (n_74_131), .C1 (n_78_129), .C2 (n_83_125) );
AOI211_X1 g_65_134 (.ZN (n_65_134), .A (n_69_132), .B (n_72_132), .C1 (n_76_130), .C2 (n_82_127) );
AOI211_X1 g_63_135 (.ZN (n_63_135), .A (n_67_133), .B (n_70_133), .C1 (n_74_131), .C2 (n_80_128) );
AOI211_X1 g_61_136 (.ZN (n_61_136), .A (n_65_134), .B (n_71_131), .C1 (n_72_132), .C2 (n_78_129) );
AOI211_X1 g_59_137 (.ZN (n_59_137), .A (n_63_135), .B (n_69_132), .C1 (n_70_133), .C2 (n_76_130) );
AOI211_X1 g_57_138 (.ZN (n_57_138), .A (n_61_136), .B (n_67_133), .C1 (n_71_131), .C2 (n_74_131) );
AOI211_X1 g_55_139 (.ZN (n_55_139), .A (n_59_137), .B (n_65_134), .C1 (n_69_132), .C2 (n_72_132) );
AOI211_X1 g_53_140 (.ZN (n_53_140), .A (n_57_138), .B (n_63_135), .C1 (n_67_133), .C2 (n_70_133) );
AOI211_X1 g_51_141 (.ZN (n_51_141), .A (n_55_139), .B (n_61_136), .C1 (n_65_134), .C2 (n_71_131) );
AOI211_X1 g_49_142 (.ZN (n_49_142), .A (n_53_140), .B (n_59_137), .C1 (n_63_135), .C2 (n_69_132) );
AOI211_X1 g_50_140 (.ZN (n_50_140), .A (n_51_141), .B (n_57_138), .C1 (n_61_136), .C2 (n_67_133) );
AOI211_X1 g_48_141 (.ZN (n_48_141), .A (n_49_142), .B (n_55_139), .C1 (n_59_137), .C2 (n_65_134) );
AOI211_X1 g_46_142 (.ZN (n_46_142), .A (n_50_140), .B (n_53_140), .C1 (n_57_138), .C2 (n_63_135) );
AOI211_X1 g_44_143 (.ZN (n_44_143), .A (n_48_141), .B (n_51_141), .C1 (n_55_139), .C2 (n_61_136) );
AOI211_X1 g_43_145 (.ZN (n_43_145), .A (n_46_142), .B (n_49_142), .C1 (n_53_140), .C2 (n_59_137) );
AOI211_X1 g_45_144 (.ZN (n_45_144), .A (n_44_143), .B (n_50_140), .C1 (n_51_141), .C2 (n_57_138) );
AOI211_X1 g_47_143 (.ZN (n_47_143), .A (n_43_145), .B (n_48_141), .C1 (n_49_142), .C2 (n_55_139) );
AOI211_X1 g_46_145 (.ZN (n_46_145), .A (n_45_144), .B (n_46_142), .C1 (n_50_140), .C2 (n_53_140) );
AOI211_X1 g_44_146 (.ZN (n_44_146), .A (n_47_143), .B (n_44_143), .C1 (n_48_141), .C2 (n_51_141) );
AOI211_X1 g_42_145 (.ZN (n_42_145), .A (n_46_145), .B (n_43_145), .C1 (n_46_142), .C2 (n_49_142) );
AOI211_X1 g_43_147 (.ZN (n_43_147), .A (n_44_146), .B (n_45_144), .C1 (n_44_143), .C2 (n_50_140) );
AOI211_X1 g_41_148 (.ZN (n_41_148), .A (n_42_145), .B (n_47_143), .C1 (n_43_145), .C2 (n_48_141) );
AOI211_X1 g_42_150 (.ZN (n_42_150), .A (n_43_147), .B (n_46_145), .C1 (n_45_144), .C2 (n_46_142) );
AOI211_X1 g_43_148 (.ZN (n_43_148), .A (n_41_148), .B (n_44_146), .C1 (n_47_143), .C2 (n_44_143) );
AOI211_X1 g_42_146 (.ZN (n_42_146), .A (n_42_150), .B (n_42_145), .C1 (n_46_145), .C2 (n_43_145) );
AOI211_X1 g_44_145 (.ZN (n_44_145), .A (n_43_148), .B (n_43_147), .C1 (n_44_146), .C2 (n_45_144) );
AOI211_X1 g_45_147 (.ZN (n_45_147), .A (n_42_146), .B (n_41_148), .C1 (n_42_145), .C2 (n_47_143) );
AOI211_X1 g_44_149 (.ZN (n_44_149), .A (n_44_145), .B (n_42_150), .C1 (n_43_147), .C2 (n_46_145) );
AOI211_X1 g_46_150 (.ZN (n_46_150), .A (n_45_147), .B (n_43_148), .C1 (n_41_148), .C2 (n_44_146) );
AOI211_X1 g_45_148 (.ZN (n_45_148), .A (n_44_149), .B (n_42_146), .C1 (n_42_150), .C2 (n_42_145) );
AOI211_X1 g_47_147 (.ZN (n_47_147), .A (n_46_150), .B (n_44_145), .C1 (n_43_148), .C2 (n_43_147) );
AOI211_X1 g_45_146 (.ZN (n_45_146), .A (n_45_148), .B (n_45_147), .C1 (n_42_146), .C2 (n_41_148) );
AOI211_X1 g_46_144 (.ZN (n_46_144), .A (n_47_147), .B (n_44_149), .C1 (n_44_145), .C2 (n_42_150) );
AOI211_X1 g_48_143 (.ZN (n_48_143), .A (n_45_146), .B (n_46_150), .C1 (n_45_147), .C2 (n_43_148) );
AOI211_X1 g_50_142 (.ZN (n_50_142), .A (n_46_144), .B (n_45_148), .C1 (n_44_149), .C2 (n_42_146) );
AOI211_X1 g_52_141 (.ZN (n_52_141), .A (n_48_143), .B (n_47_147), .C1 (n_46_150), .C2 (n_44_145) );
AOI211_X1 g_54_140 (.ZN (n_54_140), .A (n_50_142), .B (n_45_146), .C1 (n_45_148), .C2 (n_45_147) );
AOI211_X1 g_53_142 (.ZN (n_53_142), .A (n_52_141), .B (n_46_144), .C1 (n_47_147), .C2 (n_44_149) );
AOI211_X1 g_52_140 (.ZN (n_52_140), .A (n_54_140), .B (n_48_143), .C1 (n_45_146), .C2 (n_46_150) );
AOI211_X1 g_54_139 (.ZN (n_54_139), .A (n_53_142), .B (n_50_142), .C1 (n_46_144), .C2 (n_45_148) );
AOI211_X1 g_56_138 (.ZN (n_56_138), .A (n_52_140), .B (n_52_141), .C1 (n_48_143), .C2 (n_47_147) );
AOI211_X1 g_58_137 (.ZN (n_58_137), .A (n_54_139), .B (n_54_140), .C1 (n_50_142), .C2 (n_45_146) );
AOI211_X1 g_60_136 (.ZN (n_60_136), .A (n_56_138), .B (n_53_142), .C1 (n_52_141), .C2 (n_46_144) );
AOI211_X1 g_62_135 (.ZN (n_62_135), .A (n_58_137), .B (n_52_140), .C1 (n_54_140), .C2 (n_48_143) );
AOI211_X1 g_61_137 (.ZN (n_61_137), .A (n_60_136), .B (n_54_139), .C1 (n_53_142), .C2 (n_50_142) );
AOI211_X1 g_63_136 (.ZN (n_63_136), .A (n_62_135), .B (n_56_138), .C1 (n_52_140), .C2 (n_52_141) );
AOI211_X1 g_65_135 (.ZN (n_65_135), .A (n_61_137), .B (n_58_137), .C1 (n_54_139), .C2 (n_54_140) );
AOI211_X1 g_67_134 (.ZN (n_67_134), .A (n_63_136), .B (n_60_136), .C1 (n_56_138), .C2 (n_53_142) );
AOI211_X1 g_66_136 (.ZN (n_66_136), .A (n_65_135), .B (n_62_135), .C1 (n_58_137), .C2 (n_52_140) );
AOI211_X1 g_68_135 (.ZN (n_68_135), .A (n_67_134), .B (n_61_137), .C1 (n_60_136), .C2 (n_54_139) );
AOI211_X1 g_70_134 (.ZN (n_70_134), .A (n_66_136), .B (n_63_136), .C1 (n_62_135), .C2 (n_56_138) );
AOI211_X1 g_72_133 (.ZN (n_72_133), .A (n_68_135), .B (n_65_135), .C1 (n_61_137), .C2 (n_58_137) );
AOI211_X1 g_74_132 (.ZN (n_74_132), .A (n_70_134), .B (n_67_134), .C1 (n_63_136), .C2 (n_60_136) );
AOI211_X1 g_76_131 (.ZN (n_76_131), .A (n_72_133), .B (n_66_136), .C1 (n_65_135), .C2 (n_62_135) );
AOI211_X1 g_78_130 (.ZN (n_78_130), .A (n_74_132), .B (n_68_135), .C1 (n_67_134), .C2 (n_61_137) );
AOI211_X1 g_80_129 (.ZN (n_80_129), .A (n_76_131), .B (n_70_134), .C1 (n_66_136), .C2 (n_63_136) );
AOI211_X1 g_81_127 (.ZN (n_81_127), .A (n_78_130), .B (n_72_133), .C1 (n_68_135), .C2 (n_65_135) );
AOI211_X1 g_83_128 (.ZN (n_83_128), .A (n_80_129), .B (n_74_132), .C1 (n_70_134), .C2 (n_67_134) );
AOI211_X1 g_85_127 (.ZN (n_85_127), .A (n_81_127), .B (n_76_131), .C1 (n_72_133), .C2 (n_66_136) );
AOI211_X1 g_87_126 (.ZN (n_87_126), .A (n_83_128), .B (n_78_130), .C1 (n_74_132), .C2 (n_68_135) );
AOI211_X1 g_89_125 (.ZN (n_89_125), .A (n_85_127), .B (n_80_129), .C1 (n_76_131), .C2 (n_70_134) );
AOI211_X1 g_91_124 (.ZN (n_91_124), .A (n_87_126), .B (n_81_127), .C1 (n_78_130), .C2 (n_72_133) );
AOI211_X1 g_93_123 (.ZN (n_93_123), .A (n_89_125), .B (n_83_128), .C1 (n_80_129), .C2 (n_74_132) );
AOI211_X1 g_95_122 (.ZN (n_95_122), .A (n_91_124), .B (n_85_127), .C1 (n_81_127), .C2 (n_76_131) );
AOI211_X1 g_97_121 (.ZN (n_97_121), .A (n_93_123), .B (n_87_126), .C1 (n_83_128), .C2 (n_78_130) );
AOI211_X1 g_99_120 (.ZN (n_99_120), .A (n_95_122), .B (n_89_125), .C1 (n_85_127), .C2 (n_80_129) );
AOI211_X1 g_101_119 (.ZN (n_101_119), .A (n_97_121), .B (n_91_124), .C1 (n_87_126), .C2 (n_81_127) );
AOI211_X1 g_103_118 (.ZN (n_103_118), .A (n_99_120), .B (n_93_123), .C1 (n_89_125), .C2 (n_83_128) );
AOI211_X1 g_105_117 (.ZN (n_105_117), .A (n_101_119), .B (n_95_122), .C1 (n_91_124), .C2 (n_85_127) );
AOI211_X1 g_107_116 (.ZN (n_107_116), .A (n_103_118), .B (n_97_121), .C1 (n_93_123), .C2 (n_87_126) );
AOI211_X1 g_109_115 (.ZN (n_109_115), .A (n_105_117), .B (n_99_120), .C1 (n_95_122), .C2 (n_89_125) );
AOI211_X1 g_108_117 (.ZN (n_108_117), .A (n_107_116), .B (n_101_119), .C1 (n_97_121), .C2 (n_91_124) );
AOI211_X1 g_107_115 (.ZN (n_107_115), .A (n_109_115), .B (n_103_118), .C1 (n_99_120), .C2 (n_93_123) );
AOI211_X1 g_109_114 (.ZN (n_109_114), .A (n_108_117), .B (n_105_117), .C1 (n_101_119), .C2 (n_95_122) );
AOI211_X1 g_111_113 (.ZN (n_111_113), .A (n_107_115), .B (n_107_116), .C1 (n_103_118), .C2 (n_97_121) );
AOI211_X1 g_113_112 (.ZN (n_113_112), .A (n_109_114), .B (n_109_115), .C1 (n_105_117), .C2 (n_99_120) );
AOI211_X1 g_115_111 (.ZN (n_115_111), .A (n_111_113), .B (n_108_117), .C1 (n_107_116), .C2 (n_101_119) );
AOI211_X1 g_114_113 (.ZN (n_114_113), .A (n_113_112), .B (n_107_115), .C1 (n_109_115), .C2 (n_103_118) );
AOI211_X1 g_116_112 (.ZN (n_116_112), .A (n_115_111), .B (n_109_114), .C1 (n_108_117), .C2 (n_105_117) );
AOI211_X1 g_118_111 (.ZN (n_118_111), .A (n_114_113), .B (n_111_113), .C1 (n_107_115), .C2 (n_107_116) );
AOI211_X1 g_120_110 (.ZN (n_120_110), .A (n_116_112), .B (n_113_112), .C1 (n_109_114), .C2 (n_109_115) );
AOI211_X1 g_122_109 (.ZN (n_122_109), .A (n_118_111), .B (n_115_111), .C1 (n_111_113), .C2 (n_108_117) );
AOI211_X1 g_124_108 (.ZN (n_124_108), .A (n_120_110), .B (n_114_113), .C1 (n_113_112), .C2 (n_107_115) );
AOI211_X1 g_126_107 (.ZN (n_126_107), .A (n_122_109), .B (n_116_112), .C1 (n_115_111), .C2 (n_109_114) );
AOI211_X1 g_128_106 (.ZN (n_128_106), .A (n_124_108), .B (n_118_111), .C1 (n_114_113), .C2 (n_111_113) );
AOI211_X1 g_130_105 (.ZN (n_130_105), .A (n_126_107), .B (n_120_110), .C1 (n_116_112), .C2 (n_113_112) );
AOI211_X1 g_132_104 (.ZN (n_132_104), .A (n_128_106), .B (n_122_109), .C1 (n_118_111), .C2 (n_115_111) );
AOI211_X1 g_134_103 (.ZN (n_134_103), .A (n_130_105), .B (n_124_108), .C1 (n_120_110), .C2 (n_114_113) );
AOI211_X1 g_136_102 (.ZN (n_136_102), .A (n_132_104), .B (n_126_107), .C1 (n_122_109), .C2 (n_116_112) );
AOI211_X1 g_138_101 (.ZN (n_138_101), .A (n_134_103), .B (n_128_106), .C1 (n_124_108), .C2 (n_118_111) );
AOI211_X1 g_140_100 (.ZN (n_140_100), .A (n_136_102), .B (n_130_105), .C1 (n_126_107), .C2 (n_120_110) );
AOI211_X1 g_142_99 (.ZN (n_142_99), .A (n_138_101), .B (n_132_104), .C1 (n_128_106), .C2 (n_122_109) );
AOI211_X1 g_144_98 (.ZN (n_144_98), .A (n_140_100), .B (n_134_103), .C1 (n_130_105), .C2 (n_124_108) );
AOI211_X1 g_146_99 (.ZN (n_146_99), .A (n_142_99), .B (n_136_102), .C1 (n_132_104), .C2 (n_126_107) );
AOI211_X1 g_144_100 (.ZN (n_144_100), .A (n_144_98), .B (n_138_101), .C1 (n_134_103), .C2 (n_128_106) );
AOI211_X1 g_142_101 (.ZN (n_142_101), .A (n_146_99), .B (n_140_100), .C1 (n_136_102), .C2 (n_130_105) );
AOI211_X1 g_143_99 (.ZN (n_143_99), .A (n_144_100), .B (n_142_99), .C1 (n_138_101), .C2 (n_132_104) );
AOI211_X1 g_144_101 (.ZN (n_144_101), .A (n_142_101), .B (n_144_98), .C1 (n_140_100), .C2 (n_134_103) );
AOI211_X1 g_146_102 (.ZN (n_146_102), .A (n_143_99), .B (n_146_99), .C1 (n_142_99), .C2 (n_136_102) );
AOI211_X1 g_145_100 (.ZN (n_145_100), .A (n_144_101), .B (n_144_100), .C1 (n_144_98), .C2 (n_138_101) );
AOI211_X1 g_147_101 (.ZN (n_147_101), .A (n_146_102), .B (n_142_101), .C1 (n_146_99), .C2 (n_140_100) );
AOI211_X1 g_148_103 (.ZN (n_148_103), .A (n_145_100), .B (n_143_99), .C1 (n_144_100), .C2 (n_142_99) );
AOI211_X1 g_146_104 (.ZN (n_146_104), .A (n_147_101), .B (n_144_101), .C1 (n_142_101), .C2 (n_144_98) );
AOI211_X1 g_145_102 (.ZN (n_145_102), .A (n_148_103), .B (n_146_102), .C1 (n_143_99), .C2 (n_146_99) );
AOI211_X1 g_143_101 (.ZN (n_143_101), .A (n_146_104), .B (n_145_100), .C1 (n_144_101), .C2 (n_144_100) );
AOI211_X1 g_141_100 (.ZN (n_141_100), .A (n_145_102), .B (n_147_101), .C1 (n_146_102), .C2 (n_142_101) );
AOI211_X1 g_139_101 (.ZN (n_139_101), .A (n_143_101), .B (n_148_103), .C1 (n_145_100), .C2 (n_143_99) );
AOI211_X1 g_137_102 (.ZN (n_137_102), .A (n_141_100), .B (n_146_104), .C1 (n_147_101), .C2 (n_144_101) );
AOI211_X1 g_135_103 (.ZN (n_135_103), .A (n_139_101), .B (n_145_102), .C1 (n_148_103), .C2 (n_146_102) );
AOI211_X1 g_133_104 (.ZN (n_133_104), .A (n_137_102), .B (n_143_101), .C1 (n_146_104), .C2 (n_145_100) );
AOI211_X1 g_131_105 (.ZN (n_131_105), .A (n_135_103), .B (n_141_100), .C1 (n_145_102), .C2 (n_147_101) );
AOI211_X1 g_129_106 (.ZN (n_129_106), .A (n_133_104), .B (n_139_101), .C1 (n_143_101), .C2 (n_148_103) );
AOI211_X1 g_127_107 (.ZN (n_127_107), .A (n_131_105), .B (n_137_102), .C1 (n_141_100), .C2 (n_146_104) );
AOI211_X1 g_125_108 (.ZN (n_125_108), .A (n_129_106), .B (n_135_103), .C1 (n_139_101), .C2 (n_145_102) );
AOI211_X1 g_123_109 (.ZN (n_123_109), .A (n_127_107), .B (n_133_104), .C1 (n_137_102), .C2 (n_143_101) );
AOI211_X1 g_121_110 (.ZN (n_121_110), .A (n_125_108), .B (n_131_105), .C1 (n_135_103), .C2 (n_141_100) );
AOI211_X1 g_119_111 (.ZN (n_119_111), .A (n_123_109), .B (n_129_106), .C1 (n_133_104), .C2 (n_139_101) );
AOI211_X1 g_117_112 (.ZN (n_117_112), .A (n_121_110), .B (n_127_107), .C1 (n_131_105), .C2 (n_137_102) );
AOI211_X1 g_115_113 (.ZN (n_115_113), .A (n_119_111), .B (n_125_108), .C1 (n_129_106), .C2 (n_135_103) );
AOI211_X1 g_113_114 (.ZN (n_113_114), .A (n_117_112), .B (n_123_109), .C1 (n_127_107), .C2 (n_133_104) );
AOI211_X1 g_111_115 (.ZN (n_111_115), .A (n_115_113), .B (n_121_110), .C1 (n_125_108), .C2 (n_131_105) );
AOI211_X1 g_109_116 (.ZN (n_109_116), .A (n_113_114), .B (n_119_111), .C1 (n_123_109), .C2 (n_129_106) );
AOI211_X1 g_107_117 (.ZN (n_107_117), .A (n_111_115), .B (n_117_112), .C1 (n_121_110), .C2 (n_127_107) );
AOI211_X1 g_105_116 (.ZN (n_105_116), .A (n_109_116), .B (n_115_113), .C1 (n_119_111), .C2 (n_125_108) );
AOI211_X1 g_103_117 (.ZN (n_103_117), .A (n_107_117), .B (n_113_114), .C1 (n_117_112), .C2 (n_123_109) );
AOI211_X1 g_101_118 (.ZN (n_101_118), .A (n_105_116), .B (n_111_115), .C1 (n_115_113), .C2 (n_121_110) );
AOI211_X1 g_99_119 (.ZN (n_99_119), .A (n_103_117), .B (n_109_116), .C1 (n_113_114), .C2 (n_119_111) );
AOI211_X1 g_97_120 (.ZN (n_97_120), .A (n_101_118), .B (n_107_117), .C1 (n_111_115), .C2 (n_117_112) );
AOI211_X1 g_95_121 (.ZN (n_95_121), .A (n_99_119), .B (n_105_116), .C1 (n_109_116), .C2 (n_115_113) );
AOI211_X1 g_93_122 (.ZN (n_93_122), .A (n_97_120), .B (n_103_117), .C1 (n_107_117), .C2 (n_113_114) );
AOI211_X1 g_91_123 (.ZN (n_91_123), .A (n_95_121), .B (n_101_118), .C1 (n_105_116), .C2 (n_111_115) );
AOI211_X1 g_89_124 (.ZN (n_89_124), .A (n_93_122), .B (n_99_119), .C1 (n_103_117), .C2 (n_109_116) );
AOI211_X1 g_88_126 (.ZN (n_88_126), .A (n_91_123), .B (n_97_120), .C1 (n_101_118), .C2 (n_107_117) );
AOI211_X1 g_90_125 (.ZN (n_90_125), .A (n_89_124), .B (n_95_121), .C1 (n_99_119), .C2 (n_105_116) );
AOI211_X1 g_92_124 (.ZN (n_92_124), .A (n_88_126), .B (n_93_122), .C1 (n_97_120), .C2 (n_103_117) );
AOI211_X1 g_94_123 (.ZN (n_94_123), .A (n_90_125), .B (n_91_123), .C1 (n_95_121), .C2 (n_101_118) );
AOI211_X1 g_96_122 (.ZN (n_96_122), .A (n_92_124), .B (n_89_124), .C1 (n_93_122), .C2 (n_99_119) );
AOI211_X1 g_98_121 (.ZN (n_98_121), .A (n_94_123), .B (n_88_126), .C1 (n_91_123), .C2 (n_97_120) );
AOI211_X1 g_100_120 (.ZN (n_100_120), .A (n_96_122), .B (n_90_125), .C1 (n_89_124), .C2 (n_95_121) );
AOI211_X1 g_102_119 (.ZN (n_102_119), .A (n_98_121), .B (n_92_124), .C1 (n_88_126), .C2 (n_93_122) );
AOI211_X1 g_104_118 (.ZN (n_104_118), .A (n_100_120), .B (n_94_123), .C1 (n_90_125), .C2 (n_91_123) );
AOI211_X1 g_106_117 (.ZN (n_106_117), .A (n_102_119), .B (n_96_122), .C1 (n_92_124), .C2 (n_89_124) );
AOI211_X1 g_108_116 (.ZN (n_108_116), .A (n_104_118), .B (n_98_121), .C1 (n_94_123), .C2 (n_88_126) );
AOI211_X1 g_110_115 (.ZN (n_110_115), .A (n_106_117), .B (n_100_120), .C1 (n_96_122), .C2 (n_90_125) );
AOI211_X1 g_112_114 (.ZN (n_112_114), .A (n_108_116), .B (n_102_119), .C1 (n_98_121), .C2 (n_92_124) );
AOI211_X1 g_111_116 (.ZN (n_111_116), .A (n_110_115), .B (n_104_118), .C1 (n_100_120), .C2 (n_94_123) );
AOI211_X1 g_113_115 (.ZN (n_113_115), .A (n_112_114), .B (n_106_117), .C1 (n_102_119), .C2 (n_96_122) );
AOI211_X1 g_115_114 (.ZN (n_115_114), .A (n_111_116), .B (n_108_116), .C1 (n_104_118), .C2 (n_98_121) );
AOI211_X1 g_113_113 (.ZN (n_113_113), .A (n_113_115), .B (n_110_115), .C1 (n_106_117), .C2 (n_100_120) );
AOI211_X1 g_115_112 (.ZN (n_115_112), .A (n_115_114), .B (n_112_114), .C1 (n_108_116), .C2 (n_102_119) );
AOI211_X1 g_117_111 (.ZN (n_117_111), .A (n_113_113), .B (n_111_116), .C1 (n_110_115), .C2 (n_104_118) );
AOI211_X1 g_119_110 (.ZN (n_119_110), .A (n_115_112), .B (n_113_115), .C1 (n_112_114), .C2 (n_106_117) );
AOI211_X1 g_121_109 (.ZN (n_121_109), .A (n_117_111), .B (n_115_114), .C1 (n_111_116), .C2 (n_108_116) );
AOI211_X1 g_123_108 (.ZN (n_123_108), .A (n_119_110), .B (n_113_113), .C1 (n_113_115), .C2 (n_110_115) );
AOI211_X1 g_125_107 (.ZN (n_125_107), .A (n_121_109), .B (n_115_112), .C1 (n_115_114), .C2 (n_112_114) );
AOI211_X1 g_127_106 (.ZN (n_127_106), .A (n_123_108), .B (n_117_111), .C1 (n_113_113), .C2 (n_111_116) );
AOI211_X1 g_126_108 (.ZN (n_126_108), .A (n_125_107), .B (n_119_110), .C1 (n_115_112), .C2 (n_113_115) );
AOI211_X1 g_128_107 (.ZN (n_128_107), .A (n_127_106), .B (n_121_109), .C1 (n_117_111), .C2 (n_115_114) );
AOI211_X1 g_127_109 (.ZN (n_127_109), .A (n_126_108), .B (n_123_108), .C1 (n_119_110), .C2 (n_113_113) );
AOI211_X1 g_129_108 (.ZN (n_129_108), .A (n_128_107), .B (n_125_107), .C1 (n_121_109), .C2 (n_115_112) );
AOI211_X1 g_131_107 (.ZN (n_131_107), .A (n_127_109), .B (n_127_106), .C1 (n_123_108), .C2 (n_117_111) );
AOI211_X1 g_133_106 (.ZN (n_133_106), .A (n_129_108), .B (n_126_108), .C1 (n_125_107), .C2 (n_119_110) );
AOI211_X1 g_135_105 (.ZN (n_135_105), .A (n_131_107), .B (n_128_107), .C1 (n_127_106), .C2 (n_121_109) );
AOI211_X1 g_137_104 (.ZN (n_137_104), .A (n_133_106), .B (n_127_109), .C1 (n_126_108), .C2 (n_123_108) );
AOI211_X1 g_139_103 (.ZN (n_139_103), .A (n_135_105), .B (n_129_108), .C1 (n_128_107), .C2 (n_125_107) );
AOI211_X1 g_141_102 (.ZN (n_141_102), .A (n_137_104), .B (n_131_107), .C1 (n_127_109), .C2 (n_127_106) );
AOI211_X1 g_143_103 (.ZN (n_143_103), .A (n_139_103), .B (n_133_106), .C1 (n_129_108), .C2 (n_126_108) );
AOI211_X1 g_144_105 (.ZN (n_144_105), .A (n_141_102), .B (n_135_105), .C1 (n_131_107), .C2 (n_128_107) );
AOI211_X1 g_146_106 (.ZN (n_146_106), .A (n_143_103), .B (n_137_104), .C1 (n_133_106), .C2 (n_127_109) );
AOI211_X1 g_148_107 (.ZN (n_148_107), .A (n_144_105), .B (n_139_103), .C1 (n_135_105), .C2 (n_129_108) );
AOI211_X1 g_147_105 (.ZN (n_147_105), .A (n_146_106), .B (n_141_102), .C1 (n_137_104), .C2 (n_131_107) );
AOI211_X1 g_145_104 (.ZN (n_145_104), .A (n_148_107), .B (n_143_103), .C1 (n_139_103), .C2 (n_133_106) );
AOI211_X1 g_144_102 (.ZN (n_144_102), .A (n_147_105), .B (n_144_105), .C1 (n_141_102), .C2 (n_135_105) );
AOI211_X1 g_143_100 (.ZN (n_143_100), .A (n_145_104), .B (n_146_106), .C1 (n_143_103), .C2 (n_137_104) );
AOI211_X1 g_145_101 (.ZN (n_145_101), .A (n_144_102), .B (n_148_107), .C1 (n_144_105), .C2 (n_139_103) );
AOI211_X1 g_146_103 (.ZN (n_146_103), .A (n_143_100), .B (n_147_105), .C1 (n_146_106), .C2 (n_141_102) );
AOI211_X1 g_144_104 (.ZN (n_144_104), .A (n_145_101), .B (n_145_104), .C1 (n_148_107), .C2 (n_143_103) );
AOI211_X1 g_143_102 (.ZN (n_143_102), .A (n_146_103), .B (n_144_102), .C1 (n_147_105), .C2 (n_144_105) );
AOI211_X1 g_141_101 (.ZN (n_141_101), .A (n_144_104), .B (n_143_100), .C1 (n_145_104), .C2 (n_146_106) );
AOI211_X1 g_139_102 (.ZN (n_139_102), .A (n_143_102), .B (n_145_101), .C1 (n_144_102), .C2 (n_148_107) );
AOI211_X1 g_137_103 (.ZN (n_137_103), .A (n_141_101), .B (n_146_103), .C1 (n_143_100), .C2 (n_147_105) );
AOI211_X1 g_135_104 (.ZN (n_135_104), .A (n_139_102), .B (n_144_104), .C1 (n_145_101), .C2 (n_145_104) );
AOI211_X1 g_133_105 (.ZN (n_133_105), .A (n_137_103), .B (n_143_102), .C1 (n_146_103), .C2 (n_144_102) );
AOI211_X1 g_131_106 (.ZN (n_131_106), .A (n_135_104), .B (n_141_101), .C1 (n_144_104), .C2 (n_143_100) );
AOI211_X1 g_129_107 (.ZN (n_129_107), .A (n_133_105), .B (n_139_102), .C1 (n_143_102), .C2 (n_145_101) );
AOI211_X1 g_127_108 (.ZN (n_127_108), .A (n_131_106), .B (n_137_103), .C1 (n_141_101), .C2 (n_146_103) );
AOI211_X1 g_125_109 (.ZN (n_125_109), .A (n_129_107), .B (n_135_104), .C1 (n_139_102), .C2 (n_144_104) );
AOI211_X1 g_123_110 (.ZN (n_123_110), .A (n_127_108), .B (n_133_105), .C1 (n_137_103), .C2 (n_143_102) );
AOI211_X1 g_121_111 (.ZN (n_121_111), .A (n_125_109), .B (n_131_106), .C1 (n_135_104), .C2 (n_141_101) );
AOI211_X1 g_119_112 (.ZN (n_119_112), .A (n_123_110), .B (n_129_107), .C1 (n_133_105), .C2 (n_139_102) );
AOI211_X1 g_117_113 (.ZN (n_117_113), .A (n_121_111), .B (n_127_108), .C1 (n_131_106), .C2 (n_137_103) );
AOI211_X1 g_116_115 (.ZN (n_116_115), .A (n_119_112), .B (n_125_109), .C1 (n_129_107), .C2 (n_135_104) );
AOI211_X1 g_114_114 (.ZN (n_114_114), .A (n_117_113), .B (n_123_110), .C1 (n_127_108), .C2 (n_133_105) );
AOI211_X1 g_116_113 (.ZN (n_116_113), .A (n_116_115), .B (n_121_111), .C1 (n_125_109), .C2 (n_131_106) );
AOI211_X1 g_118_112 (.ZN (n_118_112), .A (n_114_114), .B (n_119_112), .C1 (n_123_110), .C2 (n_129_107) );
AOI211_X1 g_120_111 (.ZN (n_120_111), .A (n_116_113), .B (n_117_113), .C1 (n_121_111), .C2 (n_127_108) );
AOI211_X1 g_122_110 (.ZN (n_122_110), .A (n_118_112), .B (n_116_115), .C1 (n_119_112), .C2 (n_125_109) );
AOI211_X1 g_124_109 (.ZN (n_124_109), .A (n_120_111), .B (n_114_114), .C1 (n_117_113), .C2 (n_123_110) );
AOI211_X1 g_123_111 (.ZN (n_123_111), .A (n_122_110), .B (n_116_113), .C1 (n_116_115), .C2 (n_121_111) );
AOI211_X1 g_125_110 (.ZN (n_125_110), .A (n_124_109), .B (n_118_112), .C1 (n_114_114), .C2 (n_119_112) );
AOI211_X1 g_124_112 (.ZN (n_124_112), .A (n_123_111), .B (n_120_111), .C1 (n_116_113), .C2 (n_117_113) );
AOI211_X1 g_122_111 (.ZN (n_122_111), .A (n_125_110), .B (n_122_110), .C1 (n_118_112), .C2 (n_116_115) );
AOI211_X1 g_124_110 (.ZN (n_124_110), .A (n_124_112), .B (n_124_109), .C1 (n_120_111), .C2 (n_114_114) );
AOI211_X1 g_126_109 (.ZN (n_126_109), .A (n_122_111), .B (n_123_111), .C1 (n_122_110), .C2 (n_116_113) );
AOI211_X1 g_128_108 (.ZN (n_128_108), .A (n_124_110), .B (n_125_110), .C1 (n_124_109), .C2 (n_118_112) );
AOI211_X1 g_130_107 (.ZN (n_130_107), .A (n_126_109), .B (n_124_112), .C1 (n_123_111), .C2 (n_120_111) );
AOI211_X1 g_132_106 (.ZN (n_132_106), .A (n_128_108), .B (n_122_111), .C1 (n_125_110), .C2 (n_122_110) );
AOI211_X1 g_134_105 (.ZN (n_134_105), .A (n_130_107), .B (n_124_110), .C1 (n_124_112), .C2 (n_124_109) );
AOI211_X1 g_136_104 (.ZN (n_136_104), .A (n_132_106), .B (n_126_109), .C1 (n_122_111), .C2 (n_123_111) );
AOI211_X1 g_138_103 (.ZN (n_138_103), .A (n_134_105), .B (n_128_108), .C1 (n_124_110), .C2 (n_125_110) );
AOI211_X1 g_140_102 (.ZN (n_140_102), .A (n_136_104), .B (n_130_107), .C1 (n_126_109), .C2 (n_124_112) );
AOI211_X1 g_142_103 (.ZN (n_142_103), .A (n_138_103), .B (n_132_106), .C1 (n_128_108), .C2 (n_122_111) );
AOI211_X1 g_140_104 (.ZN (n_140_104), .A (n_140_102), .B (n_134_105), .C1 (n_130_107), .C2 (n_124_110) );
AOI211_X1 g_138_105 (.ZN (n_138_105), .A (n_142_103), .B (n_136_104), .C1 (n_132_106), .C2 (n_126_109) );
AOI211_X1 g_136_106 (.ZN (n_136_106), .A (n_140_104), .B (n_138_103), .C1 (n_134_105), .C2 (n_128_108) );
AOI211_X1 g_134_107 (.ZN (n_134_107), .A (n_138_105), .B (n_140_102), .C1 (n_136_104), .C2 (n_130_107) );
AOI211_X1 g_132_108 (.ZN (n_132_108), .A (n_136_106), .B (n_142_103), .C1 (n_138_103), .C2 (n_132_106) );
AOI211_X1 g_130_109 (.ZN (n_130_109), .A (n_134_107), .B (n_140_104), .C1 (n_140_102), .C2 (n_134_105) );
AOI211_X1 g_128_110 (.ZN (n_128_110), .A (n_132_108), .B (n_138_105), .C1 (n_142_103), .C2 (n_136_104) );
AOI211_X1 g_126_111 (.ZN (n_126_111), .A (n_130_109), .B (n_136_106), .C1 (n_140_104), .C2 (n_138_103) );
AOI211_X1 g_125_113 (.ZN (n_125_113), .A (n_128_110), .B (n_134_107), .C1 (n_138_105), .C2 (n_140_102) );
AOI211_X1 g_124_111 (.ZN (n_124_111), .A (n_126_111), .B (n_132_108), .C1 (n_136_106), .C2 (n_142_103) );
AOI211_X1 g_126_110 (.ZN (n_126_110), .A (n_125_113), .B (n_130_109), .C1 (n_134_107), .C2 (n_140_104) );
AOI211_X1 g_128_109 (.ZN (n_128_109), .A (n_124_111), .B (n_128_110), .C1 (n_132_108), .C2 (n_138_105) );
AOI211_X1 g_130_108 (.ZN (n_130_108), .A (n_126_110), .B (n_126_111), .C1 (n_130_109), .C2 (n_136_106) );
AOI211_X1 g_132_107 (.ZN (n_132_107), .A (n_128_109), .B (n_125_113), .C1 (n_128_110), .C2 (n_134_107) );
AOI211_X1 g_134_106 (.ZN (n_134_106), .A (n_130_108), .B (n_124_111), .C1 (n_126_111), .C2 (n_132_108) );
AOI211_X1 g_136_105 (.ZN (n_136_105), .A (n_132_107), .B (n_126_110), .C1 (n_125_113), .C2 (n_130_109) );
AOI211_X1 g_138_104 (.ZN (n_138_104), .A (n_134_106), .B (n_128_109), .C1 (n_124_111), .C2 (n_128_110) );
AOI211_X1 g_140_103 (.ZN (n_140_103), .A (n_136_105), .B (n_130_108), .C1 (n_126_110), .C2 (n_126_111) );
AOI211_X1 g_142_102 (.ZN (n_142_102), .A (n_138_104), .B (n_132_107), .C1 (n_128_109), .C2 (n_125_113) );
AOI211_X1 g_144_103 (.ZN (n_144_103), .A (n_140_103), .B (n_134_106), .C1 (n_130_108), .C2 (n_124_111) );
AOI211_X1 g_142_104 (.ZN (n_142_104), .A (n_142_102), .B (n_136_105), .C1 (n_132_107), .C2 (n_126_110) );
AOI211_X1 g_140_105 (.ZN (n_140_105), .A (n_144_103), .B (n_138_104), .C1 (n_134_106), .C2 (n_128_109) );
AOI211_X1 g_141_103 (.ZN (n_141_103), .A (n_142_104), .B (n_140_103), .C1 (n_136_105), .C2 (n_130_108) );
AOI211_X1 g_139_104 (.ZN (n_139_104), .A (n_140_105), .B (n_142_102), .C1 (n_138_104), .C2 (n_132_107) );
AOI211_X1 g_137_105 (.ZN (n_137_105), .A (n_141_103), .B (n_144_103), .C1 (n_140_103), .C2 (n_134_106) );
AOI211_X1 g_135_106 (.ZN (n_135_106), .A (n_139_104), .B (n_142_104), .C1 (n_142_102), .C2 (n_136_105) );
AOI211_X1 g_133_107 (.ZN (n_133_107), .A (n_137_105), .B (n_140_105), .C1 (n_144_103), .C2 (n_138_104) );
AOI211_X1 g_131_108 (.ZN (n_131_108), .A (n_135_106), .B (n_141_103), .C1 (n_142_104), .C2 (n_140_103) );
AOI211_X1 g_129_109 (.ZN (n_129_109), .A (n_133_107), .B (n_139_104), .C1 (n_140_105), .C2 (n_142_102) );
AOI211_X1 g_127_110 (.ZN (n_127_110), .A (n_131_108), .B (n_137_105), .C1 (n_141_103), .C2 (n_144_103) );
AOI211_X1 g_125_111 (.ZN (n_125_111), .A (n_129_109), .B (n_135_106), .C1 (n_139_104), .C2 (n_142_104) );
AOI211_X1 g_123_112 (.ZN (n_123_112), .A (n_127_110), .B (n_133_107), .C1 (n_137_105), .C2 (n_140_105) );
AOI211_X1 g_121_113 (.ZN (n_121_113), .A (n_125_111), .B (n_131_108), .C1 (n_135_106), .C2 (n_141_103) );
AOI211_X1 g_119_114 (.ZN (n_119_114), .A (n_123_112), .B (n_129_109), .C1 (n_133_107), .C2 (n_139_104) );
AOI211_X1 g_120_112 (.ZN (n_120_112), .A (n_121_113), .B (n_127_110), .C1 (n_131_108), .C2 (n_137_105) );
AOI211_X1 g_118_113 (.ZN (n_118_113), .A (n_119_114), .B (n_125_111), .C1 (n_129_109), .C2 (n_135_106) );
AOI211_X1 g_116_114 (.ZN (n_116_114), .A (n_120_112), .B (n_123_112), .C1 (n_127_110), .C2 (n_133_107) );
AOI211_X1 g_114_115 (.ZN (n_114_115), .A (n_118_113), .B (n_121_113), .C1 (n_125_111), .C2 (n_131_108) );
AOI211_X1 g_112_116 (.ZN (n_112_116), .A (n_116_114), .B (n_119_114), .C1 (n_123_112), .C2 (n_129_109) );
AOI211_X1 g_110_117 (.ZN (n_110_117), .A (n_114_115), .B (n_120_112), .C1 (n_121_113), .C2 (n_127_110) );
AOI211_X1 g_108_118 (.ZN (n_108_118), .A (n_112_116), .B (n_118_113), .C1 (n_119_114), .C2 (n_125_111) );
AOI211_X1 g_106_119 (.ZN (n_106_119), .A (n_110_117), .B (n_116_114), .C1 (n_120_112), .C2 (n_123_112) );
AOI211_X1 g_104_120 (.ZN (n_104_120), .A (n_108_118), .B (n_114_115), .C1 (n_118_113), .C2 (n_121_113) );
AOI211_X1 g_105_118 (.ZN (n_105_118), .A (n_106_119), .B (n_112_116), .C1 (n_116_114), .C2 (n_119_114) );
AOI211_X1 g_103_119 (.ZN (n_103_119), .A (n_104_120), .B (n_110_117), .C1 (n_114_115), .C2 (n_120_112) );
AOI211_X1 g_101_120 (.ZN (n_101_120), .A (n_105_118), .B (n_108_118), .C1 (n_112_116), .C2 (n_118_113) );
AOI211_X1 g_99_121 (.ZN (n_99_121), .A (n_103_119), .B (n_106_119), .C1 (n_110_117), .C2 (n_116_114) );
AOI211_X1 g_97_122 (.ZN (n_97_122), .A (n_101_120), .B (n_104_120), .C1 (n_108_118), .C2 (n_114_115) );
AOI211_X1 g_95_123 (.ZN (n_95_123), .A (n_99_121), .B (n_105_118), .C1 (n_106_119), .C2 (n_112_116) );
AOI211_X1 g_93_124 (.ZN (n_93_124), .A (n_97_122), .B (n_103_119), .C1 (n_104_120), .C2 (n_110_117) );
AOI211_X1 g_91_125 (.ZN (n_91_125), .A (n_95_123), .B (n_101_120), .C1 (n_105_118), .C2 (n_108_118) );
AOI211_X1 g_89_126 (.ZN (n_89_126), .A (n_93_124), .B (n_99_121), .C1 (n_103_119), .C2 (n_106_119) );
AOI211_X1 g_87_127 (.ZN (n_87_127), .A (n_91_125), .B (n_97_122), .C1 (n_101_120), .C2 (n_104_120) );
AOI211_X1 g_85_126 (.ZN (n_85_126), .A (n_89_126), .B (n_95_123), .C1 (n_99_121), .C2 (n_105_118) );
AOI211_X1 g_83_127 (.ZN (n_83_127), .A (n_87_127), .B (n_93_124), .C1 (n_97_122), .C2 (n_103_119) );
AOI211_X1 g_81_128 (.ZN (n_81_128), .A (n_85_126), .B (n_91_125), .C1 (n_95_123), .C2 (n_101_120) );
AOI211_X1 g_79_129 (.ZN (n_79_129), .A (n_83_127), .B (n_89_126), .C1 (n_93_124), .C2 (n_99_121) );
AOI211_X1 g_77_130 (.ZN (n_77_130), .A (n_81_128), .B (n_87_127), .C1 (n_91_125), .C2 (n_97_122) );
AOI211_X1 g_76_132 (.ZN (n_76_132), .A (n_79_129), .B (n_85_126), .C1 (n_89_126), .C2 (n_95_123) );
AOI211_X1 g_78_131 (.ZN (n_78_131), .A (n_77_130), .B (n_83_127), .C1 (n_87_127), .C2 (n_93_124) );
AOI211_X1 g_80_130 (.ZN (n_80_130), .A (n_76_132), .B (n_81_128), .C1 (n_85_126), .C2 (n_91_125) );
AOI211_X1 g_82_129 (.ZN (n_82_129), .A (n_78_131), .B (n_79_129), .C1 (n_83_127), .C2 (n_89_126) );
AOI211_X1 g_84_128 (.ZN (n_84_128), .A (n_80_130), .B (n_77_130), .C1 (n_81_128), .C2 (n_87_127) );
AOI211_X1 g_86_129 (.ZN (n_86_129), .A (n_82_129), .B (n_76_132), .C1 (n_79_129), .C2 (n_85_126) );
AOI211_X1 g_88_128 (.ZN (n_88_128), .A (n_84_128), .B (n_78_131), .C1 (n_77_130), .C2 (n_83_127) );
AOI211_X1 g_90_127 (.ZN (n_90_127), .A (n_86_129), .B (n_80_130), .C1 (n_76_132), .C2 (n_81_128) );
AOI211_X1 g_92_126 (.ZN (n_92_126), .A (n_88_128), .B (n_82_129), .C1 (n_78_131), .C2 (n_79_129) );
AOI211_X1 g_94_125 (.ZN (n_94_125), .A (n_90_127), .B (n_84_128), .C1 (n_80_130), .C2 (n_77_130) );
AOI211_X1 g_96_124 (.ZN (n_96_124), .A (n_92_126), .B (n_86_129), .C1 (n_82_129), .C2 (n_76_132) );
AOI211_X1 g_98_123 (.ZN (n_98_123), .A (n_94_125), .B (n_88_128), .C1 (n_84_128), .C2 (n_78_131) );
AOI211_X1 g_100_122 (.ZN (n_100_122), .A (n_96_124), .B (n_90_127), .C1 (n_86_129), .C2 (n_80_130) );
AOI211_X1 g_102_121 (.ZN (n_102_121), .A (n_98_123), .B (n_92_126), .C1 (n_88_128), .C2 (n_82_129) );
AOI211_X1 g_101_123 (.ZN (n_101_123), .A (n_100_122), .B (n_94_125), .C1 (n_90_127), .C2 (n_84_128) );
AOI211_X1 g_100_121 (.ZN (n_100_121), .A (n_102_121), .B (n_96_124), .C1 (n_92_126), .C2 (n_86_129) );
AOI211_X1 g_102_120 (.ZN (n_102_120), .A (n_101_123), .B (n_98_123), .C1 (n_94_125), .C2 (n_88_128) );
AOI211_X1 g_104_119 (.ZN (n_104_119), .A (n_100_121), .B (n_100_122), .C1 (n_96_124), .C2 (n_90_127) );
AOI211_X1 g_106_118 (.ZN (n_106_118), .A (n_102_120), .B (n_102_121), .C1 (n_98_123), .C2 (n_92_126) );
AOI211_X1 g_105_120 (.ZN (n_105_120), .A (n_104_119), .B (n_101_123), .C1 (n_100_122), .C2 (n_94_125) );
AOI211_X1 g_107_119 (.ZN (n_107_119), .A (n_106_118), .B (n_100_121), .C1 (n_102_121), .C2 (n_96_124) );
AOI211_X1 g_109_118 (.ZN (n_109_118), .A (n_105_120), .B (n_102_120), .C1 (n_101_123), .C2 (n_98_123) );
AOI211_X1 g_110_116 (.ZN (n_110_116), .A (n_107_119), .B (n_104_119), .C1 (n_100_121), .C2 (n_100_122) );
AOI211_X1 g_112_115 (.ZN (n_112_115), .A (n_109_118), .B (n_106_118), .C1 (n_102_120), .C2 (n_102_121) );
AOI211_X1 g_111_117 (.ZN (n_111_117), .A (n_110_116), .B (n_105_120), .C1 (n_104_119), .C2 (n_101_123) );
AOI211_X1 g_113_116 (.ZN (n_113_116), .A (n_112_115), .B (n_107_119), .C1 (n_106_118), .C2 (n_100_121) );
AOI211_X1 g_115_115 (.ZN (n_115_115), .A (n_111_117), .B (n_109_118), .C1 (n_105_120), .C2 (n_102_120) );
AOI211_X1 g_117_114 (.ZN (n_117_114), .A (n_113_116), .B (n_110_116), .C1 (n_107_119), .C2 (n_104_119) );
AOI211_X1 g_119_113 (.ZN (n_119_113), .A (n_115_115), .B (n_112_115), .C1 (n_109_118), .C2 (n_106_118) );
AOI211_X1 g_121_112 (.ZN (n_121_112), .A (n_117_114), .B (n_111_117), .C1 (n_110_116), .C2 (n_105_120) );
AOI211_X1 g_120_114 (.ZN (n_120_114), .A (n_119_113), .B (n_113_116), .C1 (n_112_115), .C2 (n_107_119) );
AOI211_X1 g_122_113 (.ZN (n_122_113), .A (n_121_112), .B (n_115_115), .C1 (n_111_117), .C2 (n_109_118) );
AOI211_X1 g_121_115 (.ZN (n_121_115), .A (n_120_114), .B (n_117_114), .C1 (n_113_116), .C2 (n_110_116) );
AOI211_X1 g_123_114 (.ZN (n_123_114), .A (n_122_113), .B (n_119_113), .C1 (n_115_115), .C2 (n_112_115) );
AOI211_X1 g_122_112 (.ZN (n_122_112), .A (n_121_115), .B (n_121_112), .C1 (n_117_114), .C2 (n_111_117) );
AOI211_X1 g_120_113 (.ZN (n_120_113), .A (n_123_114), .B (n_120_114), .C1 (n_119_113), .C2 (n_113_116) );
AOI211_X1 g_118_114 (.ZN (n_118_114), .A (n_122_112), .B (n_122_113), .C1 (n_121_112), .C2 (n_115_115) );
AOI211_X1 g_117_116 (.ZN (n_117_116), .A (n_120_113), .B (n_121_115), .C1 (n_120_114), .C2 (n_117_114) );
AOI211_X1 g_119_115 (.ZN (n_119_115), .A (n_118_114), .B (n_123_114), .C1 (n_122_113), .C2 (n_119_113) );
AOI211_X1 g_121_114 (.ZN (n_121_114), .A (n_117_116), .B (n_122_112), .C1 (n_121_115), .C2 (n_121_112) );
AOI211_X1 g_123_113 (.ZN (n_123_113), .A (n_119_115), .B (n_120_113), .C1 (n_123_114), .C2 (n_120_114) );
AOI211_X1 g_125_112 (.ZN (n_125_112), .A (n_121_114), .B (n_118_114), .C1 (n_122_112), .C2 (n_122_113) );
AOI211_X1 g_127_111 (.ZN (n_127_111), .A (n_123_113), .B (n_117_116), .C1 (n_120_113), .C2 (n_121_115) );
AOI211_X1 g_129_110 (.ZN (n_129_110), .A (n_125_112), .B (n_119_115), .C1 (n_118_114), .C2 (n_123_114) );
AOI211_X1 g_131_109 (.ZN (n_131_109), .A (n_127_111), .B (n_121_114), .C1 (n_117_116), .C2 (n_122_112) );
AOI211_X1 g_133_108 (.ZN (n_133_108), .A (n_129_110), .B (n_123_113), .C1 (n_119_115), .C2 (n_120_113) );
AOI211_X1 g_135_107 (.ZN (n_135_107), .A (n_131_109), .B (n_125_112), .C1 (n_121_114), .C2 (n_118_114) );
AOI211_X1 g_137_106 (.ZN (n_137_106), .A (n_133_108), .B (n_127_111), .C1 (n_123_113), .C2 (n_117_116) );
AOI211_X1 g_139_105 (.ZN (n_139_105), .A (n_135_107), .B (n_129_110), .C1 (n_125_112), .C2 (n_119_115) );
AOI211_X1 g_141_104 (.ZN (n_141_104), .A (n_137_106), .B (n_131_109), .C1 (n_127_111), .C2 (n_121_114) );
AOI211_X1 g_143_105 (.ZN (n_143_105), .A (n_139_105), .B (n_133_108), .C1 (n_129_110), .C2 (n_123_113) );
AOI211_X1 g_145_106 (.ZN (n_145_106), .A (n_141_104), .B (n_135_107), .C1 (n_131_109), .C2 (n_125_112) );
AOI211_X1 g_146_108 (.ZN (n_146_108), .A (n_143_105), .B (n_137_106), .C1 (n_133_108), .C2 (n_127_111) );
AOI211_X1 g_144_107 (.ZN (n_144_107), .A (n_145_106), .B (n_139_105), .C1 (n_135_107), .C2 (n_129_110) );
AOI211_X1 g_145_105 (.ZN (n_145_105), .A (n_146_108), .B (n_141_104), .C1 (n_137_106), .C2 (n_131_109) );
AOI211_X1 g_143_104 (.ZN (n_143_104), .A (n_144_107), .B (n_143_105), .C1 (n_139_105), .C2 (n_133_108) );
AOI211_X1 g_142_106 (.ZN (n_142_106), .A (n_145_105), .B (n_145_106), .C1 (n_141_104), .C2 (n_135_107) );
AOI211_X1 g_140_107 (.ZN (n_140_107), .A (n_143_104), .B (n_146_108), .C1 (n_143_105), .C2 (n_137_106) );
AOI211_X1 g_141_105 (.ZN (n_141_105), .A (n_142_106), .B (n_144_107), .C1 (n_145_106), .C2 (n_139_105) );
AOI211_X1 g_143_106 (.ZN (n_143_106), .A (n_140_107), .B (n_145_105), .C1 (n_146_108), .C2 (n_141_104) );
AOI211_X1 g_142_108 (.ZN (n_142_108), .A (n_141_105), .B (n_143_104), .C1 (n_144_107), .C2 (n_143_105) );
AOI211_X1 g_141_106 (.ZN (n_141_106), .A (n_143_106), .B (n_142_106), .C1 (n_145_105), .C2 (n_145_106) );
AOI211_X1 g_139_107 (.ZN (n_139_107), .A (n_142_108), .B (n_140_107), .C1 (n_143_104), .C2 (n_146_108) );
AOI211_X1 g_137_108 (.ZN (n_137_108), .A (n_141_106), .B (n_141_105), .C1 (n_142_106), .C2 (n_144_107) );
AOI211_X1 g_138_106 (.ZN (n_138_106), .A (n_139_107), .B (n_143_106), .C1 (n_140_107), .C2 (n_145_105) );
AOI211_X1 g_136_107 (.ZN (n_136_107), .A (n_137_108), .B (n_142_108), .C1 (n_141_105), .C2 (n_143_104) );
AOI211_X1 g_134_108 (.ZN (n_134_108), .A (n_138_106), .B (n_141_106), .C1 (n_143_106), .C2 (n_142_106) );
AOI211_X1 g_132_109 (.ZN (n_132_109), .A (n_136_107), .B (n_139_107), .C1 (n_142_108), .C2 (n_140_107) );
AOI211_X1 g_130_110 (.ZN (n_130_110), .A (n_134_108), .B (n_137_108), .C1 (n_141_106), .C2 (n_141_105) );
AOI211_X1 g_128_111 (.ZN (n_128_111), .A (n_132_109), .B (n_138_106), .C1 (n_139_107), .C2 (n_143_106) );
AOI211_X1 g_126_112 (.ZN (n_126_112), .A (n_130_110), .B (n_136_107), .C1 (n_137_108), .C2 (n_142_108) );
AOI211_X1 g_124_113 (.ZN (n_124_113), .A (n_128_111), .B (n_134_108), .C1 (n_138_106), .C2 (n_141_106) );
AOI211_X1 g_122_114 (.ZN (n_122_114), .A (n_126_112), .B (n_132_109), .C1 (n_136_107), .C2 (n_139_107) );
AOI211_X1 g_120_115 (.ZN (n_120_115), .A (n_124_113), .B (n_130_110), .C1 (n_134_108), .C2 (n_137_108) );
AOI211_X1 g_118_116 (.ZN (n_118_116), .A (n_122_114), .B (n_128_111), .C1 (n_132_109), .C2 (n_138_106) );
AOI211_X1 g_120_117 (.ZN (n_120_117), .A (n_120_115), .B (n_126_112), .C1 (n_130_110), .C2 (n_136_107) );
AOI211_X1 g_122_116 (.ZN (n_122_116), .A (n_118_116), .B (n_124_113), .C1 (n_128_111), .C2 (n_134_108) );
AOI211_X1 g_124_115 (.ZN (n_124_115), .A (n_120_117), .B (n_122_114), .C1 (n_126_112), .C2 (n_132_109) );
AOI211_X1 g_126_114 (.ZN (n_126_114), .A (n_122_116), .B (n_120_115), .C1 (n_124_113), .C2 (n_130_110) );
AOI211_X1 g_127_112 (.ZN (n_127_112), .A (n_124_115), .B (n_118_116), .C1 (n_122_114), .C2 (n_128_111) );
AOI211_X1 g_129_111 (.ZN (n_129_111), .A (n_126_114), .B (n_120_117), .C1 (n_120_115), .C2 (n_126_112) );
AOI211_X1 g_131_110 (.ZN (n_131_110), .A (n_127_112), .B (n_122_116), .C1 (n_118_116), .C2 (n_124_113) );
AOI211_X1 g_133_109 (.ZN (n_133_109), .A (n_129_111), .B (n_124_115), .C1 (n_120_117), .C2 (n_122_114) );
AOI211_X1 g_135_108 (.ZN (n_135_108), .A (n_131_110), .B (n_126_114), .C1 (n_122_116), .C2 (n_120_115) );
AOI211_X1 g_137_107 (.ZN (n_137_107), .A (n_133_109), .B (n_127_112), .C1 (n_124_115), .C2 (n_118_116) );
AOI211_X1 g_139_106 (.ZN (n_139_106), .A (n_135_108), .B (n_129_111), .C1 (n_126_114), .C2 (n_120_117) );
AOI211_X1 g_138_108 (.ZN (n_138_108), .A (n_137_107), .B (n_131_110), .C1 (n_127_112), .C2 (n_122_116) );
AOI211_X1 g_136_109 (.ZN (n_136_109), .A (n_139_106), .B (n_133_109), .C1 (n_129_111), .C2 (n_124_115) );
AOI211_X1 g_134_110 (.ZN (n_134_110), .A (n_138_108), .B (n_135_108), .C1 (n_131_110), .C2 (n_126_114) );
AOI211_X1 g_132_111 (.ZN (n_132_111), .A (n_136_109), .B (n_137_107), .C1 (n_133_109), .C2 (n_127_112) );
AOI211_X1 g_130_112 (.ZN (n_130_112), .A (n_134_110), .B (n_139_106), .C1 (n_135_108), .C2 (n_129_111) );
AOI211_X1 g_128_113 (.ZN (n_128_113), .A (n_132_111), .B (n_138_108), .C1 (n_137_107), .C2 (n_131_110) );
AOI211_X1 g_127_115 (.ZN (n_127_115), .A (n_130_112), .B (n_136_109), .C1 (n_139_106), .C2 (n_133_109) );
AOI211_X1 g_126_113 (.ZN (n_126_113), .A (n_128_113), .B (n_134_110), .C1 (n_138_108), .C2 (n_135_108) );
AOI211_X1 g_128_112 (.ZN (n_128_112), .A (n_127_115), .B (n_132_111), .C1 (n_136_109), .C2 (n_137_107) );
AOI211_X1 g_130_111 (.ZN (n_130_111), .A (n_126_113), .B (n_130_112), .C1 (n_134_110), .C2 (n_139_106) );
AOI211_X1 g_132_110 (.ZN (n_132_110), .A (n_128_112), .B (n_128_113), .C1 (n_132_111), .C2 (n_138_108) );
AOI211_X1 g_134_109 (.ZN (n_134_109), .A (n_130_111), .B (n_127_115), .C1 (n_130_112), .C2 (n_136_109) );
AOI211_X1 g_136_108 (.ZN (n_136_108), .A (n_132_110), .B (n_126_113), .C1 (n_128_113), .C2 (n_134_110) );
AOI211_X1 g_138_107 (.ZN (n_138_107), .A (n_134_109), .B (n_128_112), .C1 (n_127_115), .C2 (n_132_111) );
AOI211_X1 g_140_106 (.ZN (n_140_106), .A (n_136_108), .B (n_130_111), .C1 (n_126_113), .C2 (n_130_112) );
AOI211_X1 g_142_105 (.ZN (n_142_105), .A (n_138_107), .B (n_132_110), .C1 (n_128_112), .C2 (n_128_113) );
AOI211_X1 g_141_107 (.ZN (n_141_107), .A (n_140_106), .B (n_134_109), .C1 (n_130_111), .C2 (n_127_115) );
AOI211_X1 g_139_108 (.ZN (n_139_108), .A (n_142_105), .B (n_136_108), .C1 (n_132_110), .C2 (n_126_113) );
AOI211_X1 g_137_109 (.ZN (n_137_109), .A (n_141_107), .B (n_138_107), .C1 (n_134_109), .C2 (n_128_112) );
AOI211_X1 g_135_110 (.ZN (n_135_110), .A (n_139_108), .B (n_140_106), .C1 (n_136_108), .C2 (n_130_111) );
AOI211_X1 g_133_111 (.ZN (n_133_111), .A (n_137_109), .B (n_142_105), .C1 (n_138_107), .C2 (n_132_110) );
AOI211_X1 g_131_112 (.ZN (n_131_112), .A (n_135_110), .B (n_141_107), .C1 (n_140_106), .C2 (n_134_109) );
AOI211_X1 g_129_113 (.ZN (n_129_113), .A (n_133_111), .B (n_139_108), .C1 (n_142_105), .C2 (n_136_108) );
AOI211_X1 g_127_114 (.ZN (n_127_114), .A (n_131_112), .B (n_137_109), .C1 (n_141_107), .C2 (n_138_107) );
AOI211_X1 g_125_115 (.ZN (n_125_115), .A (n_129_113), .B (n_135_110), .C1 (n_139_108), .C2 (n_140_106) );
AOI211_X1 g_123_116 (.ZN (n_123_116), .A (n_127_114), .B (n_133_111), .C1 (n_137_109), .C2 (n_142_105) );
AOI211_X1 g_124_114 (.ZN (n_124_114), .A (n_125_115), .B (n_131_112), .C1 (n_135_110), .C2 (n_141_107) );
AOI211_X1 g_122_115 (.ZN (n_122_115), .A (n_123_116), .B (n_129_113), .C1 (n_133_111), .C2 (n_139_108) );
AOI211_X1 g_120_116 (.ZN (n_120_116), .A (n_124_114), .B (n_127_114), .C1 (n_131_112), .C2 (n_137_109) );
AOI211_X1 g_118_115 (.ZN (n_118_115), .A (n_122_115), .B (n_125_115), .C1 (n_129_113), .C2 (n_135_110) );
AOI211_X1 g_116_116 (.ZN (n_116_116), .A (n_120_116), .B (n_123_116), .C1 (n_127_114), .C2 (n_133_111) );
AOI211_X1 g_114_117 (.ZN (n_114_117), .A (n_118_115), .B (n_124_114), .C1 (n_125_115), .C2 (n_131_112) );
AOI211_X1 g_112_118 (.ZN (n_112_118), .A (n_116_116), .B (n_122_115), .C1 (n_123_116), .C2 (n_129_113) );
AOI211_X1 g_110_119 (.ZN (n_110_119), .A (n_114_117), .B (n_120_116), .C1 (n_124_114), .C2 (n_127_114) );
AOI211_X1 g_109_117 (.ZN (n_109_117), .A (n_112_118), .B (n_118_115), .C1 (n_122_115), .C2 (n_125_115) );
AOI211_X1 g_107_118 (.ZN (n_107_118), .A (n_110_119), .B (n_116_116), .C1 (n_120_116), .C2 (n_123_116) );
AOI211_X1 g_105_119 (.ZN (n_105_119), .A (n_109_117), .B (n_114_117), .C1 (n_118_115), .C2 (n_124_114) );
AOI211_X1 g_103_120 (.ZN (n_103_120), .A (n_107_118), .B (n_112_118), .C1 (n_116_116), .C2 (n_122_115) );
AOI211_X1 g_101_121 (.ZN (n_101_121), .A (n_105_119), .B (n_110_119), .C1 (n_114_117), .C2 (n_120_116) );
AOI211_X1 g_99_122 (.ZN (n_99_122), .A (n_103_120), .B (n_109_117), .C1 (n_112_118), .C2 (n_118_115) );
AOI211_X1 g_97_123 (.ZN (n_97_123), .A (n_101_121), .B (n_107_118), .C1 (n_110_119), .C2 (n_116_116) );
AOI211_X1 g_95_124 (.ZN (n_95_124), .A (n_99_122), .B (n_105_119), .C1 (n_109_117), .C2 (n_114_117) );
AOI211_X1 g_93_125 (.ZN (n_93_125), .A (n_97_123), .B (n_103_120), .C1 (n_107_118), .C2 (n_112_118) );
AOI211_X1 g_91_126 (.ZN (n_91_126), .A (n_95_124), .B (n_101_121), .C1 (n_105_119), .C2 (n_110_119) );
AOI211_X1 g_89_127 (.ZN (n_89_127), .A (n_93_125), .B (n_99_122), .C1 (n_103_120), .C2 (n_109_117) );
AOI211_X1 g_87_128 (.ZN (n_87_128), .A (n_91_126), .B (n_97_123), .C1 (n_101_121), .C2 (n_107_118) );
AOI211_X1 g_85_129 (.ZN (n_85_129), .A (n_89_127), .B (n_95_124), .C1 (n_99_122), .C2 (n_105_119) );
AOI211_X1 g_84_127 (.ZN (n_84_127), .A (n_87_128), .B (n_93_125), .C1 (n_97_123), .C2 (n_103_120) );
AOI211_X1 g_82_128 (.ZN (n_82_128), .A (n_85_129), .B (n_91_126), .C1 (n_95_124), .C2 (n_101_121) );
AOI211_X1 g_81_130 (.ZN (n_81_130), .A (n_84_127), .B (n_89_127), .C1 (n_93_125), .C2 (n_99_122) );
AOI211_X1 g_83_129 (.ZN (n_83_129), .A (n_82_128), .B (n_87_128), .C1 (n_91_126), .C2 (n_97_123) );
AOI211_X1 g_85_128 (.ZN (n_85_128), .A (n_81_130), .B (n_85_129), .C1 (n_89_127), .C2 (n_95_124) );
AOI211_X1 g_84_130 (.ZN (n_84_130), .A (n_83_129), .B (n_84_127), .C1 (n_87_128), .C2 (n_93_125) );
AOI211_X1 g_82_131 (.ZN (n_82_131), .A (n_85_128), .B (n_82_128), .C1 (n_85_129), .C2 (n_91_126) );
AOI211_X1 g_81_129 (.ZN (n_81_129), .A (n_84_130), .B (n_81_130), .C1 (n_84_127), .C2 (n_89_127) );
AOI211_X1 g_79_130 (.ZN (n_79_130), .A (n_82_131), .B (n_83_129), .C1 (n_82_128), .C2 (n_87_128) );
AOI211_X1 g_77_131 (.ZN (n_77_131), .A (n_81_129), .B (n_85_128), .C1 (n_81_130), .C2 (n_85_129) );
AOI211_X1 g_75_132 (.ZN (n_75_132), .A (n_79_130), .B (n_84_130), .C1 (n_83_129), .C2 (n_84_127) );
AOI211_X1 g_73_133 (.ZN (n_73_133), .A (n_77_131), .B (n_82_131), .C1 (n_85_128), .C2 (n_82_128) );
AOI211_X1 g_71_134 (.ZN (n_71_134), .A (n_75_132), .B (n_81_129), .C1 (n_84_130), .C2 (n_81_130) );
AOI211_X1 g_69_135 (.ZN (n_69_135), .A (n_73_133), .B (n_79_130), .C1 (n_82_131), .C2 (n_83_129) );
AOI211_X1 g_67_136 (.ZN (n_67_136), .A (n_71_134), .B (n_77_131), .C1 (n_81_129), .C2 (n_85_128) );
AOI211_X1 g_68_134 (.ZN (n_68_134), .A (n_69_135), .B (n_75_132), .C1 (n_79_130), .C2 (n_84_130) );
AOI211_X1 g_66_135 (.ZN (n_66_135), .A (n_67_136), .B (n_73_133), .C1 (n_77_131), .C2 (n_82_131) );
AOI211_X1 g_64_136 (.ZN (n_64_136), .A (n_68_134), .B (n_71_134), .C1 (n_75_132), .C2 (n_81_129) );
AOI211_X1 g_62_137 (.ZN (n_62_137), .A (n_66_135), .B (n_69_135), .C1 (n_73_133), .C2 (n_79_130) );
AOI211_X1 g_60_138 (.ZN (n_60_138), .A (n_64_136), .B (n_67_136), .C1 (n_71_134), .C2 (n_77_131) );
AOI211_X1 g_58_139 (.ZN (n_58_139), .A (n_62_137), .B (n_68_134), .C1 (n_69_135), .C2 (n_75_132) );
AOI211_X1 g_56_140 (.ZN (n_56_140), .A (n_60_138), .B (n_66_135), .C1 (n_67_136), .C2 (n_73_133) );
AOI211_X1 g_54_141 (.ZN (n_54_141), .A (n_58_139), .B (n_64_136), .C1 (n_68_134), .C2 (n_71_134) );
AOI211_X1 g_52_142 (.ZN (n_52_142), .A (n_56_140), .B (n_62_137), .C1 (n_66_135), .C2 (n_69_135) );
AOI211_X1 g_50_141 (.ZN (n_50_141), .A (n_54_141), .B (n_60_138), .C1 (n_64_136), .C2 (n_67_136) );
AOI211_X1 g_48_142 (.ZN (n_48_142), .A (n_52_142), .B (n_58_139), .C1 (n_62_137), .C2 (n_68_134) );
AOI211_X1 g_46_143 (.ZN (n_46_143), .A (n_50_141), .B (n_56_140), .C1 (n_60_138), .C2 (n_66_135) );
AOI211_X1 g_45_145 (.ZN (n_45_145), .A (n_48_142), .B (n_54_141), .C1 (n_58_139), .C2 (n_64_136) );
AOI211_X1 g_44_147 (.ZN (n_44_147), .A (n_46_143), .B (n_52_142), .C1 (n_56_140), .C2 (n_62_137) );
AOI211_X1 g_46_148 (.ZN (n_46_148), .A (n_45_145), .B (n_50_141), .C1 (n_54_141), .C2 (n_60_138) );
AOI211_X1 g_47_146 (.ZN (n_47_146), .A (n_44_147), .B (n_48_142), .C1 (n_52_142), .C2 (n_58_139) );
AOI211_X1 g_48_144 (.ZN (n_48_144), .A (n_46_148), .B (n_46_143), .C1 (n_50_141), .C2 (n_56_140) );
AOI211_X1 g_50_143 (.ZN (n_50_143), .A (n_47_146), .B (n_45_145), .C1 (n_48_142), .C2 (n_54_141) );
AOI211_X1 g_49_145 (.ZN (n_49_145), .A (n_48_144), .B (n_44_147), .C1 (n_46_143), .C2 (n_52_142) );
AOI211_X1 g_47_144 (.ZN (n_47_144), .A (n_50_143), .B (n_46_148), .C1 (n_45_145), .C2 (n_50_141) );
AOI211_X1 g_46_146 (.ZN (n_46_146), .A (n_49_145), .B (n_47_146), .C1 (n_44_147), .C2 (n_48_142) );
AOI211_X1 g_47_148 (.ZN (n_47_148), .A (n_47_144), .B (n_48_144), .C1 (n_46_148), .C2 (n_46_143) );
AOI211_X1 g_48_146 (.ZN (n_48_146), .A (n_46_146), .B (n_50_143), .C1 (n_47_146), .C2 (n_45_145) );
AOI211_X1 g_49_148 (.ZN (n_49_148), .A (n_47_148), .B (n_49_145), .C1 (n_48_144), .C2 (n_44_147) );
AOI211_X1 g_50_150 (.ZN (n_50_150), .A (n_48_146), .B (n_47_144), .C1 (n_50_143), .C2 (n_46_148) );
AOI211_X1 g_48_149 (.ZN (n_48_149), .A (n_49_148), .B (n_46_146), .C1 (n_49_145), .C2 (n_47_146) );
AOI211_X1 g_49_147 (.ZN (n_49_147), .A (n_50_150), .B (n_47_148), .C1 (n_47_144), .C2 (n_48_144) );
AOI211_X1 g_48_145 (.ZN (n_48_145), .A (n_48_149), .B (n_48_146), .C1 (n_46_146), .C2 (n_50_143) );
AOI211_X1 g_49_143 (.ZN (n_49_143), .A (n_49_147), .B (n_49_148), .C1 (n_47_148), .C2 (n_49_145) );
AOI211_X1 g_51_142 (.ZN (n_51_142), .A (n_48_145), .B (n_50_150), .C1 (n_48_146), .C2 (n_47_144) );
AOI211_X1 g_53_141 (.ZN (n_53_141), .A (n_49_143), .B (n_48_149), .C1 (n_49_148), .C2 (n_46_146) );
AOI211_X1 g_55_140 (.ZN (n_55_140), .A (n_51_142), .B (n_49_147), .C1 (n_50_150), .C2 (n_47_148) );
AOI211_X1 g_57_139 (.ZN (n_57_139), .A (n_53_141), .B (n_48_145), .C1 (n_48_149), .C2 (n_48_146) );
AOI211_X1 g_59_138 (.ZN (n_59_138), .A (n_55_140), .B (n_49_143), .C1 (n_49_147), .C2 (n_49_148) );
AOI211_X1 g_58_140 (.ZN (n_58_140), .A (n_57_139), .B (n_51_142), .C1 (n_48_145), .C2 (n_50_150) );
AOI211_X1 g_60_139 (.ZN (n_60_139), .A (n_59_138), .B (n_53_141), .C1 (n_49_143), .C2 (n_48_149) );
AOI211_X1 g_62_138 (.ZN (n_62_138), .A (n_58_140), .B (n_55_140), .C1 (n_51_142), .C2 (n_49_147) );
AOI211_X1 g_64_137 (.ZN (n_64_137), .A (n_60_139), .B (n_57_139), .C1 (n_53_141), .C2 (n_48_145) );
AOI211_X1 g_63_139 (.ZN (n_63_139), .A (n_62_138), .B (n_59_138), .C1 (n_55_140), .C2 (n_49_143) );
AOI211_X1 g_61_138 (.ZN (n_61_138), .A (n_64_137), .B (n_58_140), .C1 (n_57_139), .C2 (n_51_142) );
AOI211_X1 g_63_137 (.ZN (n_63_137), .A (n_63_139), .B (n_60_139), .C1 (n_59_138), .C2 (n_53_141) );
AOI211_X1 g_65_136 (.ZN (n_65_136), .A (n_61_138), .B (n_62_138), .C1 (n_58_140), .C2 (n_55_140) );
AOI211_X1 g_67_135 (.ZN (n_67_135), .A (n_63_137), .B (n_64_137), .C1 (n_60_139), .C2 (n_57_139) );
AOI211_X1 g_69_134 (.ZN (n_69_134), .A (n_65_136), .B (n_63_139), .C1 (n_62_138), .C2 (n_59_138) );
AOI211_X1 g_71_133 (.ZN (n_71_133), .A (n_67_135), .B (n_61_138), .C1 (n_64_137), .C2 (n_58_140) );
AOI211_X1 g_73_132 (.ZN (n_73_132), .A (n_69_134), .B (n_63_137), .C1 (n_63_139), .C2 (n_60_139) );
AOI211_X1 g_72_134 (.ZN (n_72_134), .A (n_71_133), .B (n_65_136), .C1 (n_61_138), .C2 (n_62_138) );
AOI211_X1 g_74_133 (.ZN (n_74_133), .A (n_73_132), .B (n_67_135), .C1 (n_63_137), .C2 (n_64_137) );
AOI211_X1 g_73_135 (.ZN (n_73_135), .A (n_72_134), .B (n_69_134), .C1 (n_65_136), .C2 (n_63_139) );
AOI211_X1 g_75_134 (.ZN (n_75_134), .A (n_74_133), .B (n_71_133), .C1 (n_67_135), .C2 (n_61_138) );
AOI211_X1 g_77_133 (.ZN (n_77_133), .A (n_73_135), .B (n_73_132), .C1 (n_69_134), .C2 (n_63_137) );
AOI211_X1 g_79_132 (.ZN (n_79_132), .A (n_75_134), .B (n_72_134), .C1 (n_71_133), .C2 (n_65_136) );
AOI211_X1 g_81_131 (.ZN (n_81_131), .A (n_77_133), .B (n_74_133), .C1 (n_73_132), .C2 (n_67_135) );
AOI211_X1 g_83_130 (.ZN (n_83_130), .A (n_79_132), .B (n_73_135), .C1 (n_72_134), .C2 (n_69_134) );
AOI211_X1 g_82_132 (.ZN (n_82_132), .A (n_81_131), .B (n_75_134), .C1 (n_74_133), .C2 (n_71_133) );
AOI211_X1 g_80_131 (.ZN (n_80_131), .A (n_83_130), .B (n_77_133), .C1 (n_73_135), .C2 (n_73_132) );
AOI211_X1 g_82_130 (.ZN (n_82_130), .A (n_82_132), .B (n_79_132), .C1 (n_75_134), .C2 (n_72_134) );
AOI211_X1 g_84_129 (.ZN (n_84_129), .A (n_80_131), .B (n_81_131), .C1 (n_77_133), .C2 (n_74_133) );
AOI211_X1 g_86_128 (.ZN (n_86_128), .A (n_82_130), .B (n_83_130), .C1 (n_79_132), .C2 (n_73_135) );
AOI211_X1 g_88_127 (.ZN (n_88_127), .A (n_84_129), .B (n_82_132), .C1 (n_81_131), .C2 (n_75_134) );
AOI211_X1 g_90_126 (.ZN (n_90_126), .A (n_86_128), .B (n_80_131), .C1 (n_83_130), .C2 (n_77_133) );
AOI211_X1 g_92_125 (.ZN (n_92_125), .A (n_88_127), .B (n_82_130), .C1 (n_82_132), .C2 (n_79_132) );
AOI211_X1 g_94_124 (.ZN (n_94_124), .A (n_90_126), .B (n_84_129), .C1 (n_80_131), .C2 (n_81_131) );
AOI211_X1 g_96_123 (.ZN (n_96_123), .A (n_92_125), .B (n_86_128), .C1 (n_82_130), .C2 (n_83_130) );
AOI211_X1 g_98_122 (.ZN (n_98_122), .A (n_94_124), .B (n_88_127), .C1 (n_84_129), .C2 (n_82_132) );
AOI211_X1 g_99_124 (.ZN (n_99_124), .A (n_96_123), .B (n_90_126), .C1 (n_86_128), .C2 (n_80_131) );
AOI211_X1 g_97_125 (.ZN (n_97_125), .A (n_98_122), .B (n_92_125), .C1 (n_88_127), .C2 (n_82_130) );
AOI211_X1 g_95_126 (.ZN (n_95_126), .A (n_99_124), .B (n_94_124), .C1 (n_90_126), .C2 (n_84_129) );
AOI211_X1 g_93_127 (.ZN (n_93_127), .A (n_97_125), .B (n_96_123), .C1 (n_92_125), .C2 (n_86_128) );
AOI211_X1 g_91_128 (.ZN (n_91_128), .A (n_95_126), .B (n_98_122), .C1 (n_94_124), .C2 (n_88_127) );
AOI211_X1 g_89_129 (.ZN (n_89_129), .A (n_93_127), .B (n_99_124), .C1 (n_96_123), .C2 (n_90_126) );
AOI211_X1 g_87_130 (.ZN (n_87_130), .A (n_91_128), .B (n_97_125), .C1 (n_98_122), .C2 (n_92_125) );
AOI211_X1 g_85_131 (.ZN (n_85_131), .A (n_89_129), .B (n_95_126), .C1 (n_99_124), .C2 (n_94_124) );
AOI211_X1 g_83_132 (.ZN (n_83_132), .A (n_87_130), .B (n_93_127), .C1 (n_97_125), .C2 (n_96_123) );
AOI211_X1 g_81_133 (.ZN (n_81_133), .A (n_85_131), .B (n_91_128), .C1 (n_95_126), .C2 (n_98_122) );
AOI211_X1 g_79_134 (.ZN (n_79_134), .A (n_83_132), .B (n_89_129), .C1 (n_93_127), .C2 (n_99_124) );
AOI211_X1 g_80_132 (.ZN (n_80_132), .A (n_81_133), .B (n_87_130), .C1 (n_91_128), .C2 (n_97_125) );
AOI211_X1 g_78_133 (.ZN (n_78_133), .A (n_79_134), .B (n_85_131), .C1 (n_89_129), .C2 (n_95_126) );
AOI211_X1 g_79_131 (.ZN (n_79_131), .A (n_80_132), .B (n_83_132), .C1 (n_87_130), .C2 (n_93_127) );
AOI211_X1 g_77_132 (.ZN (n_77_132), .A (n_78_133), .B (n_81_133), .C1 (n_85_131), .C2 (n_91_128) );
AOI211_X1 g_75_133 (.ZN (n_75_133), .A (n_79_131), .B (n_79_134), .C1 (n_83_132), .C2 (n_89_129) );
AOI211_X1 g_73_134 (.ZN (n_73_134), .A (n_77_132), .B (n_80_132), .C1 (n_81_133), .C2 (n_87_130) );
AOI211_X1 g_71_135 (.ZN (n_71_135), .A (n_75_133), .B (n_78_133), .C1 (n_79_134), .C2 (n_85_131) );
AOI211_X1 g_69_136 (.ZN (n_69_136), .A (n_73_134), .B (n_79_131), .C1 (n_80_132), .C2 (n_83_132) );
AOI211_X1 g_67_137 (.ZN (n_67_137), .A (n_71_135), .B (n_77_132), .C1 (n_78_133), .C2 (n_81_133) );
AOI211_X1 g_65_138 (.ZN (n_65_138), .A (n_69_136), .B (n_75_133), .C1 (n_79_131), .C2 (n_79_134) );
AOI211_X1 g_64_140 (.ZN (n_64_140), .A (n_67_137), .B (n_73_134), .C1 (n_77_132), .C2 (n_80_132) );
AOI211_X1 g_63_138 (.ZN (n_63_138), .A (n_65_138), .B (n_71_135), .C1 (n_75_133), .C2 (n_78_133) );
AOI211_X1 g_65_137 (.ZN (n_65_137), .A (n_64_140), .B (n_69_136), .C1 (n_73_134), .C2 (n_79_131) );
AOI211_X1 g_64_139 (.ZN (n_64_139), .A (n_63_138), .B (n_67_137), .C1 (n_71_135), .C2 (n_77_132) );
AOI211_X1 g_66_138 (.ZN (n_66_138), .A (n_65_137), .B (n_65_138), .C1 (n_69_136), .C2 (n_75_133) );
AOI211_X1 g_68_137 (.ZN (n_68_137), .A (n_64_139), .B (n_64_140), .C1 (n_67_137), .C2 (n_73_134) );
AOI211_X1 g_70_136 (.ZN (n_70_136), .A (n_66_138), .B (n_63_138), .C1 (n_65_138), .C2 (n_71_135) );
AOI211_X1 g_72_135 (.ZN (n_72_135), .A (n_68_137), .B (n_65_137), .C1 (n_64_140), .C2 (n_69_136) );
AOI211_X1 g_74_134 (.ZN (n_74_134), .A (n_70_136), .B (n_64_139), .C1 (n_63_138), .C2 (n_67_137) );
AOI211_X1 g_76_133 (.ZN (n_76_133), .A (n_72_135), .B (n_66_138), .C1 (n_65_137), .C2 (n_65_138) );
AOI211_X1 g_78_132 (.ZN (n_78_132), .A (n_74_134), .B (n_68_137), .C1 (n_64_139), .C2 (n_64_140) );
AOI211_X1 g_80_133 (.ZN (n_80_133), .A (n_76_133), .B (n_70_136), .C1 (n_66_138), .C2 (n_63_138) );
AOI211_X1 g_78_134 (.ZN (n_78_134), .A (n_78_132), .B (n_72_135), .C1 (n_68_137), .C2 (n_65_137) );
AOI211_X1 g_76_135 (.ZN (n_76_135), .A (n_80_133), .B (n_74_134), .C1 (n_70_136), .C2 (n_64_139) );
AOI211_X1 g_74_136 (.ZN (n_74_136), .A (n_78_134), .B (n_76_133), .C1 (n_72_135), .C2 (n_66_138) );
AOI211_X1 g_72_137 (.ZN (n_72_137), .A (n_76_135), .B (n_78_132), .C1 (n_74_134), .C2 (n_68_137) );
AOI211_X1 g_70_138 (.ZN (n_70_138), .A (n_74_136), .B (n_80_133), .C1 (n_76_133), .C2 (n_70_136) );
AOI211_X1 g_71_136 (.ZN (n_71_136), .A (n_72_137), .B (n_78_134), .C1 (n_78_132), .C2 (n_72_135) );
AOI211_X1 g_69_137 (.ZN (n_69_137), .A (n_70_138), .B (n_76_135), .C1 (n_80_133), .C2 (n_74_134) );
AOI211_X1 g_70_135 (.ZN (n_70_135), .A (n_71_136), .B (n_74_136), .C1 (n_78_134), .C2 (n_76_133) );
AOI211_X1 g_68_136 (.ZN (n_68_136), .A (n_69_137), .B (n_72_137), .C1 (n_76_135), .C2 (n_78_132) );
AOI211_X1 g_66_137 (.ZN (n_66_137), .A (n_70_135), .B (n_70_138), .C1 (n_74_136), .C2 (n_80_133) );
AOI211_X1 g_64_138 (.ZN (n_64_138), .A (n_68_136), .B (n_71_136), .C1 (n_72_137), .C2 (n_78_134) );
AOI211_X1 g_62_139 (.ZN (n_62_139), .A (n_66_137), .B (n_69_137), .C1 (n_70_138), .C2 (n_76_135) );
AOI211_X1 g_60_140 (.ZN (n_60_140), .A (n_64_138), .B (n_70_135), .C1 (n_71_136), .C2 (n_74_136) );
AOI211_X1 g_58_141 (.ZN (n_58_141), .A (n_62_139), .B (n_68_136), .C1 (n_69_137), .C2 (n_72_137) );
AOI211_X1 g_59_139 (.ZN (n_59_139), .A (n_60_140), .B (n_66_137), .C1 (n_70_135), .C2 (n_70_138) );
AOI211_X1 g_57_140 (.ZN (n_57_140), .A (n_58_141), .B (n_64_138), .C1 (n_68_136), .C2 (n_71_136) );
AOI211_X1 g_55_141 (.ZN (n_55_141), .A (n_59_139), .B (n_62_139), .C1 (n_66_137), .C2 (n_69_137) );
AOI211_X1 g_54_143 (.ZN (n_54_143), .A (n_57_140), .B (n_60_140), .C1 (n_64_138), .C2 (n_70_135) );
AOI211_X1 g_56_142 (.ZN (n_56_142), .A (n_55_141), .B (n_58_141), .C1 (n_62_139), .C2 (n_68_136) );
AOI211_X1 g_55_144 (.ZN (n_55_144), .A (n_54_143), .B (n_59_139), .C1 (n_60_140), .C2 (n_66_137) );
AOI211_X1 g_54_142 (.ZN (n_54_142), .A (n_56_142), .B (n_57_140), .C1 (n_58_141), .C2 (n_64_138) );
AOI211_X1 g_56_141 (.ZN (n_56_141), .A (n_55_144), .B (n_55_141), .C1 (n_59_139), .C2 (n_62_139) );
AOI211_X1 g_55_143 (.ZN (n_55_143), .A (n_54_142), .B (n_54_143), .C1 (n_57_140), .C2 (n_60_140) );
AOI211_X1 g_57_142 (.ZN (n_57_142), .A (n_56_141), .B (n_56_142), .C1 (n_55_141), .C2 (n_58_141) );
AOI211_X1 g_59_141 (.ZN (n_59_141), .A (n_55_143), .B (n_55_144), .C1 (n_54_143), .C2 (n_59_139) );
AOI211_X1 g_61_140 (.ZN (n_61_140), .A (n_57_142), .B (n_54_142), .C1 (n_56_142), .C2 (n_57_140) );
AOI211_X1 g_63_141 (.ZN (n_63_141), .A (n_59_141), .B (n_56_141), .C1 (n_55_144), .C2 (n_55_141) );
AOI211_X1 g_65_140 (.ZN (n_65_140), .A (n_61_140), .B (n_55_143), .C1 (n_54_142), .C2 (n_54_143) );
AOI211_X1 g_67_139 (.ZN (n_67_139), .A (n_63_141), .B (n_57_142), .C1 (n_56_141), .C2 (n_56_142) );
AOI211_X1 g_69_138 (.ZN (n_69_138), .A (n_65_140), .B (n_59_141), .C1 (n_55_143), .C2 (n_55_144) );
AOI211_X1 g_71_137 (.ZN (n_71_137), .A (n_67_139), .B (n_61_140), .C1 (n_57_142), .C2 (n_54_142) );
AOI211_X1 g_73_136 (.ZN (n_73_136), .A (n_69_138), .B (n_63_141), .C1 (n_59_141), .C2 (n_56_141) );
AOI211_X1 g_75_135 (.ZN (n_75_135), .A (n_71_137), .B (n_65_140), .C1 (n_61_140), .C2 (n_55_143) );
AOI211_X1 g_77_134 (.ZN (n_77_134), .A (n_73_136), .B (n_67_139), .C1 (n_63_141), .C2 (n_57_142) );
AOI211_X1 g_79_133 (.ZN (n_79_133), .A (n_75_135), .B (n_69_138), .C1 (n_65_140), .C2 (n_59_141) );
AOI211_X1 g_81_132 (.ZN (n_81_132), .A (n_77_134), .B (n_71_137), .C1 (n_67_139), .C2 (n_61_140) );
AOI211_X1 g_83_131 (.ZN (n_83_131), .A (n_79_133), .B (n_73_136), .C1 (n_69_138), .C2 (n_63_141) );
AOI211_X1 g_85_130 (.ZN (n_85_130), .A (n_81_132), .B (n_75_135), .C1 (n_71_137), .C2 (n_65_140) );
AOI211_X1 g_87_129 (.ZN (n_87_129), .A (n_83_131), .B (n_77_134), .C1 (n_73_136), .C2 (n_67_139) );
AOI211_X1 g_89_128 (.ZN (n_89_128), .A (n_85_130), .B (n_79_133), .C1 (n_75_135), .C2 (n_69_138) );
AOI211_X1 g_91_127 (.ZN (n_91_127), .A (n_87_129), .B (n_81_132), .C1 (n_77_134), .C2 (n_71_137) );
AOI211_X1 g_93_126 (.ZN (n_93_126), .A (n_89_128), .B (n_83_131), .C1 (n_79_133), .C2 (n_73_136) );
AOI211_X1 g_95_125 (.ZN (n_95_125), .A (n_91_127), .B (n_85_130), .C1 (n_81_132), .C2 (n_75_135) );
AOI211_X1 g_97_124 (.ZN (n_97_124), .A (n_93_126), .B (n_87_129), .C1 (n_83_131), .C2 (n_77_134) );
AOI211_X1 g_99_123 (.ZN (n_99_123), .A (n_95_125), .B (n_89_128), .C1 (n_85_130), .C2 (n_79_133) );
AOI211_X1 g_101_122 (.ZN (n_101_122), .A (n_97_124), .B (n_91_127), .C1 (n_87_129), .C2 (n_81_132) );
AOI211_X1 g_103_121 (.ZN (n_103_121), .A (n_99_123), .B (n_93_126), .C1 (n_89_128), .C2 (n_83_131) );
AOI211_X1 g_102_123 (.ZN (n_102_123), .A (n_101_122), .B (n_95_125), .C1 (n_91_127), .C2 (n_85_130) );
AOI211_X1 g_104_122 (.ZN (n_104_122), .A (n_103_121), .B (n_97_124), .C1 (n_93_126), .C2 (n_87_129) );
AOI211_X1 g_106_121 (.ZN (n_106_121), .A (n_102_123), .B (n_99_123), .C1 (n_95_125), .C2 (n_89_128) );
AOI211_X1 g_108_120 (.ZN (n_108_120), .A (n_104_122), .B (n_101_122), .C1 (n_97_124), .C2 (n_91_127) );
AOI211_X1 g_107_122 (.ZN (n_107_122), .A (n_106_121), .B (n_103_121), .C1 (n_99_123), .C2 (n_93_126) );
AOI211_X1 g_106_120 (.ZN (n_106_120), .A (n_108_120), .B (n_102_123), .C1 (n_101_122), .C2 (n_95_125) );
AOI211_X1 g_108_119 (.ZN (n_108_119), .A (n_107_122), .B (n_104_122), .C1 (n_103_121), .C2 (n_97_124) );
AOI211_X1 g_110_118 (.ZN (n_110_118), .A (n_106_120), .B (n_106_121), .C1 (n_102_123), .C2 (n_99_123) );
AOI211_X1 g_112_117 (.ZN (n_112_117), .A (n_108_119), .B (n_108_120), .C1 (n_104_122), .C2 (n_101_122) );
AOI211_X1 g_114_116 (.ZN (n_114_116), .A (n_110_118), .B (n_107_122), .C1 (n_106_121), .C2 (n_103_121) );
AOI211_X1 g_113_118 (.ZN (n_113_118), .A (n_112_117), .B (n_106_120), .C1 (n_108_120), .C2 (n_102_123) );
AOI211_X1 g_115_117 (.ZN (n_115_117), .A (n_114_116), .B (n_108_119), .C1 (n_107_122), .C2 (n_104_122) );
AOI211_X1 g_117_118 (.ZN (n_117_118), .A (n_113_118), .B (n_110_118), .C1 (n_106_120), .C2 (n_106_121) );
AOI211_X1 g_119_117 (.ZN (n_119_117), .A (n_115_117), .B (n_112_117), .C1 (n_108_119), .C2 (n_108_120) );
AOI211_X1 g_121_116 (.ZN (n_121_116), .A (n_117_118), .B (n_114_116), .C1 (n_110_118), .C2 (n_107_122) );
AOI211_X1 g_123_115 (.ZN (n_123_115), .A (n_119_117), .B (n_113_118), .C1 (n_112_117), .C2 (n_106_120) );
AOI211_X1 g_125_114 (.ZN (n_125_114), .A (n_121_116), .B (n_115_117), .C1 (n_114_116), .C2 (n_108_119) );
AOI211_X1 g_127_113 (.ZN (n_127_113), .A (n_123_115), .B (n_117_118), .C1 (n_113_118), .C2 (n_110_118) );
AOI211_X1 g_129_112 (.ZN (n_129_112), .A (n_125_114), .B (n_119_117), .C1 (n_115_117), .C2 (n_112_117) );
AOI211_X1 g_131_111 (.ZN (n_131_111), .A (n_127_113), .B (n_121_116), .C1 (n_117_118), .C2 (n_114_116) );
AOI211_X1 g_133_110 (.ZN (n_133_110), .A (n_129_112), .B (n_123_115), .C1 (n_119_117), .C2 (n_113_118) );
AOI211_X1 g_135_109 (.ZN (n_135_109), .A (n_131_111), .B (n_125_114), .C1 (n_121_116), .C2 (n_115_117) );
AOI211_X1 g_134_111 (.ZN (n_134_111), .A (n_133_110), .B (n_127_113), .C1 (n_123_115), .C2 (n_117_118) );
AOI211_X1 g_136_110 (.ZN (n_136_110), .A (n_135_109), .B (n_129_112), .C1 (n_125_114), .C2 (n_119_117) );
AOI211_X1 g_138_109 (.ZN (n_138_109), .A (n_134_111), .B (n_131_111), .C1 (n_127_113), .C2 (n_121_116) );
AOI211_X1 g_140_108 (.ZN (n_140_108), .A (n_136_110), .B (n_133_110), .C1 (n_129_112), .C2 (n_123_115) );
AOI211_X1 g_142_107 (.ZN (n_142_107), .A (n_138_109), .B (n_135_109), .C1 (n_131_111), .C2 (n_125_114) );
AOI211_X1 g_144_106 (.ZN (n_144_106), .A (n_140_108), .B (n_134_111), .C1 (n_133_110), .C2 (n_127_113) );
AOI211_X1 g_146_107 (.ZN (n_146_107), .A (n_142_107), .B (n_136_110), .C1 (n_135_109), .C2 (n_129_112) );
AOI211_X1 g_144_108 (.ZN (n_144_108), .A (n_144_106), .B (n_138_109), .C1 (n_134_111), .C2 (n_131_111) );
AOI211_X1 g_142_109 (.ZN (n_142_109), .A (n_146_107), .B (n_140_108), .C1 (n_136_110), .C2 (n_133_110) );
AOI211_X1 g_143_107 (.ZN (n_143_107), .A (n_144_108), .B (n_142_107), .C1 (n_138_109), .C2 (n_135_109) );
AOI211_X1 g_144_109 (.ZN (n_144_109), .A (n_142_109), .B (n_144_106), .C1 (n_140_108), .C2 (n_134_111) );
AOI211_X1 g_146_110 (.ZN (n_146_110), .A (n_143_107), .B (n_146_107), .C1 (n_142_107), .C2 (n_136_110) );
AOI211_X1 g_145_108 (.ZN (n_145_108), .A (n_144_109), .B (n_144_108), .C1 (n_144_106), .C2 (n_138_109) );
AOI211_X1 g_147_109 (.ZN (n_147_109), .A (n_146_110), .B (n_142_109), .C1 (n_146_107), .C2 (n_140_108) );
AOI211_X1 g_148_111 (.ZN (n_148_111), .A (n_145_108), .B (n_143_107), .C1 (n_144_108), .C2 (n_142_107) );
AOI211_X1 g_146_112 (.ZN (n_146_112), .A (n_147_109), .B (n_144_109), .C1 (n_142_109), .C2 (n_144_106) );
AOI211_X1 g_145_110 (.ZN (n_145_110), .A (n_148_111), .B (n_146_110), .C1 (n_143_107), .C2 (n_146_107) );
AOI211_X1 g_143_109 (.ZN (n_143_109), .A (n_146_112), .B (n_145_108), .C1 (n_144_109), .C2 (n_144_108) );
AOI211_X1 g_141_108 (.ZN (n_141_108), .A (n_145_110), .B (n_147_109), .C1 (n_146_110), .C2 (n_142_109) );
AOI211_X1 g_139_109 (.ZN (n_139_109), .A (n_143_109), .B (n_148_111), .C1 (n_145_108), .C2 (n_143_107) );
AOI211_X1 g_137_110 (.ZN (n_137_110), .A (n_141_108), .B (n_146_112), .C1 (n_147_109), .C2 (n_144_109) );
AOI211_X1 g_135_111 (.ZN (n_135_111), .A (n_139_109), .B (n_145_110), .C1 (n_148_111), .C2 (n_146_110) );
AOI211_X1 g_133_112 (.ZN (n_133_112), .A (n_137_110), .B (n_143_109), .C1 (n_146_112), .C2 (n_145_108) );
AOI211_X1 g_131_113 (.ZN (n_131_113), .A (n_135_111), .B (n_141_108), .C1 (n_145_110), .C2 (n_147_109) );
AOI211_X1 g_129_114 (.ZN (n_129_114), .A (n_133_112), .B (n_139_109), .C1 (n_143_109), .C2 (n_148_111) );
AOI211_X1 g_128_116 (.ZN (n_128_116), .A (n_131_113), .B (n_137_110), .C1 (n_141_108), .C2 (n_146_112) );
AOI211_X1 g_126_115 (.ZN (n_126_115), .A (n_129_114), .B (n_135_111), .C1 (n_139_109), .C2 (n_145_110) );
AOI211_X1 g_128_114 (.ZN (n_128_114), .A (n_128_116), .B (n_133_112), .C1 (n_137_110), .C2 (n_143_109) );
AOI211_X1 g_130_113 (.ZN (n_130_113), .A (n_126_115), .B (n_131_113), .C1 (n_135_111), .C2 (n_141_108) );
AOI211_X1 g_132_112 (.ZN (n_132_112), .A (n_128_114), .B (n_129_114), .C1 (n_133_112), .C2 (n_139_109) );
AOI211_X1 g_131_114 (.ZN (n_131_114), .A (n_130_113), .B (n_128_116), .C1 (n_131_113), .C2 (n_137_110) );
AOI211_X1 g_133_113 (.ZN (n_133_113), .A (n_132_112), .B (n_126_115), .C1 (n_129_114), .C2 (n_135_111) );
AOI211_X1 g_135_112 (.ZN (n_135_112), .A (n_131_114), .B (n_128_114), .C1 (n_128_116), .C2 (n_133_112) );
AOI211_X1 g_137_111 (.ZN (n_137_111), .A (n_133_113), .B (n_130_113), .C1 (n_126_115), .C2 (n_131_113) );
AOI211_X1 g_139_110 (.ZN (n_139_110), .A (n_135_112), .B (n_132_112), .C1 (n_128_114), .C2 (n_129_114) );
AOI211_X1 g_141_109 (.ZN (n_141_109), .A (n_137_111), .B (n_131_114), .C1 (n_130_113), .C2 (n_128_116) );
AOI211_X1 g_143_108 (.ZN (n_143_108), .A (n_139_110), .B (n_133_113), .C1 (n_132_112), .C2 (n_126_115) );
AOI211_X1 g_145_109 (.ZN (n_145_109), .A (n_141_109), .B (n_135_112), .C1 (n_131_114), .C2 (n_128_114) );
AOI211_X1 g_143_110 (.ZN (n_143_110), .A (n_143_108), .B (n_137_111), .C1 (n_133_113), .C2 (n_130_113) );
AOI211_X1 g_141_111 (.ZN (n_141_111), .A (n_145_109), .B (n_139_110), .C1 (n_135_112), .C2 (n_132_112) );
AOI211_X1 g_140_109 (.ZN (n_140_109), .A (n_143_110), .B (n_141_109), .C1 (n_137_111), .C2 (n_131_114) );
AOI211_X1 g_138_110 (.ZN (n_138_110), .A (n_141_111), .B (n_143_108), .C1 (n_139_110), .C2 (n_133_113) );
AOI211_X1 g_136_111 (.ZN (n_136_111), .A (n_140_109), .B (n_145_109), .C1 (n_141_109), .C2 (n_135_112) );
AOI211_X1 g_134_112 (.ZN (n_134_112), .A (n_138_110), .B (n_143_110), .C1 (n_143_108), .C2 (n_137_111) );
AOI211_X1 g_132_113 (.ZN (n_132_113), .A (n_136_111), .B (n_141_111), .C1 (n_145_109), .C2 (n_139_110) );
AOI211_X1 g_130_114 (.ZN (n_130_114), .A (n_134_112), .B (n_140_109), .C1 (n_143_110), .C2 (n_141_109) );
AOI211_X1 g_128_115 (.ZN (n_128_115), .A (n_132_113), .B (n_138_110), .C1 (n_141_111), .C2 (n_143_108) );
AOI211_X1 g_126_116 (.ZN (n_126_116), .A (n_130_114), .B (n_136_111), .C1 (n_140_109), .C2 (n_145_109) );
AOI211_X1 g_124_117 (.ZN (n_124_117), .A (n_128_115), .B (n_134_112), .C1 (n_138_110), .C2 (n_143_110) );
AOI211_X1 g_122_118 (.ZN (n_122_118), .A (n_126_116), .B (n_132_113), .C1 (n_136_111), .C2 (n_141_111) );
AOI211_X1 g_120_119 (.ZN (n_120_119), .A (n_124_117), .B (n_130_114), .C1 (n_134_112), .C2 (n_140_109) );
AOI211_X1 g_121_117 (.ZN (n_121_117), .A (n_122_118), .B (n_128_115), .C1 (n_132_113), .C2 (n_138_110) );
AOI211_X1 g_119_116 (.ZN (n_119_116), .A (n_120_119), .B (n_126_116), .C1 (n_130_114), .C2 (n_136_111) );
AOI211_X1 g_117_115 (.ZN (n_117_115), .A (n_121_117), .B (n_124_117), .C1 (n_128_115), .C2 (n_134_112) );
AOI211_X1 g_115_116 (.ZN (n_115_116), .A (n_119_116), .B (n_122_118), .C1 (n_126_116), .C2 (n_132_113) );
AOI211_X1 g_113_117 (.ZN (n_113_117), .A (n_117_115), .B (n_120_119), .C1 (n_124_117), .C2 (n_130_114) );
AOI211_X1 g_111_118 (.ZN (n_111_118), .A (n_115_116), .B (n_121_117), .C1 (n_122_118), .C2 (n_128_115) );
AOI211_X1 g_109_119 (.ZN (n_109_119), .A (n_113_117), .B (n_119_116), .C1 (n_120_119), .C2 (n_126_116) );
AOI211_X1 g_107_120 (.ZN (n_107_120), .A (n_111_118), .B (n_117_115), .C1 (n_121_117), .C2 (n_124_117) );
AOI211_X1 g_105_121 (.ZN (n_105_121), .A (n_109_119), .B (n_115_116), .C1 (n_119_116), .C2 (n_122_118) );
AOI211_X1 g_103_122 (.ZN (n_103_122), .A (n_107_120), .B (n_113_117), .C1 (n_117_115), .C2 (n_120_119) );
AOI211_X1 g_105_123 (.ZN (n_105_123), .A (n_105_121), .B (n_111_118), .C1 (n_115_116), .C2 (n_121_117) );
AOI211_X1 g_104_121 (.ZN (n_104_121), .A (n_103_122), .B (n_109_119), .C1 (n_113_117), .C2 (n_119_116) );
AOI211_X1 g_102_122 (.ZN (n_102_122), .A (n_105_123), .B (n_107_120), .C1 (n_111_118), .C2 (n_117_115) );
AOI211_X1 g_100_123 (.ZN (n_100_123), .A (n_104_121), .B (n_105_121), .C1 (n_109_119), .C2 (n_115_116) );
AOI211_X1 g_98_124 (.ZN (n_98_124), .A (n_102_122), .B (n_103_122), .C1 (n_107_120), .C2 (n_113_117) );
AOI211_X1 g_96_125 (.ZN (n_96_125), .A (n_100_123), .B (n_105_123), .C1 (n_105_121), .C2 (n_111_118) );
AOI211_X1 g_94_126 (.ZN (n_94_126), .A (n_98_124), .B (n_104_121), .C1 (n_103_122), .C2 (n_109_119) );
AOI211_X1 g_92_127 (.ZN (n_92_127), .A (n_96_125), .B (n_102_122), .C1 (n_105_123), .C2 (n_107_120) );
AOI211_X1 g_90_128 (.ZN (n_90_128), .A (n_94_126), .B (n_100_123), .C1 (n_104_121), .C2 (n_105_121) );
AOI211_X1 g_88_129 (.ZN (n_88_129), .A (n_92_127), .B (n_98_124), .C1 (n_102_122), .C2 (n_103_122) );
AOI211_X1 g_86_130 (.ZN (n_86_130), .A (n_90_128), .B (n_96_125), .C1 (n_100_123), .C2 (n_105_123) );
AOI211_X1 g_84_131 (.ZN (n_84_131), .A (n_88_129), .B (n_94_126), .C1 (n_98_124), .C2 (n_104_121) );
AOI211_X1 g_83_133 (.ZN (n_83_133), .A (n_86_130), .B (n_92_127), .C1 (n_96_125), .C2 (n_102_122) );
AOI211_X1 g_85_132 (.ZN (n_85_132), .A (n_84_131), .B (n_90_128), .C1 (n_94_126), .C2 (n_100_123) );
AOI211_X1 g_87_131 (.ZN (n_87_131), .A (n_83_133), .B (n_88_129), .C1 (n_92_127), .C2 (n_98_124) );
AOI211_X1 g_89_130 (.ZN (n_89_130), .A (n_85_132), .B (n_86_130), .C1 (n_90_128), .C2 (n_96_125) );
AOI211_X1 g_91_129 (.ZN (n_91_129), .A (n_87_131), .B (n_84_131), .C1 (n_88_129), .C2 (n_94_126) );
AOI211_X1 g_93_128 (.ZN (n_93_128), .A (n_89_130), .B (n_83_133), .C1 (n_86_130), .C2 (n_92_127) );
AOI211_X1 g_95_127 (.ZN (n_95_127), .A (n_91_129), .B (n_85_132), .C1 (n_84_131), .C2 (n_90_128) );
AOI211_X1 g_97_126 (.ZN (n_97_126), .A (n_93_128), .B (n_87_131), .C1 (n_83_133), .C2 (n_88_129) );
AOI211_X1 g_99_125 (.ZN (n_99_125), .A (n_95_127), .B (n_89_130), .C1 (n_85_132), .C2 (n_86_130) );
AOI211_X1 g_101_124 (.ZN (n_101_124), .A (n_97_126), .B (n_91_129), .C1 (n_87_131), .C2 (n_84_131) );
AOI211_X1 g_103_123 (.ZN (n_103_123), .A (n_99_125), .B (n_93_128), .C1 (n_89_130), .C2 (n_83_133) );
AOI211_X1 g_105_122 (.ZN (n_105_122), .A (n_101_124), .B (n_95_127), .C1 (n_91_129), .C2 (n_85_132) );
AOI211_X1 g_107_121 (.ZN (n_107_121), .A (n_103_123), .B (n_97_126), .C1 (n_93_128), .C2 (n_87_131) );
AOI211_X1 g_109_120 (.ZN (n_109_120), .A (n_105_122), .B (n_99_125), .C1 (n_95_127), .C2 (n_89_130) );
AOI211_X1 g_111_119 (.ZN (n_111_119), .A (n_107_121), .B (n_101_124), .C1 (n_97_126), .C2 (n_91_129) );
AOI211_X1 g_110_121 (.ZN (n_110_121), .A (n_109_120), .B (n_103_123), .C1 (n_99_125), .C2 (n_93_128) );
AOI211_X1 g_112_120 (.ZN (n_112_120), .A (n_111_119), .B (n_105_122), .C1 (n_101_124), .C2 (n_95_127) );
AOI211_X1 g_114_119 (.ZN (n_114_119), .A (n_110_121), .B (n_107_121), .C1 (n_103_123), .C2 (n_97_126) );
AOI211_X1 g_116_118 (.ZN (n_116_118), .A (n_112_120), .B (n_109_120), .C1 (n_105_122), .C2 (n_99_125) );
AOI211_X1 g_118_117 (.ZN (n_118_117), .A (n_114_119), .B (n_111_119), .C1 (n_107_121), .C2 (n_101_124) );
AOI211_X1 g_119_119 (.ZN (n_119_119), .A (n_116_118), .B (n_110_121), .C1 (n_109_120), .C2 (n_103_123) );
AOI211_X1 g_121_118 (.ZN (n_121_118), .A (n_118_117), .B (n_112_120), .C1 (n_111_119), .C2 (n_105_122) );
AOI211_X1 g_123_117 (.ZN (n_123_117), .A (n_119_119), .B (n_114_119), .C1 (n_110_121), .C2 (n_107_121) );
AOI211_X1 g_125_116 (.ZN (n_125_116), .A (n_121_118), .B (n_116_118), .C1 (n_112_120), .C2 (n_109_120) );
AOI211_X1 g_127_117 (.ZN (n_127_117), .A (n_123_117), .B (n_118_117), .C1 (n_114_119), .C2 (n_111_119) );
AOI211_X1 g_129_116 (.ZN (n_129_116), .A (n_125_116), .B (n_119_119), .C1 (n_116_118), .C2 (n_110_121) );
AOI211_X1 g_131_115 (.ZN (n_131_115), .A (n_127_117), .B (n_121_118), .C1 (n_118_117), .C2 (n_112_120) );
AOI211_X1 g_133_114 (.ZN (n_133_114), .A (n_129_116), .B (n_123_117), .C1 (n_119_119), .C2 (n_114_119) );
AOI211_X1 g_135_113 (.ZN (n_135_113), .A (n_131_115), .B (n_125_116), .C1 (n_121_118), .C2 (n_116_118) );
AOI211_X1 g_137_112 (.ZN (n_137_112), .A (n_133_114), .B (n_127_117), .C1 (n_123_117), .C2 (n_118_117) );
AOI211_X1 g_139_111 (.ZN (n_139_111), .A (n_135_113), .B (n_129_116), .C1 (n_125_116), .C2 (n_119_119) );
AOI211_X1 g_141_110 (.ZN (n_141_110), .A (n_137_112), .B (n_131_115), .C1 (n_127_117), .C2 (n_121_118) );
AOI211_X1 g_143_111 (.ZN (n_143_111), .A (n_139_111), .B (n_133_114), .C1 (n_129_116), .C2 (n_123_117) );
AOI211_X1 g_144_113 (.ZN (n_144_113), .A (n_141_110), .B (n_135_113), .C1 (n_131_115), .C2 (n_125_116) );
AOI211_X1 g_146_114 (.ZN (n_146_114), .A (n_143_111), .B (n_137_112), .C1 (n_133_114), .C2 (n_127_117) );
AOI211_X1 g_148_115 (.ZN (n_148_115), .A (n_144_113), .B (n_139_111), .C1 (n_135_113), .C2 (n_129_116) );
AOI211_X1 g_147_113 (.ZN (n_147_113), .A (n_146_114), .B (n_141_110), .C1 (n_137_112), .C2 (n_131_115) );
AOI211_X1 g_146_111 (.ZN (n_146_111), .A (n_148_115), .B (n_143_111), .C1 (n_139_111), .C2 (n_133_114) );
AOI211_X1 g_144_110 (.ZN (n_144_110), .A (n_147_113), .B (n_144_113), .C1 (n_141_110), .C2 (n_135_113) );
AOI211_X1 g_145_112 (.ZN (n_145_112), .A (n_146_111), .B (n_146_114), .C1 (n_143_111), .C2 (n_137_112) );
AOI211_X1 g_144_114 (.ZN (n_144_114), .A (n_144_110), .B (n_148_115), .C1 (n_144_113), .C2 (n_139_111) );
AOI211_X1 g_143_112 (.ZN (n_143_112), .A (n_145_112), .B (n_147_113), .C1 (n_146_114), .C2 (n_141_110) );
AOI211_X1 g_142_110 (.ZN (n_142_110), .A (n_144_114), .B (n_146_111), .C1 (n_148_115), .C2 (n_143_111) );
AOI211_X1 g_144_111 (.ZN (n_144_111), .A (n_143_112), .B (n_144_110), .C1 (n_147_113), .C2 (n_144_113) );
AOI211_X1 g_145_113 (.ZN (n_145_113), .A (n_142_110), .B (n_145_112), .C1 (n_146_111), .C2 (n_146_114) );
AOI211_X1 g_146_115 (.ZN (n_146_115), .A (n_144_111), .B (n_144_114), .C1 (n_144_110), .C2 (n_148_115) );
AOI211_X1 g_147_117 (.ZN (n_147_117), .A (n_145_113), .B (n_143_112), .C1 (n_145_112), .C2 (n_147_113) );
AOI211_X1 g_148_119 (.ZN (n_148_119), .A (n_146_115), .B (n_142_110), .C1 (n_144_114), .C2 (n_146_111) );
AOI211_X1 g_146_118 (.ZN (n_146_118), .A (n_147_117), .B (n_144_111), .C1 (n_143_112), .C2 (n_144_110) );
AOI211_X1 g_145_116 (.ZN (n_145_116), .A (n_148_119), .B (n_145_113), .C1 (n_142_110), .C2 (n_145_112) );
AOI211_X1 g_143_115 (.ZN (n_143_115), .A (n_146_118), .B (n_146_115), .C1 (n_144_111), .C2 (n_144_114) );
AOI211_X1 g_145_114 (.ZN (n_145_114), .A (n_145_116), .B (n_147_117), .C1 (n_145_113), .C2 (n_143_112) );
AOI211_X1 g_144_112 (.ZN (n_144_112), .A (n_143_115), .B (n_148_119), .C1 (n_146_115), .C2 (n_142_110) );
AOI211_X1 g_142_113 (.ZN (n_142_113), .A (n_145_114), .B (n_146_118), .C1 (n_147_117), .C2 (n_144_111) );
AOI211_X1 g_140_112 (.ZN (n_140_112), .A (n_144_112), .B (n_145_116), .C1 (n_148_119), .C2 (n_145_113) );
AOI211_X1 g_142_111 (.ZN (n_142_111), .A (n_142_113), .B (n_143_115), .C1 (n_146_118), .C2 (n_146_115) );
AOI211_X1 g_140_110 (.ZN (n_140_110), .A (n_140_112), .B (n_145_114), .C1 (n_145_116), .C2 (n_147_117) );
AOI211_X1 g_138_111 (.ZN (n_138_111), .A (n_142_111), .B (n_144_112), .C1 (n_143_115), .C2 (n_148_119) );
AOI211_X1 g_136_112 (.ZN (n_136_112), .A (n_140_110), .B (n_142_113), .C1 (n_145_114), .C2 (n_146_118) );
AOI211_X1 g_134_113 (.ZN (n_134_113), .A (n_138_111), .B (n_140_112), .C1 (n_144_112), .C2 (n_145_116) );
AOI211_X1 g_132_114 (.ZN (n_132_114), .A (n_136_112), .B (n_142_111), .C1 (n_142_113), .C2 (n_143_115) );
AOI211_X1 g_130_115 (.ZN (n_130_115), .A (n_134_113), .B (n_140_110), .C1 (n_140_112), .C2 (n_145_114) );
AOI211_X1 g_132_116 (.ZN (n_132_116), .A (n_132_114), .B (n_138_111), .C1 (n_142_111), .C2 (n_144_112) );
AOI211_X1 g_134_115 (.ZN (n_134_115), .A (n_130_115), .B (n_136_112), .C1 (n_140_110), .C2 (n_142_113) );
AOI211_X1 g_136_114 (.ZN (n_136_114), .A (n_132_116), .B (n_134_113), .C1 (n_138_111), .C2 (n_140_112) );
AOI211_X1 g_138_113 (.ZN (n_138_113), .A (n_134_115), .B (n_132_114), .C1 (n_136_112), .C2 (n_142_111) );
AOI211_X1 g_140_114 (.ZN (n_140_114), .A (n_136_114), .B (n_130_115), .C1 (n_134_113), .C2 (n_140_110) );
AOI211_X1 g_141_112 (.ZN (n_141_112), .A (n_138_113), .B (n_132_116), .C1 (n_132_114), .C2 (n_138_111) );
AOI211_X1 g_143_113 (.ZN (n_143_113), .A (n_140_114), .B (n_134_115), .C1 (n_130_115), .C2 (n_136_112) );
AOI211_X1 g_141_114 (.ZN (n_141_114), .A (n_141_112), .B (n_136_114), .C1 (n_132_116), .C2 (n_134_113) );
AOI211_X1 g_142_112 (.ZN (n_142_112), .A (n_143_113), .B (n_138_113), .C1 (n_134_115), .C2 (n_132_114) );
AOI211_X1 g_140_111 (.ZN (n_140_111), .A (n_141_114), .B (n_140_114), .C1 (n_136_114), .C2 (n_130_115) );
AOI211_X1 g_139_113 (.ZN (n_139_113), .A (n_142_112), .B (n_141_112), .C1 (n_138_113), .C2 (n_132_116) );
AOI211_X1 g_137_114 (.ZN (n_137_114), .A (n_140_111), .B (n_143_113), .C1 (n_140_114), .C2 (n_134_115) );
AOI211_X1 g_138_112 (.ZN (n_138_112), .A (n_139_113), .B (n_141_114), .C1 (n_141_112), .C2 (n_136_114) );
AOI211_X1 g_136_113 (.ZN (n_136_113), .A (n_137_114), .B (n_142_112), .C1 (n_143_113), .C2 (n_138_113) );
AOI211_X1 g_134_114 (.ZN (n_134_114), .A (n_138_112), .B (n_140_111), .C1 (n_141_114), .C2 (n_140_114) );
AOI211_X1 g_132_115 (.ZN (n_132_115), .A (n_136_113), .B (n_139_113), .C1 (n_142_112), .C2 (n_141_112) );
AOI211_X1 g_130_116 (.ZN (n_130_116), .A (n_134_114), .B (n_137_114), .C1 (n_140_111), .C2 (n_143_113) );
AOI211_X1 g_128_117 (.ZN (n_128_117), .A (n_132_115), .B (n_138_112), .C1 (n_139_113), .C2 (n_141_114) );
AOI211_X1 g_129_115 (.ZN (n_129_115), .A (n_130_116), .B (n_136_113), .C1 (n_137_114), .C2 (n_142_112) );
AOI211_X1 g_127_116 (.ZN (n_127_116), .A (n_128_117), .B (n_134_114), .C1 (n_138_112), .C2 (n_140_111) );
AOI211_X1 g_125_117 (.ZN (n_125_117), .A (n_129_115), .B (n_132_115), .C1 (n_136_113), .C2 (n_139_113) );
AOI211_X1 g_123_118 (.ZN (n_123_118), .A (n_127_116), .B (n_130_116), .C1 (n_134_114), .C2 (n_137_114) );
AOI211_X1 g_124_116 (.ZN (n_124_116), .A (n_125_117), .B (n_128_117), .C1 (n_132_115), .C2 (n_138_112) );
AOI211_X1 g_122_117 (.ZN (n_122_117), .A (n_123_118), .B (n_129_115), .C1 (n_130_116), .C2 (n_136_113) );
AOI211_X1 g_120_118 (.ZN (n_120_118), .A (n_124_116), .B (n_127_116), .C1 (n_128_117), .C2 (n_134_114) );
AOI211_X1 g_118_119 (.ZN (n_118_119), .A (n_122_117), .B (n_125_117), .C1 (n_129_115), .C2 (n_132_115) );
AOI211_X1 g_117_117 (.ZN (n_117_117), .A (n_120_118), .B (n_123_118), .C1 (n_127_116), .C2 (n_130_116) );
AOI211_X1 g_115_118 (.ZN (n_115_118), .A (n_118_119), .B (n_124_116), .C1 (n_125_117), .C2 (n_128_117) );
AOI211_X1 g_113_119 (.ZN (n_113_119), .A (n_117_117), .B (n_122_117), .C1 (n_123_118), .C2 (n_129_115) );
AOI211_X1 g_111_120 (.ZN (n_111_120), .A (n_115_118), .B (n_120_118), .C1 (n_124_116), .C2 (n_127_116) );
AOI211_X1 g_109_121 (.ZN (n_109_121), .A (n_113_119), .B (n_118_119), .C1 (n_122_117), .C2 (n_125_117) );
AOI211_X1 g_108_123 (.ZN (n_108_123), .A (n_111_120), .B (n_117_117), .C1 (n_120_118), .C2 (n_123_118) );
AOI211_X1 g_106_122 (.ZN (n_106_122), .A (n_109_121), .B (n_115_118), .C1 (n_118_119), .C2 (n_124_116) );
AOI211_X1 g_108_121 (.ZN (n_108_121), .A (n_108_123), .B (n_113_119), .C1 (n_117_117), .C2 (n_122_117) );
AOI211_X1 g_110_120 (.ZN (n_110_120), .A (n_106_122), .B (n_111_120), .C1 (n_115_118), .C2 (n_120_118) );
AOI211_X1 g_112_119 (.ZN (n_112_119), .A (n_108_121), .B (n_109_121), .C1 (n_113_119), .C2 (n_118_119) );
AOI211_X1 g_114_118 (.ZN (n_114_118), .A (n_110_120), .B (n_108_123), .C1 (n_111_120), .C2 (n_117_117) );
AOI211_X1 g_116_117 (.ZN (n_116_117), .A (n_112_119), .B (n_106_122), .C1 (n_109_121), .C2 (n_115_118) );
AOI211_X1 g_118_118 (.ZN (n_118_118), .A (n_114_118), .B (n_108_121), .C1 (n_108_123), .C2 (n_113_119) );
AOI211_X1 g_116_119 (.ZN (n_116_119), .A (n_116_117), .B (n_110_120), .C1 (n_106_122), .C2 (n_111_120) );
AOI211_X1 g_114_120 (.ZN (n_114_120), .A (n_118_118), .B (n_112_119), .C1 (n_108_121), .C2 (n_109_121) );
AOI211_X1 g_112_121 (.ZN (n_112_121), .A (n_116_119), .B (n_114_118), .C1 (n_110_120), .C2 (n_108_123) );
AOI211_X1 g_110_122 (.ZN (n_110_122), .A (n_114_120), .B (n_116_117), .C1 (n_112_119), .C2 (n_106_122) );
AOI211_X1 g_109_124 (.ZN (n_109_124), .A (n_112_121), .B (n_118_118), .C1 (n_114_118), .C2 (n_108_121) );
AOI211_X1 g_108_122 (.ZN (n_108_122), .A (n_110_122), .B (n_116_119), .C1 (n_116_117), .C2 (n_110_120) );
AOI211_X1 g_106_123 (.ZN (n_106_123), .A (n_109_124), .B (n_114_120), .C1 (n_118_118), .C2 (n_112_119) );
AOI211_X1 g_104_124 (.ZN (n_104_124), .A (n_108_122), .B (n_112_121), .C1 (n_116_119), .C2 (n_114_118) );
AOI211_X1 g_102_125 (.ZN (n_102_125), .A (n_106_123), .B (n_110_122), .C1 (n_114_120), .C2 (n_116_117) );
AOI211_X1 g_100_124 (.ZN (n_100_124), .A (n_104_124), .B (n_109_124), .C1 (n_112_121), .C2 (n_118_118) );
AOI211_X1 g_98_125 (.ZN (n_98_125), .A (n_102_125), .B (n_108_122), .C1 (n_110_122), .C2 (n_116_119) );
AOI211_X1 g_96_126 (.ZN (n_96_126), .A (n_100_124), .B (n_106_123), .C1 (n_109_124), .C2 (n_114_120) );
AOI211_X1 g_94_127 (.ZN (n_94_127), .A (n_98_125), .B (n_104_124), .C1 (n_108_122), .C2 (n_112_121) );
AOI211_X1 g_92_128 (.ZN (n_92_128), .A (n_96_126), .B (n_102_125), .C1 (n_106_123), .C2 (n_110_122) );
AOI211_X1 g_90_129 (.ZN (n_90_129), .A (n_94_127), .B (n_100_124), .C1 (n_104_124), .C2 (n_109_124) );
AOI211_X1 g_88_130 (.ZN (n_88_130), .A (n_92_128), .B (n_98_125), .C1 (n_102_125), .C2 (n_108_122) );
AOI211_X1 g_86_131 (.ZN (n_86_131), .A (n_90_129), .B (n_96_126), .C1 (n_100_124), .C2 (n_106_123) );
AOI211_X1 g_84_132 (.ZN (n_84_132), .A (n_88_130), .B (n_94_127), .C1 (n_98_125), .C2 (n_104_124) );
AOI211_X1 g_82_133 (.ZN (n_82_133), .A (n_86_131), .B (n_92_128), .C1 (n_96_126), .C2 (n_102_125) );
AOI211_X1 g_80_134 (.ZN (n_80_134), .A (n_84_132), .B (n_90_129), .C1 (n_94_127), .C2 (n_100_124) );
AOI211_X1 g_78_135 (.ZN (n_78_135), .A (n_82_133), .B (n_88_130), .C1 (n_92_128), .C2 (n_98_125) );
AOI211_X1 g_76_134 (.ZN (n_76_134), .A (n_80_134), .B (n_86_131), .C1 (n_90_129), .C2 (n_96_126) );
AOI211_X1 g_74_135 (.ZN (n_74_135), .A (n_78_135), .B (n_84_132), .C1 (n_88_130), .C2 (n_94_127) );
AOI211_X1 g_72_136 (.ZN (n_72_136), .A (n_76_134), .B (n_82_133), .C1 (n_86_131), .C2 (n_92_128) );
AOI211_X1 g_70_137 (.ZN (n_70_137), .A (n_74_135), .B (n_80_134), .C1 (n_84_132), .C2 (n_90_129) );
AOI211_X1 g_68_138 (.ZN (n_68_138), .A (n_72_136), .B (n_78_135), .C1 (n_82_133), .C2 (n_88_130) );
AOI211_X1 g_66_139 (.ZN (n_66_139), .A (n_70_137), .B (n_76_134), .C1 (n_80_134), .C2 (n_86_131) );
AOI211_X1 g_65_141 (.ZN (n_65_141), .A (n_68_138), .B (n_74_135), .C1 (n_78_135), .C2 (n_84_132) );
AOI211_X1 g_67_140 (.ZN (n_67_140), .A (n_66_139), .B (n_72_136), .C1 (n_76_134), .C2 (n_82_133) );
AOI211_X1 g_65_139 (.ZN (n_65_139), .A (n_65_141), .B (n_70_137), .C1 (n_74_135), .C2 (n_80_134) );
AOI211_X1 g_67_138 (.ZN (n_67_138), .A (n_67_140), .B (n_68_138), .C1 (n_72_136), .C2 (n_78_135) );
AOI211_X1 g_69_139 (.ZN (n_69_139), .A (n_65_139), .B (n_66_139), .C1 (n_70_137), .C2 (n_76_134) );
AOI211_X1 g_71_138 (.ZN (n_71_138), .A (n_67_138), .B (n_65_141), .C1 (n_68_138), .C2 (n_74_135) );
AOI211_X1 g_73_137 (.ZN (n_73_137), .A (n_69_139), .B (n_67_140), .C1 (n_66_139), .C2 (n_72_136) );
AOI211_X1 g_75_136 (.ZN (n_75_136), .A (n_71_138), .B (n_65_139), .C1 (n_65_141), .C2 (n_70_137) );
AOI211_X1 g_77_135 (.ZN (n_77_135), .A (n_73_137), .B (n_67_138), .C1 (n_67_140), .C2 (n_68_138) );
AOI211_X1 g_76_137 (.ZN (n_76_137), .A (n_75_136), .B (n_69_139), .C1 (n_65_139), .C2 (n_66_139) );
AOI211_X1 g_78_136 (.ZN (n_78_136), .A (n_77_135), .B (n_71_138), .C1 (n_67_138), .C2 (n_65_141) );
AOI211_X1 g_80_135 (.ZN (n_80_135), .A (n_76_137), .B (n_73_137), .C1 (n_69_139), .C2 (n_67_140) );
AOI211_X1 g_82_134 (.ZN (n_82_134), .A (n_78_136), .B (n_75_136), .C1 (n_71_138), .C2 (n_65_139) );
AOI211_X1 g_84_133 (.ZN (n_84_133), .A (n_80_135), .B (n_77_135), .C1 (n_73_137), .C2 (n_67_138) );
AOI211_X1 g_86_132 (.ZN (n_86_132), .A (n_82_134), .B (n_76_137), .C1 (n_75_136), .C2 (n_69_139) );
AOI211_X1 g_88_131 (.ZN (n_88_131), .A (n_84_133), .B (n_78_136), .C1 (n_77_135), .C2 (n_71_138) );
AOI211_X1 g_90_130 (.ZN (n_90_130), .A (n_86_132), .B (n_80_135), .C1 (n_76_137), .C2 (n_73_137) );
AOI211_X1 g_92_129 (.ZN (n_92_129), .A (n_88_131), .B (n_82_134), .C1 (n_78_136), .C2 (n_75_136) );
AOI211_X1 g_94_128 (.ZN (n_94_128), .A (n_90_130), .B (n_84_133), .C1 (n_80_135), .C2 (n_77_135) );
AOI211_X1 g_96_127 (.ZN (n_96_127), .A (n_92_129), .B (n_86_132), .C1 (n_82_134), .C2 (n_76_137) );
AOI211_X1 g_98_126 (.ZN (n_98_126), .A (n_94_128), .B (n_88_131), .C1 (n_84_133), .C2 (n_78_136) );
AOI211_X1 g_100_125 (.ZN (n_100_125), .A (n_96_127), .B (n_90_130), .C1 (n_86_132), .C2 (n_80_135) );
AOI211_X1 g_102_124 (.ZN (n_102_124), .A (n_98_126), .B (n_92_129), .C1 (n_88_131), .C2 (n_82_134) );
AOI211_X1 g_104_123 (.ZN (n_104_123), .A (n_100_125), .B (n_94_128), .C1 (n_90_130), .C2 (n_84_133) );
AOI211_X1 g_106_124 (.ZN (n_106_124), .A (n_102_124), .B (n_96_127), .C1 (n_92_129), .C2 (n_86_132) );
AOI211_X1 g_104_125 (.ZN (n_104_125), .A (n_104_123), .B (n_98_126), .C1 (n_94_128), .C2 (n_88_131) );
AOI211_X1 g_102_126 (.ZN (n_102_126), .A (n_106_124), .B (n_100_125), .C1 (n_96_127), .C2 (n_90_130) );
AOI211_X1 g_103_124 (.ZN (n_103_124), .A (n_104_125), .B (n_102_124), .C1 (n_98_126), .C2 (n_92_129) );
AOI211_X1 g_101_125 (.ZN (n_101_125), .A (n_102_126), .B (n_104_123), .C1 (n_100_125), .C2 (n_94_128) );
AOI211_X1 g_99_126 (.ZN (n_99_126), .A (n_103_124), .B (n_106_124), .C1 (n_102_124), .C2 (n_96_127) );
AOI211_X1 g_97_127 (.ZN (n_97_127), .A (n_101_125), .B (n_104_125), .C1 (n_104_123), .C2 (n_98_126) );
AOI211_X1 g_95_128 (.ZN (n_95_128), .A (n_99_126), .B (n_102_126), .C1 (n_106_124), .C2 (n_100_125) );
AOI211_X1 g_93_129 (.ZN (n_93_129), .A (n_97_127), .B (n_103_124), .C1 (n_104_125), .C2 (n_102_124) );
AOI211_X1 g_91_130 (.ZN (n_91_130), .A (n_95_128), .B (n_101_125), .C1 (n_102_126), .C2 (n_104_123) );
AOI211_X1 g_89_131 (.ZN (n_89_131), .A (n_93_129), .B (n_99_126), .C1 (n_103_124), .C2 (n_106_124) );
AOI211_X1 g_87_132 (.ZN (n_87_132), .A (n_91_130), .B (n_97_127), .C1 (n_101_125), .C2 (n_104_125) );
AOI211_X1 g_85_133 (.ZN (n_85_133), .A (n_89_131), .B (n_95_128), .C1 (n_99_126), .C2 (n_102_126) );
AOI211_X1 g_83_134 (.ZN (n_83_134), .A (n_87_132), .B (n_93_129), .C1 (n_97_127), .C2 (n_103_124) );
AOI211_X1 g_81_135 (.ZN (n_81_135), .A (n_85_133), .B (n_91_130), .C1 (n_95_128), .C2 (n_101_125) );
AOI211_X1 g_79_136 (.ZN (n_79_136), .A (n_83_134), .B (n_89_131), .C1 (n_93_129), .C2 (n_99_126) );
AOI211_X1 g_77_137 (.ZN (n_77_137), .A (n_81_135), .B (n_87_132), .C1 (n_91_130), .C2 (n_97_127) );
AOI211_X1 g_75_138 (.ZN (n_75_138), .A (n_79_136), .B (n_85_133), .C1 (n_89_131), .C2 (n_95_128) );
AOI211_X1 g_76_136 (.ZN (n_76_136), .A (n_77_137), .B (n_83_134), .C1 (n_87_132), .C2 (n_93_129) );
AOI211_X1 g_74_137 (.ZN (n_74_137), .A (n_75_138), .B (n_81_135), .C1 (n_85_133), .C2 (n_91_130) );
AOI211_X1 g_72_138 (.ZN (n_72_138), .A (n_76_136), .B (n_79_136), .C1 (n_83_134), .C2 (n_89_131) );
AOI211_X1 g_70_139 (.ZN (n_70_139), .A (n_74_137), .B (n_77_137), .C1 (n_81_135), .C2 (n_87_132) );
AOI211_X1 g_68_140 (.ZN (n_68_140), .A (n_72_138), .B (n_75_138), .C1 (n_79_136), .C2 (n_85_133) );
AOI211_X1 g_66_141 (.ZN (n_66_141), .A (n_70_139), .B (n_76_136), .C1 (n_77_137), .C2 (n_83_134) );
AOI211_X1 g_64_142 (.ZN (n_64_142), .A (n_68_140), .B (n_74_137), .C1 (n_75_138), .C2 (n_81_135) );
AOI211_X1 g_63_140 (.ZN (n_63_140), .A (n_66_141), .B (n_72_138), .C1 (n_76_136), .C2 (n_79_136) );
AOI211_X1 g_61_139 (.ZN (n_61_139), .A (n_64_142), .B (n_70_139), .C1 (n_74_137), .C2 (n_77_137) );
AOI211_X1 g_62_141 (.ZN (n_62_141), .A (n_63_140), .B (n_68_140), .C1 (n_72_138), .C2 (n_75_138) );
AOI211_X1 g_60_142 (.ZN (n_60_142), .A (n_61_139), .B (n_66_141), .C1 (n_70_139), .C2 (n_76_136) );
AOI211_X1 g_59_140 (.ZN (n_59_140), .A (n_62_141), .B (n_64_142), .C1 (n_68_140), .C2 (n_74_137) );
AOI211_X1 g_57_141 (.ZN (n_57_141), .A (n_60_142), .B (n_63_140), .C1 (n_66_141), .C2 (n_72_138) );
AOI211_X1 g_55_142 (.ZN (n_55_142), .A (n_59_140), .B (n_61_139), .C1 (n_64_142), .C2 (n_70_139) );
AOI211_X1 g_53_143 (.ZN (n_53_143), .A (n_57_141), .B (n_62_141), .C1 (n_63_140), .C2 (n_68_140) );
AOI211_X1 g_51_144 (.ZN (n_51_144), .A (n_55_142), .B (n_60_142), .C1 (n_61_139), .C2 (n_66_141) );
AOI211_X1 g_53_145 (.ZN (n_53_145), .A (n_53_143), .B (n_59_140), .C1 (n_62_141), .C2 (n_64_142) );
AOI211_X1 g_52_143 (.ZN (n_52_143), .A (n_51_144), .B (n_57_141), .C1 (n_60_142), .C2 (n_63_140) );
AOI211_X1 g_50_144 (.ZN (n_50_144), .A (n_53_145), .B (n_55_142), .C1 (n_59_140), .C2 (n_61_139) );
AOI211_X1 g_51_146 (.ZN (n_51_146), .A (n_52_143), .B (n_53_143), .C1 (n_57_141), .C2 (n_62_141) );
AOI211_X1 g_52_144 (.ZN (n_52_144), .A (n_50_144), .B (n_51_144), .C1 (n_55_142), .C2 (n_60_142) );
AOI211_X1 g_50_145 (.ZN (n_50_145), .A (n_51_146), .B (n_53_145), .C1 (n_53_143), .C2 (n_59_140) );
AOI211_X1 g_51_143 (.ZN (n_51_143), .A (n_52_144), .B (n_52_143), .C1 (n_51_144), .C2 (n_57_141) );
AOI211_X1 g_49_144 (.ZN (n_49_144), .A (n_50_145), .B (n_50_144), .C1 (n_53_145), .C2 (n_55_142) );
AOI211_X1 g_47_145 (.ZN (n_47_145), .A (n_51_143), .B (n_51_146), .C1 (n_52_143), .C2 (n_53_143) );
AOI211_X1 g_48_147 (.ZN (n_48_147), .A (n_49_144), .B (n_52_144), .C1 (n_50_144), .C2 (n_51_144) );
AOI211_X1 g_50_146 (.ZN (n_50_146), .A (n_47_145), .B (n_50_145), .C1 (n_51_146), .C2 (n_53_145) );
AOI211_X1 g_51_148 (.ZN (n_51_148), .A (n_48_147), .B (n_51_143), .C1 (n_52_144), .C2 (n_52_143) );
AOI211_X1 g_52_146 (.ZN (n_52_146), .A (n_50_146), .B (n_49_144), .C1 (n_50_145), .C2 (n_50_144) );
AOI211_X1 g_53_144 (.ZN (n_53_144), .A (n_51_148), .B (n_47_145), .C1 (n_51_143), .C2 (n_51_146) );
AOI211_X1 g_51_145 (.ZN (n_51_145), .A (n_52_146), .B (n_48_147), .C1 (n_49_144), .C2 (n_52_144) );
AOI211_X1 g_49_146 (.ZN (n_49_146), .A (n_53_144), .B (n_50_146), .C1 (n_47_145), .C2 (n_50_145) );
AOI211_X1 g_50_148 (.ZN (n_50_148), .A (n_51_145), .B (n_51_148), .C1 (n_48_147), .C2 (n_51_143) );
AOI211_X1 g_52_147 (.ZN (n_52_147), .A (n_49_146), .B (n_52_146), .C1 (n_50_146), .C2 (n_49_144) );
AOI211_X1 g_54_146 (.ZN (n_54_146), .A (n_50_148), .B (n_53_144), .C1 (n_51_148), .C2 (n_47_145) );
AOI211_X1 g_52_145 (.ZN (n_52_145), .A (n_52_147), .B (n_51_145), .C1 (n_52_146), .C2 (n_48_147) );
AOI211_X1 g_51_147 (.ZN (n_51_147), .A (n_54_146), .B (n_49_146), .C1 (n_53_144), .C2 (n_50_146) );
AOI211_X1 g_53_148 (.ZN (n_53_148), .A (n_52_145), .B (n_50_148), .C1 (n_51_145), .C2 (n_51_148) );
AOI211_X1 g_54_150 (.ZN (n_54_150), .A (n_51_147), .B (n_52_147), .C1 (n_49_146), .C2 (n_52_146) );
AOI211_X1 g_52_149 (.ZN (n_52_149), .A (n_53_148), .B (n_54_146), .C1 (n_50_148), .C2 (n_53_144) );
AOI211_X1 g_53_147 (.ZN (n_53_147), .A (n_54_150), .B (n_52_145), .C1 (n_52_147), .C2 (n_51_145) );
AOI211_X1 g_55_148 (.ZN (n_55_148), .A (n_52_149), .B (n_51_147), .C1 (n_54_146), .C2 (n_49_146) );
AOI211_X1 g_56_146 (.ZN (n_56_146), .A (n_53_147), .B (n_53_148), .C1 (n_52_145), .C2 (n_50_148) );
AOI211_X1 g_54_145 (.ZN (n_54_145), .A (n_55_148), .B (n_54_150), .C1 (n_51_147), .C2 (n_52_147) );
AOI211_X1 g_56_144 (.ZN (n_56_144), .A (n_56_146), .B (n_52_149), .C1 (n_53_148), .C2 (n_54_146) );
AOI211_X1 g_58_143 (.ZN (n_58_143), .A (n_54_145), .B (n_53_147), .C1 (n_54_150), .C2 (n_52_145) );
AOI211_X1 g_57_145 (.ZN (n_57_145), .A (n_56_144), .B (n_55_148), .C1 (n_52_149), .C2 (n_51_147) );
AOI211_X1 g_55_146 (.ZN (n_55_146), .A (n_58_143), .B (n_56_146), .C1 (n_53_147), .C2 (n_53_148) );
AOI211_X1 g_54_144 (.ZN (n_54_144), .A (n_57_145), .B (n_54_145), .C1 (n_55_148), .C2 (n_54_150) );
AOI211_X1 g_56_143 (.ZN (n_56_143), .A (n_55_146), .B (n_56_144), .C1 (n_56_146), .C2 (n_52_149) );
AOI211_X1 g_58_142 (.ZN (n_58_142), .A (n_54_144), .B (n_58_143), .C1 (n_54_145), .C2 (n_53_147) );
AOI211_X1 g_60_141 (.ZN (n_60_141), .A (n_56_143), .B (n_57_145), .C1 (n_56_144), .C2 (n_55_148) );
AOI211_X1 g_62_140 (.ZN (n_62_140), .A (n_58_142), .B (n_55_146), .C1 (n_58_143), .C2 (n_56_146) );
AOI211_X1 g_61_142 (.ZN (n_61_142), .A (n_60_141), .B (n_54_144), .C1 (n_57_145), .C2 (n_54_145) );
AOI211_X1 g_59_143 (.ZN (n_59_143), .A (n_62_140), .B (n_56_143), .C1 (n_55_146), .C2 (n_56_144) );
AOI211_X1 g_57_144 (.ZN (n_57_144), .A (n_61_142), .B (n_58_142), .C1 (n_54_144), .C2 (n_58_143) );
AOI211_X1 g_55_145 (.ZN (n_55_145), .A (n_59_143), .B (n_60_141), .C1 (n_56_143), .C2 (n_57_145) );
AOI211_X1 g_53_146 (.ZN (n_53_146), .A (n_57_144), .B (n_62_140), .C1 (n_58_142), .C2 (n_55_146) );
AOI211_X1 g_54_148 (.ZN (n_54_148), .A (n_55_145), .B (n_61_142), .C1 (n_60_141), .C2 (n_54_144) );
AOI211_X1 g_56_147 (.ZN (n_56_147), .A (n_53_146), .B (n_59_143), .C1 (n_62_140), .C2 (n_56_143) );
AOI211_X1 g_58_148 (.ZN (n_58_148), .A (n_54_148), .B (n_57_144), .C1 (n_61_142), .C2 (n_58_142) );
AOI211_X1 g_56_149 (.ZN (n_56_149), .A (n_56_147), .B (n_55_145), .C1 (n_59_143), .C2 (n_60_141) );
AOI211_X1 g_55_147 (.ZN (n_55_147), .A (n_58_148), .B (n_53_146), .C1 (n_57_144), .C2 (n_62_140) );
AOI211_X1 g_57_146 (.ZN (n_57_146), .A (n_56_149), .B (n_54_148), .C1 (n_55_145), .C2 (n_61_142) );
AOI211_X1 g_59_145 (.ZN (n_59_145), .A (n_55_147), .B (n_56_147), .C1 (n_53_146), .C2 (n_59_143) );
AOI211_X1 g_60_147 (.ZN (n_60_147), .A (n_57_146), .B (n_58_148), .C1 (n_54_148), .C2 (n_57_144) );
AOI211_X1 g_58_146 (.ZN (n_58_146), .A (n_59_145), .B (n_56_149), .C1 (n_56_147), .C2 (n_55_145) );
AOI211_X1 g_57_148 (.ZN (n_57_148), .A (n_60_147), .B (n_55_147), .C1 (n_58_148), .C2 (n_53_146) );
AOI211_X1 g_58_150 (.ZN (n_58_150), .A (n_58_146), .B (n_57_146), .C1 (n_56_149), .C2 (n_54_148) );
AOI211_X1 g_59_148 (.ZN (n_59_148), .A (n_57_148), .B (n_59_145), .C1 (n_55_147), .C2 (n_56_147) );
AOI211_X1 g_57_147 (.ZN (n_57_147), .A (n_58_150), .B (n_60_147), .C1 (n_57_146), .C2 (n_58_148) );
AOI211_X1 g_56_145 (.ZN (n_56_145), .A (n_59_148), .B (n_58_146), .C1 (n_59_145), .C2 (n_56_149) );
AOI211_X1 g_57_143 (.ZN (n_57_143), .A (n_57_147), .B (n_57_148), .C1 (n_60_147), .C2 (n_55_147) );
AOI211_X1 g_58_145 (.ZN (n_58_145), .A (n_56_145), .B (n_58_150), .C1 (n_58_146), .C2 (n_57_146) );
AOI211_X1 g_59_147 (.ZN (n_59_147), .A (n_57_143), .B (n_59_148), .C1 (n_57_148), .C2 (n_59_145) );
AOI211_X1 g_60_149 (.ZN (n_60_149), .A (n_58_145), .B (n_57_147), .C1 (n_58_150), .C2 (n_60_147) );
AOI211_X1 g_62_150 (.ZN (n_62_150), .A (n_59_147), .B (n_56_145), .C1 (n_59_148), .C2 (n_58_146) );
AOI211_X1 g_61_148 (.ZN (n_61_148), .A (n_60_149), .B (n_57_143), .C1 (n_57_147), .C2 (n_57_148) );
AOI211_X1 g_60_146 (.ZN (n_60_146), .A (n_62_150), .B (n_58_145), .C1 (n_56_145), .C2 (n_58_150) );
AOI211_X1 g_59_144 (.ZN (n_59_144), .A (n_61_148), .B (n_59_147), .C1 (n_57_143), .C2 (n_59_148) );
AOI211_X1 g_61_143 (.ZN (n_61_143), .A (n_60_146), .B (n_60_149), .C1 (n_58_145), .C2 (n_57_147) );
AOI211_X1 g_59_142 (.ZN (n_59_142), .A (n_59_144), .B (n_62_150), .C1 (n_59_147), .C2 (n_56_145) );
AOI211_X1 g_61_141 (.ZN (n_61_141), .A (n_61_143), .B (n_61_148), .C1 (n_60_149), .C2 (n_57_143) );
AOI211_X1 g_63_142 (.ZN (n_63_142), .A (n_59_142), .B (n_60_146), .C1 (n_62_150), .C2 (n_58_145) );
AOI211_X1 g_62_144 (.ZN (n_62_144), .A (n_61_141), .B (n_59_144), .C1 (n_61_148), .C2 (n_59_147) );
AOI211_X1 g_60_143 (.ZN (n_60_143), .A (n_63_142), .B (n_61_143), .C1 (n_60_146), .C2 (n_60_149) );
AOI211_X1 g_58_144 (.ZN (n_58_144), .A (n_62_144), .B (n_59_142), .C1 (n_59_144), .C2 (n_62_150) );
AOI211_X1 g_60_145 (.ZN (n_60_145), .A (n_60_143), .B (n_61_141), .C1 (n_61_143), .C2 (n_61_148) );
AOI211_X1 g_61_147 (.ZN (n_61_147), .A (n_58_144), .B (n_63_142), .C1 (n_59_142), .C2 (n_60_146) );
AOI211_X1 g_59_146 (.ZN (n_59_146), .A (n_60_145), .B (n_62_144), .C1 (n_61_141), .C2 (n_59_144) );
AOI211_X1 g_61_145 (.ZN (n_61_145), .A (n_61_147), .B (n_60_143), .C1 (n_63_142), .C2 (n_61_143) );
AOI211_X1 g_62_143 (.ZN (n_62_143), .A (n_59_146), .B (n_58_144), .C1 (n_62_144), .C2 (n_59_142) );
AOI211_X1 g_60_144 (.ZN (n_60_144), .A (n_61_145), .B (n_60_145), .C1 (n_60_143), .C2 (n_61_141) );
AOI211_X1 g_61_146 (.ZN (n_61_146), .A (n_62_143), .B (n_61_147), .C1 (n_58_144), .C2 (n_63_142) );
AOI211_X1 g_62_148 (.ZN (n_62_148), .A (n_60_144), .B (n_59_146), .C1 (n_60_145), .C2 (n_62_144) );
AOI211_X1 g_63_146 (.ZN (n_63_146), .A (n_61_146), .B (n_61_145), .C1 (n_61_147), .C2 (n_60_143) );
AOI211_X1 g_64_144 (.ZN (n_64_144), .A (n_62_148), .B (n_62_143), .C1 (n_59_146), .C2 (n_58_144) );
AOI211_X1 g_62_145 (.ZN (n_62_145), .A (n_63_146), .B (n_60_144), .C1 (n_61_145), .C2 (n_60_145) );
AOI211_X1 g_63_147 (.ZN (n_63_147), .A (n_64_144), .B (n_61_146), .C1 (n_62_143), .C2 (n_61_147) );
AOI211_X1 g_64_149 (.ZN (n_64_149), .A (n_62_145), .B (n_62_148), .C1 (n_60_144), .C2 (n_59_146) );
AOI211_X1 g_66_150 (.ZN (n_66_150), .A (n_63_147), .B (n_63_146), .C1 (n_61_146), .C2 (n_61_145) );
AOI211_X1 g_65_148 (.ZN (n_65_148), .A (n_64_149), .B (n_64_144), .C1 (n_62_148), .C2 (n_62_143) );
AOI211_X1 g_64_146 (.ZN (n_64_146), .A (n_66_150), .B (n_62_145), .C1 (n_63_146), .C2 (n_60_144) );
AOI211_X1 g_63_148 (.ZN (n_63_148), .A (n_65_148), .B (n_63_147), .C1 (n_64_144), .C2 (n_61_146) );
AOI211_X1 g_65_147 (.ZN (n_65_147), .A (n_64_146), .B (n_64_149), .C1 (n_62_145), .C2 (n_62_148) );
AOI211_X1 g_67_148 (.ZN (n_67_148), .A (n_63_148), .B (n_66_150), .C1 (n_63_147), .C2 (n_63_146) );
AOI211_X1 g_68_146 (.ZN (n_68_146), .A (n_65_147), .B (n_65_148), .C1 (n_64_149), .C2 (n_64_144) );
AOI211_X1 g_66_145 (.ZN (n_66_145), .A (n_67_148), .B (n_64_146), .C1 (n_66_150), .C2 (n_62_145) );
AOI211_X1 g_65_143 (.ZN (n_65_143), .A (n_68_146), .B (n_63_148), .C1 (n_65_148), .C2 (n_63_147) );
AOI211_X1 g_63_144 (.ZN (n_63_144), .A (n_66_145), .B (n_65_147), .C1 (n_64_146), .C2 (n_64_149) );
AOI211_X1 g_62_142 (.ZN (n_62_142), .A (n_65_143), .B (n_67_148), .C1 (n_63_148), .C2 (n_66_150) );
AOI211_X1 g_64_141 (.ZN (n_64_141), .A (n_63_144), .B (n_68_146), .C1 (n_65_147), .C2 (n_65_148) );
AOI211_X1 g_66_140 (.ZN (n_66_140), .A (n_62_142), .B (n_66_145), .C1 (n_67_148), .C2 (n_64_146) );
AOI211_X1 g_68_139 (.ZN (n_68_139), .A (n_64_141), .B (n_65_143), .C1 (n_68_146), .C2 (n_63_148) );
AOI211_X1 g_67_141 (.ZN (n_67_141), .A (n_66_140), .B (n_63_144), .C1 (n_66_145), .C2 (n_65_147) );
AOI211_X1 g_65_142 (.ZN (n_65_142), .A (n_68_139), .B (n_62_142), .C1 (n_65_143), .C2 (n_67_148) );
AOI211_X1 g_63_143 (.ZN (n_63_143), .A (n_67_141), .B (n_64_141), .C1 (n_63_144), .C2 (n_68_146) );
AOI211_X1 g_61_144 (.ZN (n_61_144), .A (n_65_142), .B (n_66_140), .C1 (n_62_142), .C2 (n_66_145) );
AOI211_X1 g_62_146 (.ZN (n_62_146), .A (n_63_143), .B (n_68_139), .C1 (n_64_141), .C2 (n_65_143) );
AOI211_X1 g_64_145 (.ZN (n_64_145), .A (n_61_144), .B (n_67_141), .C1 (n_66_140), .C2 (n_63_144) );
AOI211_X1 g_66_146 (.ZN (n_66_146), .A (n_62_146), .B (n_65_142), .C1 (n_68_139), .C2 (n_62_142) );
AOI211_X1 g_64_147 (.ZN (n_64_147), .A (n_64_145), .B (n_63_143), .C1 (n_67_141), .C2 (n_64_141) );
AOI211_X1 g_63_145 (.ZN (n_63_145), .A (n_66_146), .B (n_61_144), .C1 (n_65_142), .C2 (n_66_140) );
AOI211_X1 g_65_144 (.ZN (n_65_144), .A (n_64_147), .B (n_62_146), .C1 (n_63_143), .C2 (n_68_139) );
AOI211_X1 g_67_143 (.ZN (n_67_143), .A (n_63_145), .B (n_64_145), .C1 (n_61_144), .C2 (n_67_141) );
AOI211_X1 g_68_141 (.ZN (n_68_141), .A (n_65_144), .B (n_66_146), .C1 (n_62_146), .C2 (n_65_142) );
AOI211_X1 g_66_142 (.ZN (n_66_142), .A (n_67_143), .B (n_64_147), .C1 (n_64_145), .C2 (n_63_143) );
AOI211_X1 g_64_143 (.ZN (n_64_143), .A (n_68_141), .B (n_63_145), .C1 (n_66_146), .C2 (n_61_144) );
AOI211_X1 g_65_145 (.ZN (n_65_145), .A (n_66_142), .B (n_65_144), .C1 (n_64_147), .C2 (n_62_146) );
AOI211_X1 g_67_144 (.ZN (n_67_144), .A (n_64_143), .B (n_67_143), .C1 (n_63_145), .C2 (n_64_145) );
AOI211_X1 g_68_142 (.ZN (n_68_142), .A (n_65_145), .B (n_68_141), .C1 (n_65_144), .C2 (n_66_146) );
AOI211_X1 g_66_143 (.ZN (n_66_143), .A (n_67_144), .B (n_66_142), .C1 (n_67_143), .C2 (n_64_147) );
AOI211_X1 g_67_145 (.ZN (n_67_145), .A (n_68_142), .B (n_64_143), .C1 (n_68_141), .C2 (n_63_145) );
AOI211_X1 g_65_146 (.ZN (n_65_146), .A (n_66_143), .B (n_65_145), .C1 (n_66_142), .C2 (n_65_144) );
AOI211_X1 g_66_148 (.ZN (n_66_148), .A (n_67_145), .B (n_67_144), .C1 (n_64_143), .C2 (n_67_143) );
AOI211_X1 g_68_147 (.ZN (n_68_147), .A (n_65_146), .B (n_68_142), .C1 (n_65_145), .C2 (n_68_141) );
AOI211_X1 g_69_145 (.ZN (n_69_145), .A (n_66_148), .B (n_66_143), .C1 (n_67_144), .C2 (n_66_142) );
AOI211_X1 g_67_146 (.ZN (n_67_146), .A (n_68_147), .B (n_67_145), .C1 (n_68_142), .C2 (n_64_143) );
AOI211_X1 g_66_144 (.ZN (n_66_144), .A (n_69_145), .B (n_65_146), .C1 (n_66_143), .C2 (n_65_145) );
AOI211_X1 g_68_143 (.ZN (n_68_143), .A (n_67_146), .B (n_66_148), .C1 (n_67_145), .C2 (n_67_144) );
AOI211_X1 g_69_141 (.ZN (n_69_141), .A (n_66_144), .B (n_68_147), .C1 (n_65_146), .C2 (n_68_142) );
AOI211_X1 g_67_142 (.ZN (n_67_142), .A (n_68_143), .B (n_69_145), .C1 (n_66_148), .C2 (n_66_143) );
AOI211_X1 g_68_144 (.ZN (n_68_144), .A (n_69_141), .B (n_67_146), .C1 (n_68_147), .C2 (n_67_145) );
AOI211_X1 g_70_143 (.ZN (n_70_143), .A (n_67_142), .B (n_66_144), .C1 (n_69_145), .C2 (n_65_146) );
AOI211_X1 g_71_141 (.ZN (n_71_141), .A (n_68_144), .B (n_68_143), .C1 (n_67_146), .C2 (n_66_148) );
AOI211_X1 g_69_140 (.ZN (n_69_140), .A (n_70_143), .B (n_69_141), .C1 (n_66_144), .C2 (n_68_147) );
AOI211_X1 g_71_139 (.ZN (n_71_139), .A (n_71_141), .B (n_67_142), .C1 (n_68_143), .C2 (n_69_145) );
AOI211_X1 g_73_138 (.ZN (n_73_138), .A (n_69_140), .B (n_68_144), .C1 (n_69_141), .C2 (n_67_146) );
AOI211_X1 g_75_137 (.ZN (n_75_137), .A (n_71_139), .B (n_70_143), .C1 (n_67_142), .C2 (n_66_144) );
AOI211_X1 g_77_136 (.ZN (n_77_136), .A (n_73_138), .B (n_71_141), .C1 (n_68_144), .C2 (n_68_143) );
AOI211_X1 g_79_135 (.ZN (n_79_135), .A (n_75_137), .B (n_69_140), .C1 (n_70_143), .C2 (n_69_141) );
AOI211_X1 g_81_134 (.ZN (n_81_134), .A (n_77_136), .B (n_71_139), .C1 (n_71_141), .C2 (n_67_142) );
AOI211_X1 g_80_136 (.ZN (n_80_136), .A (n_79_135), .B (n_73_138), .C1 (n_69_140), .C2 (n_68_144) );
AOI211_X1 g_82_135 (.ZN (n_82_135), .A (n_81_134), .B (n_75_137), .C1 (n_71_139), .C2 (n_70_143) );
AOI211_X1 g_84_134 (.ZN (n_84_134), .A (n_80_136), .B (n_77_136), .C1 (n_73_138), .C2 (n_71_141) );
AOI211_X1 g_86_133 (.ZN (n_86_133), .A (n_82_135), .B (n_79_135), .C1 (n_75_137), .C2 (n_69_140) );
AOI211_X1 g_88_132 (.ZN (n_88_132), .A (n_84_134), .B (n_81_134), .C1 (n_77_136), .C2 (n_71_139) );
AOI211_X1 g_90_131 (.ZN (n_90_131), .A (n_86_133), .B (n_80_136), .C1 (n_79_135), .C2 (n_73_138) );
AOI211_X1 g_92_130 (.ZN (n_92_130), .A (n_88_132), .B (n_82_135), .C1 (n_81_134), .C2 (n_75_137) );
AOI211_X1 g_94_129 (.ZN (n_94_129), .A (n_90_131), .B (n_84_134), .C1 (n_80_136), .C2 (n_77_136) );
AOI211_X1 g_96_128 (.ZN (n_96_128), .A (n_92_130), .B (n_86_133), .C1 (n_82_135), .C2 (n_79_135) );
AOI211_X1 g_98_127 (.ZN (n_98_127), .A (n_94_129), .B (n_88_132), .C1 (n_84_134), .C2 (n_81_134) );
AOI211_X1 g_100_126 (.ZN (n_100_126), .A (n_96_128), .B (n_90_131), .C1 (n_86_133), .C2 (n_80_136) );
AOI211_X1 g_99_128 (.ZN (n_99_128), .A (n_98_127), .B (n_92_130), .C1 (n_88_132), .C2 (n_82_135) );
AOI211_X1 g_101_127 (.ZN (n_101_127), .A (n_100_126), .B (n_94_129), .C1 (n_90_131), .C2 (n_84_134) );
AOI211_X1 g_103_126 (.ZN (n_103_126), .A (n_99_128), .B (n_96_128), .C1 (n_92_130), .C2 (n_86_133) );
AOI211_X1 g_105_125 (.ZN (n_105_125), .A (n_101_127), .B (n_98_127), .C1 (n_94_129), .C2 (n_88_132) );
AOI211_X1 g_107_124 (.ZN (n_107_124), .A (n_103_126), .B (n_100_126), .C1 (n_96_128), .C2 (n_90_131) );
AOI211_X1 g_109_123 (.ZN (n_109_123), .A (n_105_125), .B (n_99_128), .C1 (n_98_127), .C2 (n_92_130) );
AOI211_X1 g_111_122 (.ZN (n_111_122), .A (n_107_124), .B (n_101_127), .C1 (n_100_126), .C2 (n_94_129) );
AOI211_X1 g_113_121 (.ZN (n_113_121), .A (n_109_123), .B (n_103_126), .C1 (n_99_128), .C2 (n_96_128) );
AOI211_X1 g_115_120 (.ZN (n_115_120), .A (n_111_122), .B (n_105_125), .C1 (n_101_127), .C2 (n_98_127) );
AOI211_X1 g_117_119 (.ZN (n_117_119), .A (n_113_121), .B (n_107_124), .C1 (n_103_126), .C2 (n_100_126) );
AOI211_X1 g_119_118 (.ZN (n_119_118), .A (n_115_120), .B (n_109_123), .C1 (n_105_125), .C2 (n_99_128) );
AOI211_X1 g_118_120 (.ZN (n_118_120), .A (n_117_119), .B (n_111_122), .C1 (n_107_124), .C2 (n_101_127) );
AOI211_X1 g_116_121 (.ZN (n_116_121), .A (n_119_118), .B (n_113_121), .C1 (n_109_123), .C2 (n_103_126) );
AOI211_X1 g_115_119 (.ZN (n_115_119), .A (n_118_120), .B (n_115_120), .C1 (n_111_122), .C2 (n_105_125) );
AOI211_X1 g_113_120 (.ZN (n_113_120), .A (n_116_121), .B (n_117_119), .C1 (n_113_121), .C2 (n_107_124) );
AOI211_X1 g_111_121 (.ZN (n_111_121), .A (n_115_119), .B (n_119_118), .C1 (n_115_120), .C2 (n_109_123) );
AOI211_X1 g_109_122 (.ZN (n_109_122), .A (n_113_120), .B (n_118_120), .C1 (n_117_119), .C2 (n_111_122) );
AOI211_X1 g_107_123 (.ZN (n_107_123), .A (n_111_121), .B (n_116_121), .C1 (n_119_118), .C2 (n_113_121) );
AOI211_X1 g_105_124 (.ZN (n_105_124), .A (n_109_122), .B (n_115_119), .C1 (n_118_120), .C2 (n_115_120) );
AOI211_X1 g_103_125 (.ZN (n_103_125), .A (n_107_123), .B (n_113_120), .C1 (n_116_121), .C2 (n_117_119) );
AOI211_X1 g_101_126 (.ZN (n_101_126), .A (n_105_124), .B (n_111_121), .C1 (n_115_119), .C2 (n_119_118) );
AOI211_X1 g_99_127 (.ZN (n_99_127), .A (n_103_125), .B (n_109_122), .C1 (n_113_120), .C2 (n_118_120) );
AOI211_X1 g_97_128 (.ZN (n_97_128), .A (n_101_126), .B (n_107_123), .C1 (n_111_121), .C2 (n_116_121) );
AOI211_X1 g_95_129 (.ZN (n_95_129), .A (n_99_127), .B (n_105_124), .C1 (n_109_122), .C2 (n_115_119) );
AOI211_X1 g_93_130 (.ZN (n_93_130), .A (n_97_128), .B (n_103_125), .C1 (n_107_123), .C2 (n_113_120) );
AOI211_X1 g_91_131 (.ZN (n_91_131), .A (n_95_129), .B (n_101_126), .C1 (n_105_124), .C2 (n_111_121) );
AOI211_X1 g_89_132 (.ZN (n_89_132), .A (n_93_130), .B (n_99_127), .C1 (n_103_125), .C2 (n_109_122) );
AOI211_X1 g_87_133 (.ZN (n_87_133), .A (n_91_131), .B (n_97_128), .C1 (n_101_126), .C2 (n_107_123) );
AOI211_X1 g_85_134 (.ZN (n_85_134), .A (n_89_132), .B (n_95_129), .C1 (n_99_127), .C2 (n_105_124) );
AOI211_X1 g_83_135 (.ZN (n_83_135), .A (n_87_133), .B (n_93_130), .C1 (n_97_128), .C2 (n_103_125) );
AOI211_X1 g_81_136 (.ZN (n_81_136), .A (n_85_134), .B (n_91_131), .C1 (n_95_129), .C2 (n_101_126) );
AOI211_X1 g_79_137 (.ZN (n_79_137), .A (n_83_135), .B (n_89_132), .C1 (n_93_130), .C2 (n_99_127) );
AOI211_X1 g_77_138 (.ZN (n_77_138), .A (n_81_136), .B (n_87_133), .C1 (n_91_131), .C2 (n_97_128) );
AOI211_X1 g_75_139 (.ZN (n_75_139), .A (n_79_137), .B (n_85_134), .C1 (n_89_132), .C2 (n_95_129) );
AOI211_X1 g_73_140 (.ZN (n_73_140), .A (n_77_138), .B (n_83_135), .C1 (n_87_133), .C2 (n_93_130) );
AOI211_X1 g_74_138 (.ZN (n_74_138), .A (n_75_139), .B (n_81_136), .C1 (n_85_134), .C2 (n_91_131) );
AOI211_X1 g_72_139 (.ZN (n_72_139), .A (n_73_140), .B (n_79_137), .C1 (n_83_135), .C2 (n_89_132) );
AOI211_X1 g_70_140 (.ZN (n_70_140), .A (n_74_138), .B (n_77_138), .C1 (n_81_136), .C2 (n_87_133) );
AOI211_X1 g_69_142 (.ZN (n_69_142), .A (n_72_139), .B (n_75_139), .C1 (n_79_137), .C2 (n_85_134) );
AOI211_X1 g_70_144 (.ZN (n_70_144), .A (n_70_140), .B (n_73_140), .C1 (n_77_138), .C2 (n_83_135) );
AOI211_X1 g_68_145 (.ZN (n_68_145), .A (n_69_142), .B (n_74_138), .C1 (n_75_139), .C2 (n_81_136) );
AOI211_X1 g_67_147 (.ZN (n_67_147), .A (n_70_144), .B (n_72_139), .C1 (n_73_140), .C2 (n_79_137) );
AOI211_X1 g_69_146 (.ZN (n_69_146), .A (n_68_145), .B (n_70_140), .C1 (n_74_138), .C2 (n_77_138) );
AOI211_X1 g_70_148 (.ZN (n_70_148), .A (n_67_147), .B (n_69_142), .C1 (n_72_139), .C2 (n_75_139) );
AOI211_X1 g_68_149 (.ZN (n_68_149), .A (n_69_146), .B (n_70_144), .C1 (n_70_140), .C2 (n_73_140) );
AOI211_X1 g_69_147 (.ZN (n_69_147), .A (n_70_148), .B (n_68_145), .C1 (n_69_142), .C2 (n_74_138) );
AOI211_X1 g_71_146 (.ZN (n_71_146), .A (n_68_149), .B (n_67_147), .C1 (n_70_144), .C2 (n_72_139) );
AOI211_X1 g_73_145 (.ZN (n_73_145), .A (n_69_147), .B (n_69_146), .C1 (n_68_145), .C2 (n_70_140) );
AOI211_X1 g_72_147 (.ZN (n_72_147), .A (n_71_146), .B (n_70_148), .C1 (n_67_147), .C2 (n_69_142) );
AOI211_X1 g_71_145 (.ZN (n_71_145), .A (n_73_145), .B (n_68_149), .C1 (n_69_146), .C2 (n_70_144) );
AOI211_X1 g_69_144 (.ZN (n_69_144), .A (n_72_147), .B (n_69_147), .C1 (n_70_148), .C2 (n_68_145) );
AOI211_X1 g_70_142 (.ZN (n_70_142), .A (n_71_145), .B (n_71_146), .C1 (n_68_149), .C2 (n_67_147) );
AOI211_X1 g_71_140 (.ZN (n_71_140), .A (n_69_144), .B (n_73_145), .C1 (n_69_147), .C2 (n_69_146) );
AOI211_X1 g_73_139 (.ZN (n_73_139), .A (n_70_142), .B (n_72_147), .C1 (n_71_146), .C2 (n_70_148) );
AOI211_X1 g_72_141 (.ZN (n_72_141), .A (n_71_140), .B (n_71_145), .C1 (n_73_145), .C2 (n_68_149) );
AOI211_X1 g_74_140 (.ZN (n_74_140), .A (n_73_139), .B (n_69_144), .C1 (n_72_147), .C2 (n_69_147) );
AOI211_X1 g_76_139 (.ZN (n_76_139), .A (n_72_141), .B (n_70_142), .C1 (n_71_145), .C2 (n_71_146) );
AOI211_X1 g_78_138 (.ZN (n_78_138), .A (n_74_140), .B (n_71_140), .C1 (n_69_144), .C2 (n_73_145) );
AOI211_X1 g_80_137 (.ZN (n_80_137), .A (n_76_139), .B (n_73_139), .C1 (n_70_142), .C2 (n_72_147) );
AOI211_X1 g_82_136 (.ZN (n_82_136), .A (n_78_138), .B (n_72_141), .C1 (n_71_140), .C2 (n_71_145) );
AOI211_X1 g_84_135 (.ZN (n_84_135), .A (n_80_137), .B (n_74_140), .C1 (n_73_139), .C2 (n_69_144) );
AOI211_X1 g_86_134 (.ZN (n_86_134), .A (n_82_136), .B (n_76_139), .C1 (n_72_141), .C2 (n_70_142) );
AOI211_X1 g_88_133 (.ZN (n_88_133), .A (n_84_135), .B (n_78_138), .C1 (n_74_140), .C2 (n_71_140) );
AOI211_X1 g_90_132 (.ZN (n_90_132), .A (n_86_134), .B (n_80_137), .C1 (n_76_139), .C2 (n_73_139) );
AOI211_X1 g_92_131 (.ZN (n_92_131), .A (n_88_133), .B (n_82_136), .C1 (n_78_138), .C2 (n_72_141) );
AOI211_X1 g_94_130 (.ZN (n_94_130), .A (n_90_132), .B (n_84_135), .C1 (n_80_137), .C2 (n_74_140) );
AOI211_X1 g_96_129 (.ZN (n_96_129), .A (n_92_131), .B (n_86_134), .C1 (n_82_136), .C2 (n_76_139) );
AOI211_X1 g_98_128 (.ZN (n_98_128), .A (n_94_130), .B (n_88_133), .C1 (n_84_135), .C2 (n_78_138) );
AOI211_X1 g_100_127 (.ZN (n_100_127), .A (n_96_129), .B (n_90_132), .C1 (n_86_134), .C2 (n_80_137) );
AOI211_X1 g_99_129 (.ZN (n_99_129), .A (n_98_128), .B (n_92_131), .C1 (n_88_133), .C2 (n_82_136) );
AOI211_X1 g_101_128 (.ZN (n_101_128), .A (n_100_127), .B (n_94_130), .C1 (n_90_132), .C2 (n_84_135) );
AOI211_X1 g_103_127 (.ZN (n_103_127), .A (n_99_129), .B (n_96_129), .C1 (n_92_131), .C2 (n_86_134) );
AOI211_X1 g_105_126 (.ZN (n_105_126), .A (n_101_128), .B (n_98_128), .C1 (n_94_130), .C2 (n_88_133) );
AOI211_X1 g_107_125 (.ZN (n_107_125), .A (n_103_127), .B (n_100_127), .C1 (n_96_129), .C2 (n_90_132) );
AOI211_X1 g_106_127 (.ZN (n_106_127), .A (n_105_126), .B (n_99_129), .C1 (n_98_128), .C2 (n_92_131) );
AOI211_X1 g_104_126 (.ZN (n_104_126), .A (n_107_125), .B (n_101_128), .C1 (n_100_127), .C2 (n_94_130) );
AOI211_X1 g_106_125 (.ZN (n_106_125), .A (n_106_127), .B (n_103_127), .C1 (n_99_129), .C2 (n_96_129) );
AOI211_X1 g_108_124 (.ZN (n_108_124), .A (n_104_126), .B (n_105_126), .C1 (n_101_128), .C2 (n_98_128) );
AOI211_X1 g_110_123 (.ZN (n_110_123), .A (n_106_125), .B (n_107_125), .C1 (n_103_127), .C2 (n_100_127) );
AOI211_X1 g_112_122 (.ZN (n_112_122), .A (n_108_124), .B (n_106_127), .C1 (n_105_126), .C2 (n_99_129) );
AOI211_X1 g_114_121 (.ZN (n_114_121), .A (n_110_123), .B (n_104_126), .C1 (n_107_125), .C2 (n_101_128) );
AOI211_X1 g_116_120 (.ZN (n_116_120), .A (n_112_122), .B (n_106_125), .C1 (n_106_127), .C2 (n_103_127) );
AOI211_X1 g_115_122 (.ZN (n_115_122), .A (n_114_121), .B (n_108_124), .C1 (n_104_126), .C2 (n_105_126) );
AOI211_X1 g_117_121 (.ZN (n_117_121), .A (n_116_120), .B (n_110_123), .C1 (n_106_125), .C2 (n_107_125) );
AOI211_X1 g_119_120 (.ZN (n_119_120), .A (n_115_122), .B (n_112_122), .C1 (n_108_124), .C2 (n_106_127) );
AOI211_X1 g_121_119 (.ZN (n_121_119), .A (n_117_121), .B (n_114_121), .C1 (n_110_123), .C2 (n_104_126) );
AOI211_X1 g_120_121 (.ZN (n_120_121), .A (n_119_120), .B (n_116_120), .C1 (n_112_122), .C2 (n_106_125) );
AOI211_X1 g_122_120 (.ZN (n_122_120), .A (n_121_119), .B (n_115_122), .C1 (n_114_121), .C2 (n_108_124) );
AOI211_X1 g_124_119 (.ZN (n_124_119), .A (n_120_121), .B (n_117_121), .C1 (n_116_120), .C2 (n_110_123) );
AOI211_X1 g_126_118 (.ZN (n_126_118), .A (n_122_120), .B (n_119_120), .C1 (n_115_122), .C2 (n_112_122) );
AOI211_X1 g_128_119 (.ZN (n_128_119), .A (n_124_119), .B (n_121_119), .C1 (n_117_121), .C2 (n_114_121) );
AOI211_X1 g_129_117 (.ZN (n_129_117), .A (n_126_118), .B (n_120_121), .C1 (n_119_120), .C2 (n_116_120) );
AOI211_X1 g_131_116 (.ZN (n_131_116), .A (n_128_119), .B (n_122_120), .C1 (n_121_119), .C2 (n_115_122) );
AOI211_X1 g_133_115 (.ZN (n_133_115), .A (n_129_117), .B (n_124_119), .C1 (n_120_121), .C2 (n_117_121) );
AOI211_X1 g_135_114 (.ZN (n_135_114), .A (n_131_116), .B (n_126_118), .C1 (n_122_120), .C2 (n_119_120) );
AOI211_X1 g_137_113 (.ZN (n_137_113), .A (n_133_115), .B (n_128_119), .C1 (n_124_119), .C2 (n_121_119) );
AOI211_X1 g_139_112 (.ZN (n_139_112), .A (n_135_114), .B (n_129_117), .C1 (n_126_118), .C2 (n_120_121) );
AOI211_X1 g_141_113 (.ZN (n_141_113), .A (n_137_113), .B (n_131_116), .C1 (n_128_119), .C2 (n_122_120) );
AOI211_X1 g_143_114 (.ZN (n_143_114), .A (n_139_112), .B (n_133_115), .C1 (n_129_117), .C2 (n_124_119) );
AOI211_X1 g_144_116 (.ZN (n_144_116), .A (n_141_113), .B (n_135_114), .C1 (n_131_116), .C2 (n_126_118) );
AOI211_X1 g_142_115 (.ZN (n_142_115), .A (n_143_114), .B (n_137_113), .C1 (n_133_115), .C2 (n_128_119) );
AOI211_X1 g_140_116 (.ZN (n_140_116), .A (n_144_116), .B (n_139_112), .C1 (n_135_114), .C2 (n_129_117) );
AOI211_X1 g_139_114 (.ZN (n_139_114), .A (n_142_115), .B (n_141_113), .C1 (n_137_113), .C2 (n_131_116) );
AOI211_X1 g_137_115 (.ZN (n_137_115), .A (n_140_116), .B (n_143_114), .C1 (n_139_112), .C2 (n_133_115) );
AOI211_X1 g_135_116 (.ZN (n_135_116), .A (n_139_114), .B (n_144_116), .C1 (n_141_113), .C2 (n_135_114) );
AOI211_X1 g_133_117 (.ZN (n_133_117), .A (n_137_115), .B (n_142_115), .C1 (n_143_114), .C2 (n_137_113) );
AOI211_X1 g_131_118 (.ZN (n_131_118), .A (n_135_116), .B (n_140_116), .C1 (n_144_116), .C2 (n_139_112) );
AOI211_X1 g_129_119 (.ZN (n_129_119), .A (n_133_117), .B (n_139_114), .C1 (n_142_115), .C2 (n_141_113) );
AOI211_X1 g_130_117 (.ZN (n_130_117), .A (n_131_118), .B (n_137_115), .C1 (n_140_116), .C2 (n_143_114) );
AOI211_X1 g_128_118 (.ZN (n_128_118), .A (n_129_119), .B (n_135_116), .C1 (n_139_114), .C2 (n_144_116) );
AOI211_X1 g_126_117 (.ZN (n_126_117), .A (n_130_117), .B (n_133_117), .C1 (n_137_115), .C2 (n_142_115) );
AOI211_X1 g_124_118 (.ZN (n_124_118), .A (n_128_118), .B (n_131_118), .C1 (n_135_116), .C2 (n_140_116) );
AOI211_X1 g_122_119 (.ZN (n_122_119), .A (n_126_117), .B (n_129_119), .C1 (n_133_117), .C2 (n_139_114) );
AOI211_X1 g_120_120 (.ZN (n_120_120), .A (n_124_118), .B (n_130_117), .C1 (n_131_118), .C2 (n_137_115) );
AOI211_X1 g_118_121 (.ZN (n_118_121), .A (n_122_119), .B (n_128_118), .C1 (n_129_119), .C2 (n_135_116) );
AOI211_X1 g_116_122 (.ZN (n_116_122), .A (n_120_120), .B (n_126_117), .C1 (n_130_117), .C2 (n_133_117) );
AOI211_X1 g_117_120 (.ZN (n_117_120), .A (n_118_121), .B (n_124_118), .C1 (n_128_118), .C2 (n_131_118) );
AOI211_X1 g_115_121 (.ZN (n_115_121), .A (n_116_122), .B (n_122_119), .C1 (n_126_117), .C2 (n_129_119) );
AOI211_X1 g_113_122 (.ZN (n_113_122), .A (n_117_120), .B (n_120_120), .C1 (n_124_118), .C2 (n_130_117) );
AOI211_X1 g_111_123 (.ZN (n_111_123), .A (n_115_121), .B (n_118_121), .C1 (n_122_119), .C2 (n_128_118) );
AOI211_X1 g_110_125 (.ZN (n_110_125), .A (n_113_122), .B (n_116_122), .C1 (n_120_120), .C2 (n_126_117) );
AOI211_X1 g_108_126 (.ZN (n_108_126), .A (n_111_123), .B (n_117_120), .C1 (n_118_121), .C2 (n_124_118) );
AOI211_X1 g_107_128 (.ZN (n_107_128), .A (n_110_125), .B (n_115_121), .C1 (n_116_122), .C2 (n_122_119) );
AOI211_X1 g_106_126 (.ZN (n_106_126), .A (n_108_126), .B (n_113_122), .C1 (n_117_120), .C2 (n_120_120) );
AOI211_X1 g_108_125 (.ZN (n_108_125), .A (n_107_128), .B (n_111_123), .C1 (n_115_121), .C2 (n_118_121) );
AOI211_X1 g_110_124 (.ZN (n_110_124), .A (n_106_126), .B (n_110_125), .C1 (n_113_122), .C2 (n_116_122) );
AOI211_X1 g_112_123 (.ZN (n_112_123), .A (n_108_125), .B (n_108_126), .C1 (n_111_123), .C2 (n_117_120) );
AOI211_X1 g_114_122 (.ZN (n_114_122), .A (n_110_124), .B (n_107_128), .C1 (n_110_125), .C2 (n_115_121) );
AOI211_X1 g_113_124 (.ZN (n_113_124), .A (n_112_123), .B (n_106_126), .C1 (n_108_126), .C2 (n_113_122) );
AOI211_X1 g_115_123 (.ZN (n_115_123), .A (n_114_122), .B (n_108_125), .C1 (n_107_128), .C2 (n_111_123) );
AOI211_X1 g_117_122 (.ZN (n_117_122), .A (n_113_124), .B (n_110_124), .C1 (n_106_126), .C2 (n_110_125) );
AOI211_X1 g_119_121 (.ZN (n_119_121), .A (n_115_123), .B (n_112_123), .C1 (n_108_125), .C2 (n_108_126) );
AOI211_X1 g_121_120 (.ZN (n_121_120), .A (n_117_122), .B (n_114_122), .C1 (n_110_124), .C2 (n_107_128) );
AOI211_X1 g_123_119 (.ZN (n_123_119), .A (n_119_121), .B (n_113_124), .C1 (n_112_123), .C2 (n_106_126) );
AOI211_X1 g_125_118 (.ZN (n_125_118), .A (n_121_120), .B (n_115_123), .C1 (n_114_122), .C2 (n_108_125) );
AOI211_X1 g_124_120 (.ZN (n_124_120), .A (n_123_119), .B (n_117_122), .C1 (n_113_124), .C2 (n_110_124) );
AOI211_X1 g_126_119 (.ZN (n_126_119), .A (n_125_118), .B (n_119_121), .C1 (n_115_123), .C2 (n_112_123) );
AOI211_X1 g_125_121 (.ZN (n_125_121), .A (n_124_120), .B (n_121_120), .C1 (n_117_122), .C2 (n_114_122) );
AOI211_X1 g_127_120 (.ZN (n_127_120), .A (n_126_119), .B (n_123_119), .C1 (n_119_121), .C2 (n_113_124) );
AOI211_X1 g_125_119 (.ZN (n_125_119), .A (n_125_121), .B (n_125_118), .C1 (n_121_120), .C2 (n_115_123) );
AOI211_X1 g_127_118 (.ZN (n_127_118), .A (n_127_120), .B (n_124_120), .C1 (n_123_119), .C2 (n_117_122) );
AOI211_X1 g_126_120 (.ZN (n_126_120), .A (n_125_119), .B (n_126_119), .C1 (n_125_118), .C2 (n_119_121) );
AOI211_X1 g_124_121 (.ZN (n_124_121), .A (n_127_118), .B (n_125_121), .C1 (n_124_120), .C2 (n_121_120) );
AOI211_X1 g_122_122 (.ZN (n_122_122), .A (n_126_120), .B (n_127_120), .C1 (n_126_119), .C2 (n_123_119) );
AOI211_X1 g_123_120 (.ZN (n_123_120), .A (n_124_121), .B (n_125_119), .C1 (n_125_121), .C2 (n_125_118) );
AOI211_X1 g_121_121 (.ZN (n_121_121), .A (n_122_122), .B (n_127_118), .C1 (n_127_120), .C2 (n_124_120) );
AOI211_X1 g_119_122 (.ZN (n_119_122), .A (n_123_120), .B (n_126_120), .C1 (n_125_119), .C2 (n_126_119) );
AOI211_X1 g_117_123 (.ZN (n_117_123), .A (n_121_121), .B (n_124_121), .C1 (n_127_118), .C2 (n_125_121) );
AOI211_X1 g_115_124 (.ZN (n_115_124), .A (n_119_122), .B (n_122_122), .C1 (n_126_120), .C2 (n_127_120) );
AOI211_X1 g_113_123 (.ZN (n_113_123), .A (n_117_123), .B (n_123_120), .C1 (n_124_121), .C2 (n_125_119) );
AOI211_X1 g_111_124 (.ZN (n_111_124), .A (n_115_124), .B (n_121_121), .C1 (n_122_122), .C2 (n_127_118) );
AOI211_X1 g_109_125 (.ZN (n_109_125), .A (n_113_123), .B (n_119_122), .C1 (n_123_120), .C2 (n_126_120) );
AOI211_X1 g_107_126 (.ZN (n_107_126), .A (n_111_124), .B (n_117_123), .C1 (n_121_121), .C2 (n_124_121) );
AOI211_X1 g_105_127 (.ZN (n_105_127), .A (n_109_125), .B (n_115_124), .C1 (n_119_122), .C2 (n_122_122) );
AOI211_X1 g_103_128 (.ZN (n_103_128), .A (n_107_126), .B (n_113_123), .C1 (n_117_123), .C2 (n_123_120) );
AOI211_X1 g_101_129 (.ZN (n_101_129), .A (n_105_127), .B (n_111_124), .C1 (n_115_124), .C2 (n_121_121) );
AOI211_X1 g_102_127 (.ZN (n_102_127), .A (n_103_128), .B (n_109_125), .C1 (n_113_123), .C2 (n_119_122) );
AOI211_X1 g_100_128 (.ZN (n_100_128), .A (n_101_129), .B (n_107_126), .C1 (n_111_124), .C2 (n_117_123) );
AOI211_X1 g_98_129 (.ZN (n_98_129), .A (n_102_127), .B (n_105_127), .C1 (n_109_125), .C2 (n_115_124) );
AOI211_X1 g_96_130 (.ZN (n_96_130), .A (n_100_128), .B (n_103_128), .C1 (n_107_126), .C2 (n_113_123) );
AOI211_X1 g_94_131 (.ZN (n_94_131), .A (n_98_129), .B (n_101_129), .C1 (n_105_127), .C2 (n_111_124) );
AOI211_X1 g_92_132 (.ZN (n_92_132), .A (n_96_130), .B (n_102_127), .C1 (n_103_128), .C2 (n_109_125) );
AOI211_X1 g_90_133 (.ZN (n_90_133), .A (n_94_131), .B (n_100_128), .C1 (n_101_129), .C2 (n_107_126) );
AOI211_X1 g_88_134 (.ZN (n_88_134), .A (n_92_132), .B (n_98_129), .C1 (n_102_127), .C2 (n_105_127) );
AOI211_X1 g_86_135 (.ZN (n_86_135), .A (n_90_133), .B (n_96_130), .C1 (n_100_128), .C2 (n_103_128) );
AOI211_X1 g_84_136 (.ZN (n_84_136), .A (n_88_134), .B (n_94_131), .C1 (n_98_129), .C2 (n_101_129) );
AOI211_X1 g_82_137 (.ZN (n_82_137), .A (n_86_135), .B (n_92_132), .C1 (n_96_130), .C2 (n_102_127) );
AOI211_X1 g_80_138 (.ZN (n_80_138), .A (n_84_136), .B (n_90_133), .C1 (n_94_131), .C2 (n_100_128) );
AOI211_X1 g_78_137 (.ZN (n_78_137), .A (n_82_137), .B (n_88_134), .C1 (n_92_132), .C2 (n_98_129) );
AOI211_X1 g_76_138 (.ZN (n_76_138), .A (n_80_138), .B (n_86_135), .C1 (n_90_133), .C2 (n_96_130) );
AOI211_X1 g_74_139 (.ZN (n_74_139), .A (n_78_137), .B (n_84_136), .C1 (n_88_134), .C2 (n_94_131) );
AOI211_X1 g_72_140 (.ZN (n_72_140), .A (n_76_138), .B (n_82_137), .C1 (n_86_135), .C2 (n_92_132) );
AOI211_X1 g_70_141 (.ZN (n_70_141), .A (n_74_139), .B (n_80_138), .C1 (n_84_136), .C2 (n_90_133) );
AOI211_X1 g_69_143 (.ZN (n_69_143), .A (n_72_140), .B (n_78_137), .C1 (n_82_137), .C2 (n_88_134) );
AOI211_X1 g_71_142 (.ZN (n_71_142), .A (n_70_141), .B (n_76_138), .C1 (n_80_138), .C2 (n_86_135) );
AOI211_X1 g_73_141 (.ZN (n_73_141), .A (n_69_143), .B (n_74_139), .C1 (n_78_137), .C2 (n_84_136) );
AOI211_X1 g_72_143 (.ZN (n_72_143), .A (n_71_142), .B (n_72_140), .C1 (n_76_138), .C2 (n_82_137) );
AOI211_X1 g_74_142 (.ZN (n_74_142), .A (n_73_141), .B (n_70_141), .C1 (n_74_139), .C2 (n_80_138) );
AOI211_X1 g_75_140 (.ZN (n_75_140), .A (n_72_143), .B (n_69_143), .C1 (n_72_140), .C2 (n_78_137) );
AOI211_X1 g_77_139 (.ZN (n_77_139), .A (n_74_142), .B (n_71_142), .C1 (n_70_141), .C2 (n_76_138) );
AOI211_X1 g_79_138 (.ZN (n_79_138), .A (n_75_140), .B (n_73_141), .C1 (n_69_143), .C2 (n_74_139) );
AOI211_X1 g_81_137 (.ZN (n_81_137), .A (n_77_139), .B (n_72_143), .C1 (n_71_142), .C2 (n_72_140) );
AOI211_X1 g_83_136 (.ZN (n_83_136), .A (n_79_138), .B (n_74_142), .C1 (n_73_141), .C2 (n_70_141) );
AOI211_X1 g_85_135 (.ZN (n_85_135), .A (n_81_137), .B (n_75_140), .C1 (n_72_143), .C2 (n_69_143) );
AOI211_X1 g_87_134 (.ZN (n_87_134), .A (n_83_136), .B (n_77_139), .C1 (n_74_142), .C2 (n_71_142) );
AOI211_X1 g_89_133 (.ZN (n_89_133), .A (n_85_135), .B (n_79_138), .C1 (n_75_140), .C2 (n_73_141) );
AOI211_X1 g_91_132 (.ZN (n_91_132), .A (n_87_134), .B (n_81_137), .C1 (n_77_139), .C2 (n_72_143) );
AOI211_X1 g_93_131 (.ZN (n_93_131), .A (n_89_133), .B (n_83_136), .C1 (n_79_138), .C2 (n_74_142) );
AOI211_X1 g_95_130 (.ZN (n_95_130), .A (n_91_132), .B (n_85_135), .C1 (n_81_137), .C2 (n_75_140) );
AOI211_X1 g_97_129 (.ZN (n_97_129), .A (n_93_131), .B (n_87_134), .C1 (n_83_136), .C2 (n_77_139) );
AOI211_X1 g_99_130 (.ZN (n_99_130), .A (n_95_130), .B (n_89_133), .C1 (n_85_135), .C2 (n_79_138) );
AOI211_X1 g_97_131 (.ZN (n_97_131), .A (n_97_129), .B (n_91_132), .C1 (n_87_134), .C2 (n_81_137) );
AOI211_X1 g_95_132 (.ZN (n_95_132), .A (n_99_130), .B (n_93_131), .C1 (n_89_133), .C2 (n_83_136) );
AOI211_X1 g_93_133 (.ZN (n_93_133), .A (n_97_131), .B (n_95_130), .C1 (n_91_132), .C2 (n_85_135) );
AOI211_X1 g_91_134 (.ZN (n_91_134), .A (n_95_132), .B (n_97_129), .C1 (n_93_131), .C2 (n_87_134) );
AOI211_X1 g_89_135 (.ZN (n_89_135), .A (n_93_133), .B (n_99_130), .C1 (n_95_130), .C2 (n_89_133) );
AOI211_X1 g_87_136 (.ZN (n_87_136), .A (n_91_134), .B (n_97_131), .C1 (n_97_129), .C2 (n_91_132) );
AOI211_X1 g_85_137 (.ZN (n_85_137), .A (n_89_135), .B (n_95_132), .C1 (n_99_130), .C2 (n_93_131) );
AOI211_X1 g_83_138 (.ZN (n_83_138), .A (n_87_136), .B (n_93_133), .C1 (n_97_131), .C2 (n_95_130) );
AOI211_X1 g_81_139 (.ZN (n_81_139), .A (n_85_137), .B (n_91_134), .C1 (n_95_132), .C2 (n_97_129) );
AOI211_X1 g_79_140 (.ZN (n_79_140), .A (n_83_138), .B (n_89_135), .C1 (n_93_133), .C2 (n_99_130) );
AOI211_X1 g_77_141 (.ZN (n_77_141), .A (n_81_139), .B (n_87_136), .C1 (n_91_134), .C2 (n_97_131) );
AOI211_X1 g_78_139 (.ZN (n_78_139), .A (n_79_140), .B (n_85_137), .C1 (n_89_135), .C2 (n_95_132) );
AOI211_X1 g_76_140 (.ZN (n_76_140), .A (n_77_141), .B (n_83_138), .C1 (n_87_136), .C2 (n_93_133) );
AOI211_X1 g_74_141 (.ZN (n_74_141), .A (n_78_139), .B (n_81_139), .C1 (n_85_137), .C2 (n_91_134) );
AOI211_X1 g_72_142 (.ZN (n_72_142), .A (n_76_140), .B (n_79_140), .C1 (n_83_138), .C2 (n_89_135) );
AOI211_X1 g_71_144 (.ZN (n_71_144), .A (n_74_141), .B (n_77_141), .C1 (n_81_139), .C2 (n_87_136) );
AOI211_X1 g_70_146 (.ZN (n_70_146), .A (n_72_142), .B (n_78_139), .C1 (n_79_140), .C2 (n_85_137) );
AOI211_X1 g_69_148 (.ZN (n_69_148), .A (n_71_144), .B (n_76_140), .C1 (n_77_141), .C2 (n_83_138) );
AOI211_X1 g_70_150 (.ZN (n_70_150), .A (n_70_146), .B (n_74_141), .C1 (n_78_139), .C2 (n_81_139) );
AOI211_X1 g_71_148 (.ZN (n_71_148), .A (n_69_148), .B (n_72_142), .C1 (n_76_140), .C2 (n_79_140) );
AOI211_X1 g_72_146 (.ZN (n_72_146), .A (n_70_150), .B (n_71_144), .C1 (n_74_141), .C2 (n_77_141) );
AOI211_X1 g_70_145 (.ZN (n_70_145), .A (n_71_148), .B (n_70_146), .C1 (n_72_142), .C2 (n_78_139) );
AOI211_X1 g_71_143 (.ZN (n_71_143), .A (n_72_146), .B (n_69_148), .C1 (n_71_144), .C2 (n_76_140) );
AOI211_X1 g_73_144 (.ZN (n_73_144), .A (n_70_145), .B (n_70_150), .C1 (n_70_146), .C2 (n_74_141) );
AOI211_X1 g_75_143 (.ZN (n_75_143), .A (n_71_143), .B (n_71_148), .C1 (n_69_148), .C2 (n_72_142) );
AOI211_X1 g_76_141 (.ZN (n_76_141), .A (n_73_144), .B (n_72_146), .C1 (n_70_150), .C2 (n_71_144) );
AOI211_X1 g_78_140 (.ZN (n_78_140), .A (n_75_143), .B (n_70_145), .C1 (n_71_148), .C2 (n_70_146) );
AOI211_X1 g_80_139 (.ZN (n_80_139), .A (n_76_141), .B (n_71_143), .C1 (n_72_146), .C2 (n_69_148) );
AOI211_X1 g_82_138 (.ZN (n_82_138), .A (n_78_140), .B (n_73_144), .C1 (n_70_145), .C2 (n_70_150) );
AOI211_X1 g_84_137 (.ZN (n_84_137), .A (n_80_139), .B (n_75_143), .C1 (n_71_143), .C2 (n_71_148) );
AOI211_X1 g_86_136 (.ZN (n_86_136), .A (n_82_138), .B (n_76_141), .C1 (n_73_144), .C2 (n_72_146) );
AOI211_X1 g_88_135 (.ZN (n_88_135), .A (n_84_137), .B (n_78_140), .C1 (n_75_143), .C2 (n_70_145) );
AOI211_X1 g_90_134 (.ZN (n_90_134), .A (n_86_136), .B (n_80_139), .C1 (n_76_141), .C2 (n_71_143) );
AOI211_X1 g_92_133 (.ZN (n_92_133), .A (n_88_135), .B (n_82_138), .C1 (n_78_140), .C2 (n_73_144) );
AOI211_X1 g_94_132 (.ZN (n_94_132), .A (n_90_134), .B (n_84_137), .C1 (n_80_139), .C2 (n_75_143) );
AOI211_X1 g_96_131 (.ZN (n_96_131), .A (n_92_133), .B (n_86_136), .C1 (n_82_138), .C2 (n_76_141) );
AOI211_X1 g_98_130 (.ZN (n_98_130), .A (n_94_132), .B (n_88_135), .C1 (n_84_137), .C2 (n_78_140) );
AOI211_X1 g_100_129 (.ZN (n_100_129), .A (n_96_131), .B (n_90_134), .C1 (n_86_136), .C2 (n_80_139) );
AOI211_X1 g_102_128 (.ZN (n_102_128), .A (n_98_130), .B (n_92_133), .C1 (n_88_135), .C2 (n_82_138) );
AOI211_X1 g_104_127 (.ZN (n_104_127), .A (n_100_129), .B (n_94_132), .C1 (n_90_134), .C2 (n_84_137) );
AOI211_X1 g_105_129 (.ZN (n_105_129), .A (n_102_128), .B (n_96_131), .C1 (n_92_133), .C2 (n_86_136) );
AOI211_X1 g_103_130 (.ZN (n_103_130), .A (n_104_127), .B (n_98_130), .C1 (n_94_132), .C2 (n_88_135) );
AOI211_X1 g_104_128 (.ZN (n_104_128), .A (n_105_129), .B (n_100_129), .C1 (n_96_131), .C2 (n_90_134) );
AOI211_X1 g_102_129 (.ZN (n_102_129), .A (n_103_130), .B (n_102_128), .C1 (n_98_130), .C2 (n_92_133) );
AOI211_X1 g_100_130 (.ZN (n_100_130), .A (n_104_128), .B (n_104_127), .C1 (n_100_129), .C2 (n_94_132) );
AOI211_X1 g_98_131 (.ZN (n_98_131), .A (n_102_129), .B (n_105_129), .C1 (n_102_128), .C2 (n_96_131) );
AOI211_X1 g_96_132 (.ZN (n_96_132), .A (n_100_130), .B (n_103_130), .C1 (n_104_127), .C2 (n_98_130) );
AOI211_X1 g_97_130 (.ZN (n_97_130), .A (n_98_131), .B (n_104_128), .C1 (n_105_129), .C2 (n_100_129) );
AOI211_X1 g_95_131 (.ZN (n_95_131), .A (n_96_132), .B (n_102_129), .C1 (n_103_130), .C2 (n_102_128) );
AOI211_X1 g_93_132 (.ZN (n_93_132), .A (n_97_130), .B (n_100_130), .C1 (n_104_128), .C2 (n_104_127) );
AOI211_X1 g_91_133 (.ZN (n_91_133), .A (n_95_131), .B (n_98_131), .C1 (n_102_129), .C2 (n_105_129) );
AOI211_X1 g_89_134 (.ZN (n_89_134), .A (n_93_132), .B (n_96_132), .C1 (n_100_130), .C2 (n_103_130) );
AOI211_X1 g_87_135 (.ZN (n_87_135), .A (n_91_133), .B (n_97_130), .C1 (n_98_131), .C2 (n_104_128) );
AOI211_X1 g_85_136 (.ZN (n_85_136), .A (n_89_134), .B (n_95_131), .C1 (n_96_132), .C2 (n_102_129) );
AOI211_X1 g_83_137 (.ZN (n_83_137), .A (n_87_135), .B (n_93_132), .C1 (n_97_130), .C2 (n_100_130) );
AOI211_X1 g_81_138 (.ZN (n_81_138), .A (n_85_136), .B (n_91_133), .C1 (n_95_131), .C2 (n_98_131) );
AOI211_X1 g_79_139 (.ZN (n_79_139), .A (n_83_137), .B (n_89_134), .C1 (n_93_132), .C2 (n_96_132) );
AOI211_X1 g_77_140 (.ZN (n_77_140), .A (n_81_138), .B (n_87_135), .C1 (n_91_133), .C2 (n_97_130) );
AOI211_X1 g_75_141 (.ZN (n_75_141), .A (n_79_139), .B (n_85_136), .C1 (n_89_134), .C2 (n_95_131) );
AOI211_X1 g_73_142 (.ZN (n_73_142), .A (n_77_140), .B (n_83_137), .C1 (n_87_135), .C2 (n_93_132) );
AOI211_X1 g_72_144 (.ZN (n_72_144), .A (n_75_141), .B (n_81_138), .C1 (n_85_136), .C2 (n_91_133) );
AOI211_X1 g_74_143 (.ZN (n_74_143), .A (n_73_142), .B (n_79_139), .C1 (n_83_137), .C2 (n_89_134) );
AOI211_X1 g_76_142 (.ZN (n_76_142), .A (n_72_144), .B (n_77_140), .C1 (n_81_138), .C2 (n_87_135) );
AOI211_X1 g_78_141 (.ZN (n_78_141), .A (n_74_143), .B (n_75_141), .C1 (n_79_139), .C2 (n_85_136) );
AOI211_X1 g_80_140 (.ZN (n_80_140), .A (n_76_142), .B (n_73_142), .C1 (n_77_140), .C2 (n_83_137) );
AOI211_X1 g_82_139 (.ZN (n_82_139), .A (n_78_141), .B (n_72_144), .C1 (n_75_141), .C2 (n_81_138) );
AOI211_X1 g_84_138 (.ZN (n_84_138), .A (n_80_140), .B (n_74_143), .C1 (n_73_142), .C2 (n_79_139) );
AOI211_X1 g_86_137 (.ZN (n_86_137), .A (n_82_139), .B (n_76_142), .C1 (n_72_144), .C2 (n_77_140) );
AOI211_X1 g_88_136 (.ZN (n_88_136), .A (n_84_138), .B (n_78_141), .C1 (n_74_143), .C2 (n_75_141) );
AOI211_X1 g_90_135 (.ZN (n_90_135), .A (n_86_137), .B (n_80_140), .C1 (n_76_142), .C2 (n_73_142) );
AOI211_X1 g_92_134 (.ZN (n_92_134), .A (n_88_136), .B (n_82_139), .C1 (n_78_141), .C2 (n_72_144) );
AOI211_X1 g_94_133 (.ZN (n_94_133), .A (n_90_135), .B (n_84_138), .C1 (n_80_140), .C2 (n_74_143) );
AOI211_X1 g_93_135 (.ZN (n_93_135), .A (n_92_134), .B (n_86_137), .C1 (n_82_139), .C2 (n_76_142) );
AOI211_X1 g_95_134 (.ZN (n_95_134), .A (n_94_133), .B (n_88_136), .C1 (n_84_138), .C2 (n_78_141) );
AOI211_X1 g_97_133 (.ZN (n_97_133), .A (n_93_135), .B (n_90_135), .C1 (n_86_137), .C2 (n_80_140) );
AOI211_X1 g_99_132 (.ZN (n_99_132), .A (n_95_134), .B (n_92_134), .C1 (n_88_136), .C2 (n_82_139) );
AOI211_X1 g_101_131 (.ZN (n_101_131), .A (n_97_133), .B (n_94_133), .C1 (n_90_135), .C2 (n_84_138) );
AOI211_X1 g_100_133 (.ZN (n_100_133), .A (n_99_132), .B (n_93_135), .C1 (n_92_134), .C2 (n_86_137) );
AOI211_X1 g_99_131 (.ZN (n_99_131), .A (n_101_131), .B (n_95_134), .C1 (n_94_133), .C2 (n_88_136) );
AOI211_X1 g_101_130 (.ZN (n_101_130), .A (n_100_133), .B (n_97_133), .C1 (n_93_135), .C2 (n_90_135) );
AOI211_X1 g_103_129 (.ZN (n_103_129), .A (n_99_131), .B (n_99_132), .C1 (n_95_134), .C2 (n_92_134) );
AOI211_X1 g_105_128 (.ZN (n_105_128), .A (n_101_130), .B (n_101_131), .C1 (n_97_133), .C2 (n_94_133) );
AOI211_X1 g_107_127 (.ZN (n_107_127), .A (n_103_129), .B (n_100_133), .C1 (n_99_132), .C2 (n_93_135) );
AOI211_X1 g_109_126 (.ZN (n_109_126), .A (n_105_128), .B (n_99_131), .C1 (n_101_131), .C2 (n_95_134) );
AOI211_X1 g_111_125 (.ZN (n_111_125), .A (n_107_127), .B (n_101_130), .C1 (n_100_133), .C2 (n_97_133) );
AOI211_X1 g_110_127 (.ZN (n_110_127), .A (n_109_126), .B (n_103_129), .C1 (n_99_131), .C2 (n_99_132) );
AOI211_X1 g_112_126 (.ZN (n_112_126), .A (n_111_125), .B (n_105_128), .C1 (n_101_130), .C2 (n_101_131) );
AOI211_X1 g_114_125 (.ZN (n_114_125), .A (n_110_127), .B (n_107_127), .C1 (n_103_129), .C2 (n_100_133) );
AOI211_X1 g_112_124 (.ZN (n_112_124), .A (n_112_126), .B (n_109_126), .C1 (n_105_128), .C2 (n_99_131) );
AOI211_X1 g_114_123 (.ZN (n_114_123), .A (n_114_125), .B (n_111_125), .C1 (n_107_127), .C2 (n_101_130) );
AOI211_X1 g_113_125 (.ZN (n_113_125), .A (n_112_124), .B (n_110_127), .C1 (n_109_126), .C2 (n_103_129) );
AOI211_X1 g_111_126 (.ZN (n_111_126), .A (n_114_123), .B (n_112_126), .C1 (n_111_125), .C2 (n_105_128) );
AOI211_X1 g_109_127 (.ZN (n_109_127), .A (n_113_125), .B (n_114_125), .C1 (n_110_127), .C2 (n_107_127) );
AOI211_X1 g_108_129 (.ZN (n_108_129), .A (n_111_126), .B (n_112_124), .C1 (n_112_126), .C2 (n_109_126) );
AOI211_X1 g_106_128 (.ZN (n_106_128), .A (n_109_127), .B (n_114_123), .C1 (n_114_125), .C2 (n_111_125) );
AOI211_X1 g_108_127 (.ZN (n_108_127), .A (n_108_129), .B (n_113_125), .C1 (n_112_124), .C2 (n_110_127) );
AOI211_X1 g_110_126 (.ZN (n_110_126), .A (n_106_128), .B (n_111_126), .C1 (n_114_123), .C2 (n_112_126) );
AOI211_X1 g_112_125 (.ZN (n_112_125), .A (n_108_127), .B (n_109_127), .C1 (n_113_125), .C2 (n_114_125) );
AOI211_X1 g_114_124 (.ZN (n_114_124), .A (n_110_126), .B (n_108_129), .C1 (n_111_126), .C2 (n_112_124) );
AOI211_X1 g_116_123 (.ZN (n_116_123), .A (n_112_125), .B (n_106_128), .C1 (n_109_127), .C2 (n_114_123) );
AOI211_X1 g_118_122 (.ZN (n_118_122), .A (n_114_124), .B (n_108_127), .C1 (n_108_129), .C2 (n_113_125) );
AOI211_X1 g_120_123 (.ZN (n_120_123), .A (n_116_123), .B (n_110_126), .C1 (n_106_128), .C2 (n_111_126) );
AOI211_X1 g_118_124 (.ZN (n_118_124), .A (n_118_122), .B (n_112_125), .C1 (n_108_127), .C2 (n_109_127) );
AOI211_X1 g_116_125 (.ZN (n_116_125), .A (n_120_123), .B (n_114_124), .C1 (n_110_126), .C2 (n_108_129) );
AOI211_X1 g_114_126 (.ZN (n_114_126), .A (n_118_124), .B (n_116_123), .C1 (n_112_125), .C2 (n_106_128) );
AOI211_X1 g_112_127 (.ZN (n_112_127), .A (n_116_125), .B (n_118_122), .C1 (n_114_124), .C2 (n_108_127) );
AOI211_X1 g_110_128 (.ZN (n_110_128), .A (n_114_126), .B (n_120_123), .C1 (n_116_123), .C2 (n_110_126) );
AOI211_X1 g_109_130 (.ZN (n_109_130), .A (n_112_127), .B (n_118_124), .C1 (n_118_122), .C2 (n_112_125) );
AOI211_X1 g_108_128 (.ZN (n_108_128), .A (n_110_128), .B (n_116_125), .C1 (n_120_123), .C2 (n_114_124) );
AOI211_X1 g_106_129 (.ZN (n_106_129), .A (n_109_130), .B (n_114_126), .C1 (n_118_124), .C2 (n_116_123) );
AOI211_X1 g_104_130 (.ZN (n_104_130), .A (n_108_128), .B (n_112_127), .C1 (n_116_125), .C2 (n_118_122) );
AOI211_X1 g_102_131 (.ZN (n_102_131), .A (n_106_129), .B (n_110_128), .C1 (n_114_126), .C2 (n_120_123) );
AOI211_X1 g_100_132 (.ZN (n_100_132), .A (n_104_130), .B (n_109_130), .C1 (n_112_127), .C2 (n_118_124) );
AOI211_X1 g_98_133 (.ZN (n_98_133), .A (n_102_131), .B (n_108_128), .C1 (n_110_128), .C2 (n_116_125) );
AOI211_X1 g_96_134 (.ZN (n_96_134), .A (n_100_132), .B (n_106_129), .C1 (n_109_130), .C2 (n_114_126) );
AOI211_X1 g_97_132 (.ZN (n_97_132), .A (n_98_133), .B (n_104_130), .C1 (n_108_128), .C2 (n_112_127) );
AOI211_X1 g_95_133 (.ZN (n_95_133), .A (n_96_134), .B (n_102_131), .C1 (n_106_129), .C2 (n_110_128) );
AOI211_X1 g_93_134 (.ZN (n_93_134), .A (n_97_132), .B (n_100_132), .C1 (n_104_130), .C2 (n_109_130) );
AOI211_X1 g_91_135 (.ZN (n_91_135), .A (n_95_133), .B (n_98_133), .C1 (n_102_131), .C2 (n_108_128) );
AOI211_X1 g_89_136 (.ZN (n_89_136), .A (n_93_134), .B (n_96_134), .C1 (n_100_132), .C2 (n_106_129) );
AOI211_X1 g_87_137 (.ZN (n_87_137), .A (n_91_135), .B (n_97_132), .C1 (n_98_133), .C2 (n_104_130) );
AOI211_X1 g_85_138 (.ZN (n_85_138), .A (n_89_136), .B (n_95_133), .C1 (n_96_134), .C2 (n_102_131) );
AOI211_X1 g_83_139 (.ZN (n_83_139), .A (n_87_137), .B (n_93_134), .C1 (n_97_132), .C2 (n_100_132) );
AOI211_X1 g_81_140 (.ZN (n_81_140), .A (n_85_138), .B (n_91_135), .C1 (n_95_133), .C2 (n_98_133) );
AOI211_X1 g_79_141 (.ZN (n_79_141), .A (n_83_139), .B (n_89_136), .C1 (n_93_134), .C2 (n_96_134) );
AOI211_X1 g_77_142 (.ZN (n_77_142), .A (n_81_140), .B (n_87_137), .C1 (n_91_135), .C2 (n_97_132) );
AOI211_X1 g_76_144 (.ZN (n_76_144), .A (n_79_141), .B (n_85_138), .C1 (n_89_136), .C2 (n_95_133) );
AOI211_X1 g_75_142 (.ZN (n_75_142), .A (n_77_142), .B (n_83_139), .C1 (n_87_137), .C2 (n_93_134) );
AOI211_X1 g_73_143 (.ZN (n_73_143), .A (n_76_144), .B (n_81_140), .C1 (n_85_138), .C2 (n_91_135) );
AOI211_X1 g_74_145 (.ZN (n_74_145), .A (n_75_142), .B (n_79_141), .C1 (n_83_139), .C2 (n_89_136) );
AOI211_X1 g_73_147 (.ZN (n_73_147), .A (n_73_143), .B (n_77_142), .C1 (n_81_140), .C2 (n_87_137) );
AOI211_X1 g_72_145 (.ZN (n_72_145), .A (n_74_145), .B (n_76_144), .C1 (n_79_141), .C2 (n_85_138) );
AOI211_X1 g_71_147 (.ZN (n_71_147), .A (n_73_147), .B (n_75_142), .C1 (n_77_142), .C2 (n_83_139) );
AOI211_X1 g_72_149 (.ZN (n_72_149), .A (n_72_145), .B (n_73_143), .C1 (n_76_144), .C2 (n_81_140) );
AOI211_X1 g_74_150 (.ZN (n_74_150), .A (n_71_147), .B (n_74_145), .C1 (n_75_142), .C2 (n_79_141) );
AOI211_X1 g_73_148 (.ZN (n_73_148), .A (n_72_149), .B (n_73_147), .C1 (n_73_143), .C2 (n_77_142) );
AOI211_X1 g_74_146 (.ZN (n_74_146), .A (n_74_150), .B (n_72_145), .C1 (n_74_145), .C2 (n_76_144) );
AOI211_X1 g_75_148 (.ZN (n_75_148), .A (n_73_148), .B (n_71_147), .C1 (n_73_147), .C2 (n_75_142) );
AOI211_X1 g_76_146 (.ZN (n_76_146), .A (n_74_146), .B (n_72_149), .C1 (n_72_145), .C2 (n_73_143) );
AOI211_X1 g_75_144 (.ZN (n_75_144), .A (n_75_148), .B (n_74_150), .C1 (n_71_147), .C2 (n_74_145) );
AOI211_X1 g_77_143 (.ZN (n_77_143), .A (n_76_146), .B (n_73_148), .C1 (n_72_149), .C2 (n_73_147) );
AOI211_X1 g_79_142 (.ZN (n_79_142), .A (n_75_144), .B (n_74_146), .C1 (n_74_150), .C2 (n_72_145) );
AOI211_X1 g_81_141 (.ZN (n_81_141), .A (n_77_143), .B (n_75_148), .C1 (n_73_148), .C2 (n_71_147) );
AOI211_X1 g_83_140 (.ZN (n_83_140), .A (n_79_142), .B (n_76_146), .C1 (n_74_146), .C2 (n_72_149) );
AOI211_X1 g_85_139 (.ZN (n_85_139), .A (n_81_141), .B (n_75_144), .C1 (n_75_148), .C2 (n_74_150) );
AOI211_X1 g_87_138 (.ZN (n_87_138), .A (n_83_140), .B (n_77_143), .C1 (n_76_146), .C2 (n_73_148) );
AOI211_X1 g_89_137 (.ZN (n_89_137), .A (n_85_139), .B (n_79_142), .C1 (n_75_144), .C2 (n_74_146) );
AOI211_X1 g_91_136 (.ZN (n_91_136), .A (n_87_138), .B (n_81_141), .C1 (n_77_143), .C2 (n_75_148) );
AOI211_X1 g_90_138 (.ZN (n_90_138), .A (n_89_137), .B (n_83_140), .C1 (n_79_142), .C2 (n_76_146) );
AOI211_X1 g_88_137 (.ZN (n_88_137), .A (n_91_136), .B (n_85_139), .C1 (n_81_141), .C2 (n_75_144) );
AOI211_X1 g_90_136 (.ZN (n_90_136), .A (n_90_138), .B (n_87_138), .C1 (n_83_140), .C2 (n_77_143) );
AOI211_X1 g_92_135 (.ZN (n_92_135), .A (n_88_137), .B (n_89_137), .C1 (n_85_139), .C2 (n_79_142) );
AOI211_X1 g_94_134 (.ZN (n_94_134), .A (n_90_136), .B (n_91_136), .C1 (n_87_138), .C2 (n_81_141) );
AOI211_X1 g_96_133 (.ZN (n_96_133), .A (n_92_135), .B (n_90_138), .C1 (n_89_137), .C2 (n_83_140) );
AOI211_X1 g_98_132 (.ZN (n_98_132), .A (n_94_134), .B (n_88_137), .C1 (n_91_136), .C2 (n_85_139) );
AOI211_X1 g_100_131 (.ZN (n_100_131), .A (n_96_133), .B (n_90_136), .C1 (n_90_138), .C2 (n_87_138) );
AOI211_X1 g_102_130 (.ZN (n_102_130), .A (n_98_132), .B (n_92_135), .C1 (n_88_137), .C2 (n_89_137) );
AOI211_X1 g_104_129 (.ZN (n_104_129), .A (n_100_131), .B (n_94_134), .C1 (n_90_136), .C2 (n_91_136) );
AOI211_X1 g_106_130 (.ZN (n_106_130), .A (n_102_130), .B (n_96_133), .C1 (n_92_135), .C2 (n_90_138) );
AOI211_X1 g_104_131 (.ZN (n_104_131), .A (n_104_129), .B (n_98_132), .C1 (n_94_134), .C2 (n_88_137) );
AOI211_X1 g_102_132 (.ZN (n_102_132), .A (n_106_130), .B (n_100_131), .C1 (n_96_133), .C2 (n_90_136) );
AOI211_X1 g_101_134 (.ZN (n_101_134), .A (n_104_131), .B (n_102_130), .C1 (n_98_132), .C2 (n_92_135) );
AOI211_X1 g_99_133 (.ZN (n_99_133), .A (n_102_132), .B (n_104_129), .C1 (n_100_131), .C2 (n_94_134) );
AOI211_X1 g_101_132 (.ZN (n_101_132), .A (n_101_134), .B (n_106_130), .C1 (n_102_130), .C2 (n_96_133) );
AOI211_X1 g_103_131 (.ZN (n_103_131), .A (n_99_133), .B (n_104_131), .C1 (n_104_129), .C2 (n_98_132) );
AOI211_X1 g_105_130 (.ZN (n_105_130), .A (n_101_132), .B (n_102_132), .C1 (n_106_130), .C2 (n_100_131) );
AOI211_X1 g_107_129 (.ZN (n_107_129), .A (n_103_131), .B (n_101_134), .C1 (n_104_131), .C2 (n_102_130) );
AOI211_X1 g_109_128 (.ZN (n_109_128), .A (n_105_130), .B (n_99_133), .C1 (n_102_132), .C2 (n_104_129) );
AOI211_X1 g_111_127 (.ZN (n_111_127), .A (n_107_129), .B (n_101_132), .C1 (n_101_134), .C2 (n_106_130) );
AOI211_X1 g_113_126 (.ZN (n_113_126), .A (n_109_128), .B (n_103_131), .C1 (n_99_133), .C2 (n_104_131) );
AOI211_X1 g_115_125 (.ZN (n_115_125), .A (n_111_127), .B (n_105_130), .C1 (n_101_132), .C2 (n_102_132) );
AOI211_X1 g_117_124 (.ZN (n_117_124), .A (n_113_126), .B (n_107_129), .C1 (n_103_131), .C2 (n_101_134) );
AOI211_X1 g_119_123 (.ZN (n_119_123), .A (n_115_125), .B (n_109_128), .C1 (n_105_130), .C2 (n_99_133) );
AOI211_X1 g_121_122 (.ZN (n_121_122), .A (n_117_124), .B (n_111_127), .C1 (n_107_129), .C2 (n_101_132) );
AOI211_X1 g_123_121 (.ZN (n_123_121), .A (n_119_123), .B (n_113_126), .C1 (n_109_128), .C2 (n_103_131) );
AOI211_X1 g_125_120 (.ZN (n_125_120), .A (n_121_122), .B (n_115_125), .C1 (n_111_127), .C2 (n_105_130) );
AOI211_X1 g_127_119 (.ZN (n_127_119), .A (n_123_121), .B (n_117_124), .C1 (n_113_126), .C2 (n_107_129) );
AOI211_X1 g_129_118 (.ZN (n_129_118), .A (n_125_120), .B (n_119_123), .C1 (n_115_125), .C2 (n_109_128) );
AOI211_X1 g_131_117 (.ZN (n_131_117), .A (n_127_119), .B (n_121_122), .C1 (n_117_124), .C2 (n_111_127) );
AOI211_X1 g_133_116 (.ZN (n_133_116), .A (n_129_118), .B (n_123_121), .C1 (n_119_123), .C2 (n_113_126) );
AOI211_X1 g_135_115 (.ZN (n_135_115), .A (n_131_117), .B (n_125_120), .C1 (n_121_122), .C2 (n_115_125) );
AOI211_X1 g_134_117 (.ZN (n_134_117), .A (n_133_116), .B (n_127_119), .C1 (n_123_121), .C2 (n_117_124) );
AOI211_X1 g_136_116 (.ZN (n_136_116), .A (n_135_115), .B (n_129_118), .C1 (n_125_120), .C2 (n_119_123) );
AOI211_X1 g_138_115 (.ZN (n_138_115), .A (n_134_117), .B (n_131_117), .C1 (n_127_119), .C2 (n_121_122) );
AOI211_X1 g_137_117 (.ZN (n_137_117), .A (n_136_116), .B (n_133_116), .C1 (n_129_118), .C2 (n_123_121) );
AOI211_X1 g_136_115 (.ZN (n_136_115), .A (n_138_115), .B (n_135_115), .C1 (n_131_117), .C2 (n_125_120) );
AOI211_X1 g_138_114 (.ZN (n_138_114), .A (n_137_117), .B (n_134_117), .C1 (n_133_116), .C2 (n_127_119) );
AOI211_X1 g_140_113 (.ZN (n_140_113), .A (n_136_115), .B (n_136_116), .C1 (n_135_115), .C2 (n_129_118) );
AOI211_X1 g_139_115 (.ZN (n_139_115), .A (n_138_114), .B (n_138_115), .C1 (n_134_117), .C2 (n_131_117) );
AOI211_X1 g_137_116 (.ZN (n_137_116), .A (n_140_113), .B (n_137_117), .C1 (n_136_116), .C2 (n_133_116) );
AOI211_X1 g_135_117 (.ZN (n_135_117), .A (n_139_115), .B (n_136_115), .C1 (n_138_115), .C2 (n_135_115) );
AOI211_X1 g_133_118 (.ZN (n_133_118), .A (n_137_116), .B (n_138_114), .C1 (n_137_117), .C2 (n_134_117) );
AOI211_X1 g_134_116 (.ZN (n_134_116), .A (n_135_117), .B (n_140_113), .C1 (n_136_115), .C2 (n_136_116) );
AOI211_X1 g_132_117 (.ZN (n_132_117), .A (n_133_118), .B (n_139_115), .C1 (n_138_114), .C2 (n_138_115) );
AOI211_X1 g_130_118 (.ZN (n_130_118), .A (n_134_116), .B (n_137_116), .C1 (n_140_113), .C2 (n_137_117) );
AOI211_X1 g_129_120 (.ZN (n_129_120), .A (n_132_117), .B (n_135_117), .C1 (n_139_115), .C2 (n_136_115) );
AOI211_X1 g_131_119 (.ZN (n_131_119), .A (n_130_118), .B (n_133_118), .C1 (n_137_116), .C2 (n_138_114) );
AOI211_X1 g_130_121 (.ZN (n_130_121), .A (n_129_120), .B (n_134_116), .C1 (n_135_117), .C2 (n_140_113) );
AOI211_X1 g_128_120 (.ZN (n_128_120), .A (n_131_119), .B (n_132_117), .C1 (n_133_118), .C2 (n_139_115) );
AOI211_X1 g_130_119 (.ZN (n_130_119), .A (n_130_121), .B (n_130_118), .C1 (n_134_116), .C2 (n_137_116) );
AOI211_X1 g_132_118 (.ZN (n_132_118), .A (n_128_120), .B (n_129_120), .C1 (n_132_117), .C2 (n_135_117) );
AOI211_X1 g_131_120 (.ZN (n_131_120), .A (n_130_119), .B (n_131_119), .C1 (n_130_118), .C2 (n_133_118) );
AOI211_X1 g_133_119 (.ZN (n_133_119), .A (n_132_118), .B (n_130_121), .C1 (n_129_120), .C2 (n_134_116) );
AOI211_X1 g_135_118 (.ZN (n_135_118), .A (n_131_120), .B (n_128_120), .C1 (n_131_119), .C2 (n_132_117) );
AOI211_X1 g_134_120 (.ZN (n_134_120), .A (n_133_119), .B (n_130_119), .C1 (n_130_121), .C2 (n_130_118) );
AOI211_X1 g_132_119 (.ZN (n_132_119), .A (n_135_118), .B (n_132_118), .C1 (n_128_120), .C2 (n_129_120) );
AOI211_X1 g_134_118 (.ZN (n_134_118), .A (n_134_120), .B (n_131_120), .C1 (n_130_119), .C2 (n_131_119) );
AOI211_X1 g_136_117 (.ZN (n_136_117), .A (n_132_119), .B (n_133_119), .C1 (n_132_118), .C2 (n_130_121) );
AOI211_X1 g_138_116 (.ZN (n_138_116), .A (n_134_118), .B (n_135_118), .C1 (n_131_120), .C2 (n_128_120) );
AOI211_X1 g_140_115 (.ZN (n_140_115), .A (n_136_117), .B (n_134_120), .C1 (n_133_119), .C2 (n_130_119) );
AOI211_X1 g_142_114 (.ZN (n_142_114), .A (n_138_116), .B (n_132_119), .C1 (n_135_118), .C2 (n_132_118) );
AOI211_X1 g_141_116 (.ZN (n_141_116), .A (n_140_115), .B (n_134_118), .C1 (n_134_120), .C2 (n_131_120) );
AOI211_X1 g_139_117 (.ZN (n_139_117), .A (n_142_114), .B (n_136_117), .C1 (n_132_119), .C2 (n_133_119) );
AOI211_X1 g_137_118 (.ZN (n_137_118), .A (n_141_116), .B (n_138_116), .C1 (n_134_118), .C2 (n_135_118) );
AOI211_X1 g_135_119 (.ZN (n_135_119), .A (n_139_117), .B (n_140_115), .C1 (n_136_117), .C2 (n_134_120) );
AOI211_X1 g_133_120 (.ZN (n_133_120), .A (n_137_118), .B (n_142_114), .C1 (n_138_116), .C2 (n_132_119) );
AOI211_X1 g_131_121 (.ZN (n_131_121), .A (n_135_119), .B (n_141_116), .C1 (n_140_115), .C2 (n_134_118) );
AOI211_X1 g_129_122 (.ZN (n_129_122), .A (n_133_120), .B (n_139_117), .C1 (n_142_114), .C2 (n_136_117) );
AOI211_X1 g_130_120 (.ZN (n_130_120), .A (n_131_121), .B (n_137_118), .C1 (n_141_116), .C2 (n_138_116) );
AOI211_X1 g_128_121 (.ZN (n_128_121), .A (n_129_122), .B (n_135_119), .C1 (n_139_117), .C2 (n_140_115) );
AOI211_X1 g_126_122 (.ZN (n_126_122), .A (n_130_120), .B (n_133_120), .C1 (n_137_118), .C2 (n_142_114) );
AOI211_X1 g_124_123 (.ZN (n_124_123), .A (n_128_121), .B (n_131_121), .C1 (n_135_119), .C2 (n_141_116) );
AOI211_X1 g_122_124 (.ZN (n_122_124), .A (n_126_122), .B (n_129_122), .C1 (n_133_120), .C2 (n_139_117) );
AOI211_X1 g_123_122 (.ZN (n_123_122), .A (n_124_123), .B (n_130_120), .C1 (n_131_121), .C2 (n_137_118) );
AOI211_X1 g_121_123 (.ZN (n_121_123), .A (n_122_124), .B (n_128_121), .C1 (n_129_122), .C2 (n_135_119) );
AOI211_X1 g_122_121 (.ZN (n_122_121), .A (n_123_122), .B (n_126_122), .C1 (n_130_120), .C2 (n_133_120) );
AOI211_X1 g_120_122 (.ZN (n_120_122), .A (n_121_123), .B (n_124_123), .C1 (n_128_121), .C2 (n_131_121) );
AOI211_X1 g_118_123 (.ZN (n_118_123), .A (n_122_121), .B (n_122_124), .C1 (n_126_122), .C2 (n_129_122) );
AOI211_X1 g_116_124 (.ZN (n_116_124), .A (n_120_122), .B (n_123_122), .C1 (n_124_123), .C2 (n_130_120) );
AOI211_X1 g_115_126 (.ZN (n_115_126), .A (n_118_123), .B (n_121_123), .C1 (n_122_124), .C2 (n_128_121) );
AOI211_X1 g_117_125 (.ZN (n_117_125), .A (n_116_124), .B (n_122_121), .C1 (n_123_122), .C2 (n_126_122) );
AOI211_X1 g_119_124 (.ZN (n_119_124), .A (n_115_126), .B (n_120_122), .C1 (n_121_123), .C2 (n_124_123) );
AOI211_X1 g_118_126 (.ZN (n_118_126), .A (n_117_125), .B (n_118_123), .C1 (n_122_121), .C2 (n_122_124) );
AOI211_X1 g_120_125 (.ZN (n_120_125), .A (n_119_124), .B (n_116_124), .C1 (n_120_122), .C2 (n_123_122) );
AOI211_X1 g_119_127 (.ZN (n_119_127), .A (n_118_126), .B (n_115_126), .C1 (n_118_123), .C2 (n_121_123) );
AOI211_X1 g_118_125 (.ZN (n_118_125), .A (n_120_125), .B (n_117_125), .C1 (n_116_124), .C2 (n_122_121) );
AOI211_X1 g_120_124 (.ZN (n_120_124), .A (n_119_127), .B (n_119_124), .C1 (n_115_126), .C2 (n_120_122) );
AOI211_X1 g_122_123 (.ZN (n_122_123), .A (n_118_125), .B (n_118_126), .C1 (n_117_125), .C2 (n_118_123) );
AOI211_X1 g_124_122 (.ZN (n_124_122), .A (n_120_124), .B (n_120_125), .C1 (n_119_124), .C2 (n_116_124) );
AOI211_X1 g_126_121 (.ZN (n_126_121), .A (n_122_123), .B (n_119_127), .C1 (n_118_126), .C2 (n_115_126) );
AOI211_X1 g_128_122 (.ZN (n_128_122), .A (n_124_122), .B (n_118_125), .C1 (n_120_125), .C2 (n_117_125) );
AOI211_X1 g_126_123 (.ZN (n_126_123), .A (n_126_121), .B (n_120_124), .C1 (n_119_127), .C2 (n_119_124) );
AOI211_X1 g_127_121 (.ZN (n_127_121), .A (n_128_122), .B (n_122_123), .C1 (n_118_125), .C2 (n_118_126) );
AOI211_X1 g_125_122 (.ZN (n_125_122), .A (n_126_123), .B (n_124_122), .C1 (n_120_124), .C2 (n_120_125) );
AOI211_X1 g_123_123 (.ZN (n_123_123), .A (n_127_121), .B (n_126_121), .C1 (n_122_123), .C2 (n_119_127) );
AOI211_X1 g_121_124 (.ZN (n_121_124), .A (n_125_122), .B (n_128_122), .C1 (n_124_122), .C2 (n_118_125) );
AOI211_X1 g_119_125 (.ZN (n_119_125), .A (n_123_123), .B (n_126_123), .C1 (n_126_121), .C2 (n_120_124) );
AOI211_X1 g_117_126 (.ZN (n_117_126), .A (n_121_124), .B (n_127_121), .C1 (n_128_122), .C2 (n_122_123) );
AOI211_X1 g_115_127 (.ZN (n_115_127), .A (n_119_125), .B (n_125_122), .C1 (n_126_123), .C2 (n_124_122) );
AOI211_X1 g_113_128 (.ZN (n_113_128), .A (n_117_126), .B (n_123_123), .C1 (n_127_121), .C2 (n_126_121) );
AOI211_X1 g_111_129 (.ZN (n_111_129), .A (n_115_127), .B (n_121_124), .C1 (n_125_122), .C2 (n_128_122) );
AOI211_X1 g_110_131 (.ZN (n_110_131), .A (n_113_128), .B (n_119_125), .C1 (n_123_123), .C2 (n_126_123) );
AOI211_X1 g_109_129 (.ZN (n_109_129), .A (n_111_129), .B (n_117_126), .C1 (n_121_124), .C2 (n_127_121) );
AOI211_X1 g_111_128 (.ZN (n_111_128), .A (n_110_131), .B (n_115_127), .C1 (n_119_125), .C2 (n_125_122) );
AOI211_X1 g_113_127 (.ZN (n_113_127), .A (n_109_129), .B (n_113_128), .C1 (n_117_126), .C2 (n_123_123) );
AOI211_X1 g_112_129 (.ZN (n_112_129), .A (n_111_128), .B (n_111_129), .C1 (n_115_127), .C2 (n_121_124) );
AOI211_X1 g_114_128 (.ZN (n_114_128), .A (n_113_127), .B (n_110_131), .C1 (n_113_128), .C2 (n_119_125) );
AOI211_X1 g_116_127 (.ZN (n_116_127), .A (n_112_129), .B (n_109_129), .C1 (n_111_129), .C2 (n_117_126) );
AOI211_X1 g_115_129 (.ZN (n_115_129), .A (n_114_128), .B (n_111_128), .C1 (n_110_131), .C2 (n_115_127) );
AOI211_X1 g_117_128 (.ZN (n_117_128), .A (n_116_127), .B (n_113_127), .C1 (n_109_129), .C2 (n_113_128) );
AOI211_X1 g_116_126 (.ZN (n_116_126), .A (n_115_129), .B (n_112_129), .C1 (n_111_128), .C2 (n_111_129) );
AOI211_X1 g_114_127 (.ZN (n_114_127), .A (n_117_128), .B (n_114_128), .C1 (n_113_127), .C2 (n_110_131) );
AOI211_X1 g_112_128 (.ZN (n_112_128), .A (n_116_126), .B (n_116_127), .C1 (n_112_129), .C2 (n_109_129) );
AOI211_X1 g_110_129 (.ZN (n_110_129), .A (n_114_127), .B (n_115_129), .C1 (n_114_128), .C2 (n_111_128) );
AOI211_X1 g_108_130 (.ZN (n_108_130), .A (n_112_128), .B (n_117_128), .C1 (n_116_127), .C2 (n_113_127) );
AOI211_X1 g_106_131 (.ZN (n_106_131), .A (n_110_129), .B (n_116_126), .C1 (n_115_129), .C2 (n_112_129) );
AOI211_X1 g_104_132 (.ZN (n_104_132), .A (n_108_130), .B (n_114_127), .C1 (n_117_128), .C2 (n_114_128) );
AOI211_X1 g_102_133 (.ZN (n_102_133), .A (n_106_131), .B (n_112_128), .C1 (n_116_126), .C2 (n_116_127) );
AOI211_X1 g_100_134 (.ZN (n_100_134), .A (n_104_132), .B (n_110_129), .C1 (n_114_127), .C2 (n_115_129) );
AOI211_X1 g_98_135 (.ZN (n_98_135), .A (n_102_133), .B (n_108_130), .C1 (n_112_128), .C2 (n_117_128) );
AOI211_X1 g_96_136 (.ZN (n_96_136), .A (n_100_134), .B (n_106_131), .C1 (n_110_129), .C2 (n_116_126) );
AOI211_X1 g_97_134 (.ZN (n_97_134), .A (n_98_135), .B (n_104_132), .C1 (n_108_130), .C2 (n_114_127) );
AOI211_X1 g_95_135 (.ZN (n_95_135), .A (n_96_136), .B (n_102_133), .C1 (n_106_131), .C2 (n_112_128) );
AOI211_X1 g_93_136 (.ZN (n_93_136), .A (n_97_134), .B (n_100_134), .C1 (n_104_132), .C2 (n_110_129) );
AOI211_X1 g_91_137 (.ZN (n_91_137), .A (n_95_135), .B (n_98_135), .C1 (n_102_133), .C2 (n_108_130) );
AOI211_X1 g_89_138 (.ZN (n_89_138), .A (n_93_136), .B (n_96_136), .C1 (n_100_134), .C2 (n_106_131) );
AOI211_X1 g_87_139 (.ZN (n_87_139), .A (n_91_137), .B (n_97_134), .C1 (n_98_135), .C2 (n_104_132) );
AOI211_X1 g_85_140 (.ZN (n_85_140), .A (n_89_138), .B (n_95_135), .C1 (n_96_136), .C2 (n_102_133) );
AOI211_X1 g_86_138 (.ZN (n_86_138), .A (n_87_139), .B (n_93_136), .C1 (n_97_134), .C2 (n_100_134) );
AOI211_X1 g_84_139 (.ZN (n_84_139), .A (n_85_140), .B (n_91_137), .C1 (n_95_135), .C2 (n_98_135) );
AOI211_X1 g_82_140 (.ZN (n_82_140), .A (n_86_138), .B (n_89_138), .C1 (n_93_136), .C2 (n_96_136) );
AOI211_X1 g_80_141 (.ZN (n_80_141), .A (n_84_139), .B (n_87_139), .C1 (n_91_137), .C2 (n_97_134) );
AOI211_X1 g_78_142 (.ZN (n_78_142), .A (n_82_140), .B (n_85_140), .C1 (n_89_138), .C2 (n_95_135) );
AOI211_X1 g_76_143 (.ZN (n_76_143), .A (n_80_141), .B (n_86_138), .C1 (n_87_139), .C2 (n_93_136) );
AOI211_X1 g_74_144 (.ZN (n_74_144), .A (n_78_142), .B (n_84_139), .C1 (n_85_140), .C2 (n_91_137) );
AOI211_X1 g_73_146 (.ZN (n_73_146), .A (n_76_143), .B (n_82_140), .C1 (n_86_138), .C2 (n_89_138) );
AOI211_X1 g_75_145 (.ZN (n_75_145), .A (n_74_144), .B (n_80_141), .C1 (n_84_139), .C2 (n_87_139) );
AOI211_X1 g_77_144 (.ZN (n_77_144), .A (n_73_146), .B (n_78_142), .C1 (n_82_140), .C2 (n_85_140) );
AOI211_X1 g_79_143 (.ZN (n_79_143), .A (n_75_145), .B (n_76_143), .C1 (n_80_141), .C2 (n_86_138) );
AOI211_X1 g_81_142 (.ZN (n_81_142), .A (n_77_144), .B (n_74_144), .C1 (n_78_142), .C2 (n_84_139) );
AOI211_X1 g_83_141 (.ZN (n_83_141), .A (n_79_143), .B (n_73_146), .C1 (n_76_143), .C2 (n_82_140) );
AOI211_X1 g_82_143 (.ZN (n_82_143), .A (n_81_142), .B (n_75_145), .C1 (n_74_144), .C2 (n_80_141) );
AOI211_X1 g_80_142 (.ZN (n_80_142), .A (n_83_141), .B (n_77_144), .C1 (n_73_146), .C2 (n_78_142) );
AOI211_X1 g_78_143 (.ZN (n_78_143), .A (n_82_143), .B (n_79_143), .C1 (n_75_145), .C2 (n_76_143) );
AOI211_X1 g_77_145 (.ZN (n_77_145), .A (n_80_142), .B (n_81_142), .C1 (n_77_144), .C2 (n_74_144) );
AOI211_X1 g_75_146 (.ZN (n_75_146), .A (n_78_143), .B (n_83_141), .C1 (n_79_143), .C2 (n_73_146) );
AOI211_X1 g_74_148 (.ZN (n_74_148), .A (n_77_145), .B (n_82_143), .C1 (n_81_142), .C2 (n_75_145) );
AOI211_X1 g_76_147 (.ZN (n_76_147), .A (n_75_146), .B (n_80_142), .C1 (n_83_141), .C2 (n_77_144) );
AOI211_X1 g_78_148 (.ZN (n_78_148), .A (n_74_148), .B (n_78_143), .C1 (n_82_143), .C2 (n_79_143) );
AOI211_X1 g_76_149 (.ZN (n_76_149), .A (n_76_147), .B (n_77_145), .C1 (n_80_142), .C2 (n_81_142) );
AOI211_X1 g_75_147 (.ZN (n_75_147), .A (n_78_148), .B (n_75_146), .C1 (n_78_143), .C2 (n_83_141) );
AOI211_X1 g_77_146 (.ZN (n_77_146), .A (n_76_149), .B (n_74_148), .C1 (n_77_145), .C2 (n_82_143) );
AOI211_X1 g_79_145 (.ZN (n_79_145), .A (n_75_147), .B (n_76_147), .C1 (n_75_146), .C2 (n_80_142) );
AOI211_X1 g_80_143 (.ZN (n_80_143), .A (n_77_146), .B (n_78_148), .C1 (n_74_148), .C2 (n_78_143) );
AOI211_X1 g_78_144 (.ZN (n_78_144), .A (n_79_145), .B (n_76_149), .C1 (n_76_147), .C2 (n_77_145) );
AOI211_X1 g_76_145 (.ZN (n_76_145), .A (n_80_143), .B (n_75_147), .C1 (n_78_148), .C2 (n_75_146) );
AOI211_X1 g_77_147 (.ZN (n_77_147), .A (n_78_144), .B (n_77_146), .C1 (n_76_149), .C2 (n_74_148) );
AOI211_X1 g_79_146 (.ZN (n_79_146), .A (n_76_145), .B (n_79_145), .C1 (n_75_147), .C2 (n_76_147) );
AOI211_X1 g_80_144 (.ZN (n_80_144), .A (n_77_147), .B (n_80_143), .C1 (n_77_146), .C2 (n_78_148) );
AOI211_X1 g_78_145 (.ZN (n_78_145), .A (n_79_146), .B (n_78_144), .C1 (n_79_145), .C2 (n_76_149) );
AOI211_X1 g_79_147 (.ZN (n_79_147), .A (n_80_144), .B (n_76_145), .C1 (n_80_143), .C2 (n_75_147) );
AOI211_X1 g_77_148 (.ZN (n_77_148), .A (n_78_145), .B (n_77_147), .C1 (n_78_144), .C2 (n_77_146) );
AOI211_X1 g_78_150 (.ZN (n_78_150), .A (n_79_147), .B (n_79_146), .C1 (n_76_145), .C2 (n_79_145) );
AOI211_X1 g_80_149 (.ZN (n_80_149), .A (n_77_148), .B (n_80_144), .C1 (n_77_147), .C2 (n_80_143) );
AOI211_X1 g_82_150 (.ZN (n_82_150), .A (n_78_150), .B (n_78_145), .C1 (n_79_146), .C2 (n_78_144) );
AOI211_X1 g_81_148 (.ZN (n_81_148), .A (n_80_149), .B (n_79_147), .C1 (n_80_144), .C2 (n_76_145) );
AOI211_X1 g_80_146 (.ZN (n_80_146), .A (n_82_150), .B (n_77_148), .C1 (n_78_145), .C2 (n_77_147) );
AOI211_X1 g_79_148 (.ZN (n_79_148), .A (n_81_148), .B (n_78_150), .C1 (n_79_147), .C2 (n_79_146) );
AOI211_X1 g_78_146 (.ZN (n_78_146), .A (n_80_146), .B (n_80_149), .C1 (n_77_148), .C2 (n_80_144) );
AOI211_X1 g_79_144 (.ZN (n_79_144), .A (n_79_148), .B (n_82_150), .C1 (n_78_150), .C2 (n_78_145) );
AOI211_X1 g_81_145 (.ZN (n_81_145), .A (n_78_146), .B (n_81_148), .C1 (n_80_149), .C2 (n_79_147) );
AOI211_X1 g_80_147 (.ZN (n_80_147), .A (n_79_144), .B (n_80_146), .C1 (n_82_150), .C2 (n_77_148) );
AOI211_X1 g_82_148 (.ZN (n_82_148), .A (n_81_145), .B (n_79_148), .C1 (n_81_148), .C2 (n_78_150) );
AOI211_X1 g_81_146 (.ZN (n_81_146), .A (n_80_147), .B (n_78_146), .C1 (n_80_146), .C2 (n_80_149) );
AOI211_X1 g_83_145 (.ZN (n_83_145), .A (n_82_148), .B (n_79_144), .C1 (n_79_148), .C2 (n_82_150) );
AOI211_X1 g_81_144 (.ZN (n_81_144), .A (n_81_146), .B (n_81_145), .C1 (n_78_146), .C2 (n_81_148) );
AOI211_X1 g_82_142 (.ZN (n_82_142), .A (n_83_145), .B (n_80_147), .C1 (n_79_144), .C2 (n_80_146) );
AOI211_X1 g_84_141 (.ZN (n_84_141), .A (n_81_144), .B (n_82_148), .C1 (n_81_145), .C2 (n_79_148) );
AOI211_X1 g_86_140 (.ZN (n_86_140), .A (n_82_142), .B (n_81_146), .C1 (n_80_147), .C2 (n_78_146) );
AOI211_X1 g_88_139 (.ZN (n_88_139), .A (n_84_141), .B (n_83_145), .C1 (n_82_148), .C2 (n_79_144) );
AOI211_X1 g_87_141 (.ZN (n_87_141), .A (n_86_140), .B (n_81_144), .C1 (n_81_146), .C2 (n_81_145) );
AOI211_X1 g_86_139 (.ZN (n_86_139), .A (n_88_139), .B (n_82_142), .C1 (n_83_145), .C2 (n_80_147) );
AOI211_X1 g_88_138 (.ZN (n_88_138), .A (n_87_141), .B (n_84_141), .C1 (n_81_144), .C2 (n_82_148) );
AOI211_X1 g_90_137 (.ZN (n_90_137), .A (n_86_139), .B (n_86_140), .C1 (n_82_142), .C2 (n_81_146) );
AOI211_X1 g_92_136 (.ZN (n_92_136), .A (n_88_138), .B (n_88_139), .C1 (n_84_141), .C2 (n_83_145) );
AOI211_X1 g_94_135 (.ZN (n_94_135), .A (n_90_137), .B (n_87_141), .C1 (n_86_140), .C2 (n_81_144) );
AOI211_X1 g_93_137 (.ZN (n_93_137), .A (n_92_136), .B (n_86_139), .C1 (n_88_139), .C2 (n_82_142) );
AOI211_X1 g_95_136 (.ZN (n_95_136), .A (n_94_135), .B (n_88_138), .C1 (n_87_141), .C2 (n_84_141) );
AOI211_X1 g_97_135 (.ZN (n_97_135), .A (n_93_137), .B (n_90_137), .C1 (n_86_139), .C2 (n_86_140) );
AOI211_X1 g_99_134 (.ZN (n_99_134), .A (n_95_136), .B (n_92_136), .C1 (n_88_138), .C2 (n_88_139) );
AOI211_X1 g_101_133 (.ZN (n_101_133), .A (n_97_135), .B (n_94_135), .C1 (n_90_137), .C2 (n_87_141) );
AOI211_X1 g_103_132 (.ZN (n_103_132), .A (n_99_134), .B (n_93_137), .C1 (n_92_136), .C2 (n_86_139) );
AOI211_X1 g_105_131 (.ZN (n_105_131), .A (n_101_133), .B (n_95_136), .C1 (n_94_135), .C2 (n_88_138) );
AOI211_X1 g_107_130 (.ZN (n_107_130), .A (n_103_132), .B (n_97_135), .C1 (n_93_137), .C2 (n_90_137) );
AOI211_X1 g_108_132 (.ZN (n_108_132), .A (n_105_131), .B (n_99_134), .C1 (n_95_136), .C2 (n_92_136) );
AOI211_X1 g_106_133 (.ZN (n_106_133), .A (n_107_130), .B (n_101_133), .C1 (n_97_135), .C2 (n_94_135) );
AOI211_X1 g_107_131 (.ZN (n_107_131), .A (n_108_132), .B (n_103_132), .C1 (n_99_134), .C2 (n_93_137) );
AOI211_X1 g_105_132 (.ZN (n_105_132), .A (n_106_133), .B (n_105_131), .C1 (n_101_133), .C2 (n_95_136) );
AOI211_X1 g_103_133 (.ZN (n_103_133), .A (n_107_131), .B (n_107_130), .C1 (n_103_132), .C2 (n_97_135) );
AOI211_X1 g_102_135 (.ZN (n_102_135), .A (n_105_132), .B (n_108_132), .C1 (n_105_131), .C2 (n_99_134) );
AOI211_X1 g_104_134 (.ZN (n_104_134), .A (n_103_133), .B (n_106_133), .C1 (n_107_130), .C2 (n_101_133) );
AOI211_X1 g_103_136 (.ZN (n_103_136), .A (n_102_135), .B (n_107_131), .C1 (n_108_132), .C2 (n_103_132) );
AOI211_X1 g_102_134 (.ZN (n_102_134), .A (n_104_134), .B (n_105_132), .C1 (n_106_133), .C2 (n_105_131) );
AOI211_X1 g_104_133 (.ZN (n_104_133), .A (n_103_136), .B (n_103_133), .C1 (n_107_131), .C2 (n_107_130) );
AOI211_X1 g_106_132 (.ZN (n_106_132), .A (n_102_134), .B (n_102_135), .C1 (n_105_132), .C2 (n_108_132) );
AOI211_X1 g_108_131 (.ZN (n_108_131), .A (n_104_133), .B (n_104_134), .C1 (n_103_133), .C2 (n_106_133) );
AOI211_X1 g_110_130 (.ZN (n_110_130), .A (n_106_132), .B (n_103_136), .C1 (n_102_135), .C2 (n_107_131) );
AOI211_X1 g_109_132 (.ZN (n_109_132), .A (n_108_131), .B (n_102_134), .C1 (n_104_134), .C2 (n_105_132) );
AOI211_X1 g_111_131 (.ZN (n_111_131), .A (n_110_130), .B (n_104_133), .C1 (n_103_136), .C2 (n_103_133) );
AOI211_X1 g_113_130 (.ZN (n_113_130), .A (n_109_132), .B (n_106_132), .C1 (n_102_134), .C2 (n_102_135) );
AOI211_X1 g_112_132 (.ZN (n_112_132), .A (n_111_131), .B (n_108_131), .C1 (n_104_133), .C2 (n_104_134) );
AOI211_X1 g_111_130 (.ZN (n_111_130), .A (n_113_130), .B (n_110_130), .C1 (n_106_132), .C2 (n_103_136) );
AOI211_X1 g_113_129 (.ZN (n_113_129), .A (n_112_132), .B (n_109_132), .C1 (n_108_131), .C2 (n_102_134) );
AOI211_X1 g_115_128 (.ZN (n_115_128), .A (n_111_130), .B (n_111_131), .C1 (n_110_130), .C2 (n_104_133) );
AOI211_X1 g_117_127 (.ZN (n_117_127), .A (n_113_129), .B (n_113_130), .C1 (n_109_132), .C2 (n_106_132) );
AOI211_X1 g_119_126 (.ZN (n_119_126), .A (n_115_128), .B (n_112_132), .C1 (n_111_131), .C2 (n_108_131) );
AOI211_X1 g_121_125 (.ZN (n_121_125), .A (n_117_127), .B (n_111_130), .C1 (n_113_130), .C2 (n_110_130) );
AOI211_X1 g_123_124 (.ZN (n_123_124), .A (n_119_126), .B (n_113_129), .C1 (n_112_132), .C2 (n_109_132) );
AOI211_X1 g_125_123 (.ZN (n_125_123), .A (n_121_125), .B (n_115_128), .C1 (n_111_130), .C2 (n_111_131) );
AOI211_X1 g_127_122 (.ZN (n_127_122), .A (n_123_124), .B (n_117_127), .C1 (n_113_129), .C2 (n_113_130) );
AOI211_X1 g_129_121 (.ZN (n_129_121), .A (n_125_123), .B (n_119_126), .C1 (n_115_128), .C2 (n_112_132) );
AOI211_X1 g_128_123 (.ZN (n_128_123), .A (n_127_122), .B (n_121_125), .C1 (n_117_127), .C2 (n_111_130) );
AOI211_X1 g_130_122 (.ZN (n_130_122), .A (n_129_121), .B (n_123_124), .C1 (n_119_126), .C2 (n_113_129) );
AOI211_X1 g_132_121 (.ZN (n_132_121), .A (n_128_123), .B (n_125_123), .C1 (n_121_125), .C2 (n_115_128) );
AOI211_X1 g_131_123 (.ZN (n_131_123), .A (n_130_122), .B (n_127_122), .C1 (n_123_124), .C2 (n_117_127) );
AOI211_X1 g_133_122 (.ZN (n_133_122), .A (n_132_121), .B (n_129_121), .C1 (n_125_123), .C2 (n_119_126) );
AOI211_X1 g_132_120 (.ZN (n_132_120), .A (n_131_123), .B (n_128_123), .C1 (n_127_122), .C2 (n_121_125) );
AOI211_X1 g_134_119 (.ZN (n_134_119), .A (n_133_122), .B (n_130_122), .C1 (n_129_121), .C2 (n_123_124) );
AOI211_X1 g_136_118 (.ZN (n_136_118), .A (n_132_120), .B (n_132_121), .C1 (n_128_123), .C2 (n_125_123) );
AOI211_X1 g_138_117 (.ZN (n_138_117), .A (n_134_119), .B (n_131_123), .C1 (n_130_122), .C2 (n_127_122) );
AOI211_X1 g_137_119 (.ZN (n_137_119), .A (n_136_118), .B (n_133_122), .C1 (n_132_121), .C2 (n_129_121) );
AOI211_X1 g_139_118 (.ZN (n_139_118), .A (n_138_117), .B (n_132_120), .C1 (n_131_123), .C2 (n_128_123) );
AOI211_X1 g_141_117 (.ZN (n_141_117), .A (n_137_119), .B (n_134_119), .C1 (n_133_122), .C2 (n_130_122) );
AOI211_X1 g_139_116 (.ZN (n_139_116), .A (n_139_118), .B (n_136_118), .C1 (n_132_120), .C2 (n_132_121) );
AOI211_X1 g_141_115 (.ZN (n_141_115), .A (n_141_117), .B (n_138_117), .C1 (n_134_119), .C2 (n_131_123) );
AOI211_X1 g_143_116 (.ZN (n_143_116), .A (n_139_116), .B (n_137_119), .C1 (n_136_118), .C2 (n_133_122) );
AOI211_X1 g_145_117 (.ZN (n_145_117), .A (n_141_115), .B (n_139_118), .C1 (n_138_117), .C2 (n_132_120) );
AOI211_X1 g_144_115 (.ZN (n_144_115), .A (n_143_116), .B (n_141_117), .C1 (n_137_119), .C2 (n_134_119) );
AOI211_X1 g_146_116 (.ZN (n_146_116), .A (n_145_117), .B (n_139_116), .C1 (n_139_118), .C2 (n_136_118) );
AOI211_X1 g_144_117 (.ZN (n_144_117), .A (n_144_115), .B (n_141_115), .C1 (n_141_117), .C2 (n_138_117) );
AOI211_X1 g_142_116 (.ZN (n_142_116), .A (n_146_116), .B (n_143_116), .C1 (n_139_116), .C2 (n_137_119) );
AOI211_X1 g_143_118 (.ZN (n_143_118), .A (n_144_117), .B (n_145_117), .C1 (n_141_115), .C2 (n_139_118) );
AOI211_X1 g_141_119 (.ZN (n_141_119), .A (n_142_116), .B (n_144_115), .C1 (n_143_116), .C2 (n_141_117) );
AOI211_X1 g_142_117 (.ZN (n_142_117), .A (n_143_118), .B (n_146_116), .C1 (n_145_117), .C2 (n_139_116) );
AOI211_X1 g_140_118 (.ZN (n_140_118), .A (n_141_119), .B (n_144_117), .C1 (n_144_115), .C2 (n_141_115) );
AOI211_X1 g_138_119 (.ZN (n_138_119), .A (n_142_117), .B (n_142_116), .C1 (n_146_116), .C2 (n_143_116) );
AOI211_X1 g_136_120 (.ZN (n_136_120), .A (n_140_118), .B (n_143_118), .C1 (n_144_117), .C2 (n_145_117) );
AOI211_X1 g_134_121 (.ZN (n_134_121), .A (n_138_119), .B (n_141_119), .C1 (n_142_116), .C2 (n_144_115) );
AOI211_X1 g_132_122 (.ZN (n_132_122), .A (n_136_120), .B (n_142_117), .C1 (n_143_118), .C2 (n_146_116) );
AOI211_X1 g_130_123 (.ZN (n_130_123), .A (n_134_121), .B (n_140_118), .C1 (n_141_119), .C2 (n_144_117) );
AOI211_X1 g_128_124 (.ZN (n_128_124), .A (n_132_122), .B (n_138_119), .C1 (n_142_117), .C2 (n_142_116) );
AOI211_X1 g_126_125 (.ZN (n_126_125), .A (n_130_123), .B (n_136_120), .C1 (n_140_118), .C2 (n_143_118) );
AOI211_X1 g_127_123 (.ZN (n_127_123), .A (n_128_124), .B (n_134_121), .C1 (n_138_119), .C2 (n_141_119) );
AOI211_X1 g_125_124 (.ZN (n_125_124), .A (n_126_125), .B (n_132_122), .C1 (n_136_120), .C2 (n_142_117) );
AOI211_X1 g_123_125 (.ZN (n_123_125), .A (n_127_123), .B (n_130_123), .C1 (n_134_121), .C2 (n_140_118) );
AOI211_X1 g_121_126 (.ZN (n_121_126), .A (n_125_124), .B (n_128_124), .C1 (n_132_122), .C2 (n_138_119) );
AOI211_X1 g_120_128 (.ZN (n_120_128), .A (n_123_125), .B (n_126_125), .C1 (n_130_123), .C2 (n_136_120) );
AOI211_X1 g_118_127 (.ZN (n_118_127), .A (n_121_126), .B (n_127_123), .C1 (n_128_124), .C2 (n_134_121) );
AOI211_X1 g_120_126 (.ZN (n_120_126), .A (n_120_128), .B (n_125_124), .C1 (n_126_125), .C2 (n_132_122) );
AOI211_X1 g_122_125 (.ZN (n_122_125), .A (n_118_127), .B (n_123_125), .C1 (n_127_123), .C2 (n_130_123) );
AOI211_X1 g_124_124 (.ZN (n_124_124), .A (n_120_126), .B (n_121_126), .C1 (n_125_124), .C2 (n_128_124) );
AOI211_X1 g_123_126 (.ZN (n_123_126), .A (n_122_125), .B (n_120_128), .C1 (n_123_125), .C2 (n_126_125) );
AOI211_X1 g_125_125 (.ZN (n_125_125), .A (n_124_124), .B (n_118_127), .C1 (n_121_126), .C2 (n_127_123) );
AOI211_X1 g_127_124 (.ZN (n_127_124), .A (n_123_126), .B (n_120_126), .C1 (n_120_128), .C2 (n_125_124) );
AOI211_X1 g_129_123 (.ZN (n_129_123), .A (n_125_125), .B (n_122_125), .C1 (n_118_127), .C2 (n_123_125) );
AOI211_X1 g_131_122 (.ZN (n_131_122), .A (n_127_124), .B (n_124_124), .C1 (n_120_126), .C2 (n_121_126) );
AOI211_X1 g_133_121 (.ZN (n_133_121), .A (n_129_123), .B (n_123_126), .C1 (n_122_125), .C2 (n_120_128) );
AOI211_X1 g_135_120 (.ZN (n_135_120), .A (n_131_122), .B (n_125_125), .C1 (n_124_124), .C2 (n_118_127) );
AOI211_X1 g_134_122 (.ZN (n_134_122), .A (n_133_121), .B (n_127_124), .C1 (n_123_126), .C2 (n_120_126) );
AOI211_X1 g_136_121 (.ZN (n_136_121), .A (n_135_120), .B (n_129_123), .C1 (n_125_125), .C2 (n_122_125) );
AOI211_X1 g_138_120 (.ZN (n_138_120), .A (n_134_122), .B (n_131_122), .C1 (n_127_124), .C2 (n_124_124) );
AOI211_X1 g_136_119 (.ZN (n_136_119), .A (n_136_121), .B (n_133_121), .C1 (n_129_123), .C2 (n_123_126) );
AOI211_X1 g_138_118 (.ZN (n_138_118), .A (n_138_120), .B (n_135_120), .C1 (n_131_122), .C2 (n_125_125) );
AOI211_X1 g_140_117 (.ZN (n_140_117), .A (n_136_119), .B (n_134_122), .C1 (n_133_121), .C2 (n_127_124) );
AOI211_X1 g_142_118 (.ZN (n_142_118), .A (n_138_118), .B (n_136_121), .C1 (n_135_120), .C2 (n_129_123) );
AOI211_X1 g_140_119 (.ZN (n_140_119), .A (n_140_117), .B (n_138_120), .C1 (n_134_122), .C2 (n_131_122) );
AOI211_X1 g_139_121 (.ZN (n_139_121), .A (n_142_118), .B (n_136_119), .C1 (n_136_121), .C2 (n_133_121) );
AOI211_X1 g_137_120 (.ZN (n_137_120), .A (n_140_119), .B (n_138_118), .C1 (n_138_120), .C2 (n_135_120) );
AOI211_X1 g_135_121 (.ZN (n_135_121), .A (n_139_121), .B (n_140_117), .C1 (n_136_119), .C2 (n_134_122) );
AOI211_X1 g_137_122 (.ZN (n_137_122), .A (n_137_120), .B (n_142_118), .C1 (n_138_118), .C2 (n_136_121) );
AOI211_X1 g_135_123 (.ZN (n_135_123), .A (n_135_121), .B (n_140_119), .C1 (n_140_117), .C2 (n_138_120) );
AOI211_X1 g_133_124 (.ZN (n_133_124), .A (n_137_122), .B (n_139_121), .C1 (n_142_118), .C2 (n_136_119) );
AOI211_X1 g_131_125 (.ZN (n_131_125), .A (n_135_123), .B (n_137_120), .C1 (n_140_119), .C2 (n_138_118) );
AOI211_X1 g_132_123 (.ZN (n_132_123), .A (n_133_124), .B (n_135_121), .C1 (n_139_121), .C2 (n_140_117) );
AOI211_X1 g_130_124 (.ZN (n_130_124), .A (n_131_125), .B (n_137_122), .C1 (n_137_120), .C2 (n_142_118) );
AOI211_X1 g_128_125 (.ZN (n_128_125), .A (n_132_123), .B (n_135_123), .C1 (n_135_121), .C2 (n_140_119) );
AOI211_X1 g_126_124 (.ZN (n_126_124), .A (n_130_124), .B (n_133_124), .C1 (n_137_122), .C2 (n_139_121) );
AOI211_X1 g_124_125 (.ZN (n_124_125), .A (n_128_125), .B (n_131_125), .C1 (n_135_123), .C2 (n_137_120) );
AOI211_X1 g_122_126 (.ZN (n_122_126), .A (n_126_124), .B (n_132_123), .C1 (n_133_124), .C2 (n_135_121) );
AOI211_X1 g_120_127 (.ZN (n_120_127), .A (n_124_125), .B (n_130_124), .C1 (n_131_125), .C2 (n_137_122) );
AOI211_X1 g_118_128 (.ZN (n_118_128), .A (n_122_126), .B (n_128_125), .C1 (n_132_123), .C2 (n_135_123) );
AOI211_X1 g_116_129 (.ZN (n_116_129), .A (n_120_127), .B (n_126_124), .C1 (n_130_124), .C2 (n_133_124) );
AOI211_X1 g_114_130 (.ZN (n_114_130), .A (n_118_128), .B (n_124_125), .C1 (n_128_125), .C2 (n_131_125) );
AOI211_X1 g_112_131 (.ZN (n_112_131), .A (n_116_129), .B (n_122_126), .C1 (n_126_124), .C2 (n_132_123) );
AOI211_X1 g_110_132 (.ZN (n_110_132), .A (n_114_130), .B (n_120_127), .C1 (n_124_125), .C2 (n_130_124) );
AOI211_X1 g_108_133 (.ZN (n_108_133), .A (n_112_131), .B (n_118_128), .C1 (n_122_126), .C2 (n_128_125) );
AOI211_X1 g_109_131 (.ZN (n_109_131), .A (n_110_132), .B (n_116_129), .C1 (n_120_127), .C2 (n_126_124) );
AOI211_X1 g_107_132 (.ZN (n_107_132), .A (n_108_133), .B (n_114_130), .C1 (n_118_128), .C2 (n_124_125) );
AOI211_X1 g_105_133 (.ZN (n_105_133), .A (n_109_131), .B (n_112_131), .C1 (n_116_129), .C2 (n_122_126) );
AOI211_X1 g_103_134 (.ZN (n_103_134), .A (n_107_132), .B (n_110_132), .C1 (n_114_130), .C2 (n_120_127) );
AOI211_X1 g_101_135 (.ZN (n_101_135), .A (n_105_133), .B (n_108_133), .C1 (n_112_131), .C2 (n_118_128) );
AOI211_X1 g_99_136 (.ZN (n_99_136), .A (n_103_134), .B (n_109_131), .C1 (n_110_132), .C2 (n_116_129) );
AOI211_X1 g_98_134 (.ZN (n_98_134), .A (n_101_135), .B (n_107_132), .C1 (n_108_133), .C2 (n_114_130) );
AOI211_X1 g_96_135 (.ZN (n_96_135), .A (n_99_136), .B (n_105_133), .C1 (n_109_131), .C2 (n_112_131) );
AOI211_X1 g_94_136 (.ZN (n_94_136), .A (n_98_134), .B (n_103_134), .C1 (n_107_132), .C2 (n_110_132) );
AOI211_X1 g_92_137 (.ZN (n_92_137), .A (n_96_135), .B (n_101_135), .C1 (n_105_133), .C2 (n_108_133) );
AOI211_X1 g_91_139 (.ZN (n_91_139), .A (n_94_136), .B (n_99_136), .C1 (n_103_134), .C2 (n_109_131) );
AOI211_X1 g_89_140 (.ZN (n_89_140), .A (n_92_137), .B (n_98_134), .C1 (n_101_135), .C2 (n_107_132) );
AOI211_X1 g_88_142 (.ZN (n_88_142), .A (n_91_139), .B (n_96_135), .C1 (n_99_136), .C2 (n_105_133) );
AOI211_X1 g_87_140 (.ZN (n_87_140), .A (n_89_140), .B (n_94_136), .C1 (n_98_134), .C2 (n_103_134) );
AOI211_X1 g_89_139 (.ZN (n_89_139), .A (n_88_142), .B (n_92_137), .C1 (n_96_135), .C2 (n_101_135) );
AOI211_X1 g_91_138 (.ZN (n_91_138), .A (n_87_140), .B (n_91_139), .C1 (n_94_136), .C2 (n_99_136) );
AOI211_X1 g_90_140 (.ZN (n_90_140), .A (n_89_139), .B (n_89_140), .C1 (n_92_137), .C2 (n_98_134) );
AOI211_X1 g_92_139 (.ZN (n_92_139), .A (n_91_138), .B (n_88_142), .C1 (n_91_139), .C2 (n_96_135) );
AOI211_X1 g_94_138 (.ZN (n_94_138), .A (n_90_140), .B (n_87_140), .C1 (n_89_140), .C2 (n_94_136) );
AOI211_X1 g_96_137 (.ZN (n_96_137), .A (n_92_139), .B (n_89_139), .C1 (n_88_142), .C2 (n_92_137) );
AOI211_X1 g_98_136 (.ZN (n_98_136), .A (n_94_138), .B (n_91_138), .C1 (n_87_140), .C2 (n_91_139) );
AOI211_X1 g_100_135 (.ZN (n_100_135), .A (n_96_137), .B (n_90_140), .C1 (n_89_139), .C2 (n_89_140) );
AOI211_X1 g_101_137 (.ZN (n_101_137), .A (n_98_136), .B (n_92_139), .C1 (n_91_138), .C2 (n_88_142) );
AOI211_X1 g_99_138 (.ZN (n_99_138), .A (n_100_135), .B (n_94_138), .C1 (n_90_140), .C2 (n_87_140) );
AOI211_X1 g_100_136 (.ZN (n_100_136), .A (n_101_137), .B (n_96_137), .C1 (n_92_139), .C2 (n_89_139) );
AOI211_X1 g_98_137 (.ZN (n_98_137), .A (n_99_138), .B (n_98_136), .C1 (n_94_138), .C2 (n_91_138) );
AOI211_X1 g_99_135 (.ZN (n_99_135), .A (n_100_136), .B (n_100_135), .C1 (n_96_137), .C2 (n_90_140) );
AOI211_X1 g_97_136 (.ZN (n_97_136), .A (n_98_137), .B (n_101_137), .C1 (n_98_136), .C2 (n_92_139) );
AOI211_X1 g_95_137 (.ZN (n_95_137), .A (n_99_135), .B (n_99_138), .C1 (n_100_135), .C2 (n_94_138) );
AOI211_X1 g_93_138 (.ZN (n_93_138), .A (n_97_136), .B (n_100_136), .C1 (n_101_137), .C2 (n_96_137) );
AOI211_X1 g_92_140 (.ZN (n_92_140), .A (n_95_137), .B (n_98_137), .C1 (n_99_138), .C2 (n_98_136) );
AOI211_X1 g_90_139 (.ZN (n_90_139), .A (n_93_138), .B (n_99_135), .C1 (n_100_136), .C2 (n_100_135) );
AOI211_X1 g_92_138 (.ZN (n_92_138), .A (n_92_140), .B (n_97_136), .C1 (n_98_137), .C2 (n_101_137) );
AOI211_X1 g_94_137 (.ZN (n_94_137), .A (n_90_139), .B (n_95_137), .C1 (n_99_135), .C2 (n_99_138) );
AOI211_X1 g_96_138 (.ZN (n_96_138), .A (n_92_138), .B (n_93_138), .C1 (n_97_136), .C2 (n_100_136) );
AOI211_X1 g_94_139 (.ZN (n_94_139), .A (n_94_137), .B (n_92_140), .C1 (n_95_137), .C2 (n_98_137) );
AOI211_X1 g_93_141 (.ZN (n_93_141), .A (n_96_138), .B (n_90_139), .C1 (n_93_138), .C2 (n_99_135) );
AOI211_X1 g_91_140 (.ZN (n_91_140), .A (n_94_139), .B (n_92_138), .C1 (n_92_140), .C2 (n_97_136) );
AOI211_X1 g_93_139 (.ZN (n_93_139), .A (n_93_141), .B (n_94_137), .C1 (n_90_139), .C2 (n_95_137) );
AOI211_X1 g_95_138 (.ZN (n_95_138), .A (n_91_140), .B (n_96_138), .C1 (n_92_138), .C2 (n_93_138) );
AOI211_X1 g_97_137 (.ZN (n_97_137), .A (n_93_139), .B (n_94_139), .C1 (n_94_137), .C2 (n_92_140) );
AOI211_X1 g_96_139 (.ZN (n_96_139), .A (n_95_138), .B (n_93_141), .C1 (n_96_138), .C2 (n_90_139) );
AOI211_X1 g_98_138 (.ZN (n_98_138), .A (n_97_137), .B (n_91_140), .C1 (n_94_139), .C2 (n_92_138) );
AOI211_X1 g_100_137 (.ZN (n_100_137), .A (n_96_139), .B (n_93_139), .C1 (n_93_141), .C2 (n_94_137) );
AOI211_X1 g_102_136 (.ZN (n_102_136), .A (n_98_138), .B (n_95_138), .C1 (n_91_140), .C2 (n_96_138) );
AOI211_X1 g_104_135 (.ZN (n_104_135), .A (n_100_137), .B (n_97_137), .C1 (n_93_139), .C2 (n_94_139) );
AOI211_X1 g_106_134 (.ZN (n_106_134), .A (n_102_136), .B (n_96_139), .C1 (n_95_138), .C2 (n_93_141) );
AOI211_X1 g_105_136 (.ZN (n_105_136), .A (n_104_135), .B (n_98_138), .C1 (n_97_137), .C2 (n_91_140) );
AOI211_X1 g_103_135 (.ZN (n_103_135), .A (n_106_134), .B (n_100_137), .C1 (n_96_139), .C2 (n_93_139) );
AOI211_X1 g_105_134 (.ZN (n_105_134), .A (n_105_136), .B (n_102_136), .C1 (n_98_138), .C2 (n_95_138) );
AOI211_X1 g_107_133 (.ZN (n_107_133), .A (n_103_135), .B (n_104_135), .C1 (n_100_137), .C2 (n_97_137) );
AOI211_X1 g_106_135 (.ZN (n_106_135), .A (n_105_134), .B (n_106_134), .C1 (n_102_136), .C2 (n_96_139) );
AOI211_X1 g_108_134 (.ZN (n_108_134), .A (n_107_133), .B (n_105_136), .C1 (n_104_135), .C2 (n_98_138) );
AOI211_X1 g_110_133 (.ZN (n_110_133), .A (n_106_135), .B (n_103_135), .C1 (n_106_134), .C2 (n_100_137) );
AOI211_X1 g_109_135 (.ZN (n_109_135), .A (n_108_134), .B (n_105_134), .C1 (n_105_136), .C2 (n_102_136) );
AOI211_X1 g_107_134 (.ZN (n_107_134), .A (n_110_133), .B (n_107_133), .C1 (n_103_135), .C2 (n_104_135) );
AOI211_X1 g_105_135 (.ZN (n_105_135), .A (n_109_135), .B (n_106_135), .C1 (n_105_134), .C2 (n_106_134) );
AOI211_X1 g_107_136 (.ZN (n_107_136), .A (n_107_134), .B (n_108_134), .C1 (n_107_133), .C2 (n_105_136) );
AOI211_X1 g_105_137 (.ZN (n_105_137), .A (n_105_135), .B (n_110_133), .C1 (n_106_135), .C2 (n_103_135) );
AOI211_X1 g_103_138 (.ZN (n_103_138), .A (n_107_136), .B (n_109_135), .C1 (n_108_134), .C2 (n_105_134) );
AOI211_X1 g_104_136 (.ZN (n_104_136), .A (n_105_137), .B (n_107_134), .C1 (n_110_133), .C2 (n_107_133) );
AOI211_X1 g_102_137 (.ZN (n_102_137), .A (n_103_138), .B (n_105_135), .C1 (n_109_135), .C2 (n_106_135) );
AOI211_X1 g_101_139 (.ZN (n_101_139), .A (n_104_136), .B (n_107_136), .C1 (n_107_134), .C2 (n_108_134) );
AOI211_X1 g_99_140 (.ZN (n_99_140), .A (n_102_137), .B (n_105_137), .C1 (n_105_135), .C2 (n_110_133) );
AOI211_X1 g_97_139 (.ZN (n_97_139), .A (n_101_139), .B (n_103_138), .C1 (n_107_136), .C2 (n_109_135) );
AOI211_X1 g_95_140 (.ZN (n_95_140), .A (n_99_140), .B (n_104_136), .C1 (n_105_137), .C2 (n_107_134) );
AOI211_X1 g_97_141 (.ZN (n_97_141), .A (n_97_139), .B (n_102_137), .C1 (n_103_138), .C2 (n_105_135) );
AOI211_X1 g_98_139 (.ZN (n_98_139), .A (n_95_140), .B (n_101_139), .C1 (n_104_136), .C2 (n_107_136) );
AOI211_X1 g_100_138 (.ZN (n_100_138), .A (n_97_141), .B (n_99_140), .C1 (n_102_137), .C2 (n_105_137) );
AOI211_X1 g_101_136 (.ZN (n_101_136), .A (n_98_139), .B (n_97_139), .C1 (n_101_139), .C2 (n_103_138) );
AOI211_X1 g_99_137 (.ZN (n_99_137), .A (n_100_138), .B (n_95_140), .C1 (n_99_140), .C2 (n_104_136) );
AOI211_X1 g_97_138 (.ZN (n_97_138), .A (n_101_136), .B (n_97_141), .C1 (n_97_139), .C2 (n_102_137) );
AOI211_X1 g_95_139 (.ZN (n_95_139), .A (n_99_137), .B (n_98_139), .C1 (n_95_140), .C2 (n_101_139) );
AOI211_X1 g_93_140 (.ZN (n_93_140), .A (n_97_138), .B (n_100_138), .C1 (n_97_141), .C2 (n_99_140) );
AOI211_X1 g_91_141 (.ZN (n_91_141), .A (n_95_139), .B (n_101_136), .C1 (n_98_139), .C2 (n_97_139) );
AOI211_X1 g_89_142 (.ZN (n_89_142), .A (n_93_140), .B (n_99_137), .C1 (n_100_138), .C2 (n_95_140) );
AOI211_X1 g_88_140 (.ZN (n_88_140), .A (n_91_141), .B (n_97_138), .C1 (n_101_136), .C2 (n_97_141) );
AOI211_X1 g_90_141 (.ZN (n_90_141), .A (n_89_142), .B (n_95_139), .C1 (n_99_137), .C2 (n_98_139) );
AOI211_X1 g_92_142 (.ZN (n_92_142), .A (n_88_140), .B (n_93_140), .C1 (n_97_138), .C2 (n_100_138) );
AOI211_X1 g_94_141 (.ZN (n_94_141), .A (n_90_141), .B (n_91_141), .C1 (n_95_139), .C2 (n_101_136) );
AOI211_X1 g_96_140 (.ZN (n_96_140), .A (n_92_142), .B (n_89_142), .C1 (n_93_140), .C2 (n_99_137) );
AOI211_X1 g_95_142 (.ZN (n_95_142), .A (n_94_141), .B (n_88_140), .C1 (n_91_141), .C2 (n_97_138) );
AOI211_X1 g_94_140 (.ZN (n_94_140), .A (n_96_140), .B (n_90_141), .C1 (n_89_142), .C2 (n_95_139) );
AOI211_X1 g_92_141 (.ZN (n_92_141), .A (n_95_142), .B (n_92_142), .C1 (n_88_140), .C2 (n_93_140) );
AOI211_X1 g_90_142 (.ZN (n_90_142), .A (n_94_140), .B (n_94_141), .C1 (n_90_141), .C2 (n_91_141) );
AOI211_X1 g_88_141 (.ZN (n_88_141), .A (n_92_141), .B (n_96_140), .C1 (n_92_142), .C2 (n_89_142) );
AOI211_X1 g_86_142 (.ZN (n_86_142), .A (n_90_142), .B (n_95_142), .C1 (n_94_141), .C2 (n_88_140) );
AOI211_X1 g_84_143 (.ZN (n_84_143), .A (n_88_141), .B (n_94_140), .C1 (n_96_140), .C2 (n_90_141) );
AOI211_X1 g_85_141 (.ZN (n_85_141), .A (n_86_142), .B (n_92_141), .C1 (n_95_142), .C2 (n_92_142) );
AOI211_X1 g_83_142 (.ZN (n_83_142), .A (n_84_143), .B (n_90_142), .C1 (n_94_140), .C2 (n_94_141) );
AOI211_X1 g_84_140 (.ZN (n_84_140), .A (n_85_141), .B (n_88_141), .C1 (n_92_141), .C2 (n_96_140) );
AOI211_X1 g_82_141 (.ZN (n_82_141), .A (n_83_142), .B (n_86_142), .C1 (n_90_142), .C2 (n_95_142) );
AOI211_X1 g_81_143 (.ZN (n_81_143), .A (n_84_140), .B (n_84_143), .C1 (n_88_141), .C2 (n_94_140) );
AOI211_X1 g_80_145 (.ZN (n_80_145), .A (n_82_141), .B (n_85_141), .C1 (n_86_142), .C2 (n_92_141) );
AOI211_X1 g_82_144 (.ZN (n_82_144), .A (n_81_143), .B (n_83_142), .C1 (n_84_143), .C2 (n_90_142) );
AOI211_X1 g_83_146 (.ZN (n_83_146), .A (n_80_145), .B (n_84_140), .C1 (n_85_141), .C2 (n_88_141) );
AOI211_X1 g_81_147 (.ZN (n_81_147), .A (n_82_144), .B (n_82_141), .C1 (n_83_142), .C2 (n_86_142) );
AOI211_X1 g_83_148 (.ZN (n_83_148), .A (n_83_146), .B (n_81_143), .C1 (n_84_140), .C2 (n_84_143) );
AOI211_X1 g_82_146 (.ZN (n_82_146), .A (n_81_147), .B (n_80_145), .C1 (n_82_141), .C2 (n_85_141) );
AOI211_X1 g_84_147 (.ZN (n_84_147), .A (n_83_148), .B (n_82_144), .C1 (n_81_143), .C2 (n_83_142) );
AOI211_X1 g_85_145 (.ZN (n_85_145), .A (n_82_146), .B (n_83_146), .C1 (n_80_145), .C2 (n_84_140) );
AOI211_X1 g_83_144 (.ZN (n_83_144), .A (n_84_147), .B (n_81_147), .C1 (n_82_144), .C2 (n_82_141) );
AOI211_X1 g_84_142 (.ZN (n_84_142), .A (n_85_145), .B (n_83_148), .C1 (n_83_146), .C2 (n_81_143) );
AOI211_X1 g_86_141 (.ZN (n_86_141), .A (n_83_144), .B (n_82_146), .C1 (n_81_147), .C2 (n_80_145) );
AOI211_X1 g_85_143 (.ZN (n_85_143), .A (n_84_142), .B (n_84_147), .C1 (n_83_148), .C2 (n_82_144) );
AOI211_X1 g_87_142 (.ZN (n_87_142), .A (n_86_141), .B (n_85_145), .C1 (n_82_146), .C2 (n_83_146) );
AOI211_X1 g_89_141 (.ZN (n_89_141), .A (n_85_143), .B (n_83_144), .C1 (n_84_147), .C2 (n_81_147) );
AOI211_X1 g_88_143 (.ZN (n_88_143), .A (n_87_142), .B (n_84_142), .C1 (n_85_145), .C2 (n_83_148) );
AOI211_X1 g_86_144 (.ZN (n_86_144), .A (n_89_141), .B (n_86_141), .C1 (n_83_144), .C2 (n_82_146) );
AOI211_X1 g_85_142 (.ZN (n_85_142), .A (n_88_143), .B (n_85_143), .C1 (n_84_142), .C2 (n_84_147) );
AOI211_X1 g_83_143 (.ZN (n_83_143), .A (n_86_144), .B (n_87_142), .C1 (n_86_141), .C2 (n_85_145) );
AOI211_X1 g_82_145 (.ZN (n_82_145), .A (n_85_142), .B (n_89_141), .C1 (n_85_143), .C2 (n_83_144) );
AOI211_X1 g_84_144 (.ZN (n_84_144), .A (n_83_143), .B (n_88_143), .C1 (n_87_142), .C2 (n_84_142) );
AOI211_X1 g_86_143 (.ZN (n_86_143), .A (n_82_145), .B (n_86_144), .C1 (n_89_141), .C2 (n_86_141) );
AOI211_X1 g_87_145 (.ZN (n_87_145), .A (n_84_144), .B (n_85_142), .C1 (n_88_143), .C2 (n_85_143) );
AOI211_X1 g_85_144 (.ZN (n_85_144), .A (n_86_143), .B (n_83_143), .C1 (n_86_144), .C2 (n_87_142) );
AOI211_X1 g_84_146 (.ZN (n_84_146), .A (n_87_145), .B (n_82_145), .C1 (n_85_142), .C2 (n_89_141) );
AOI211_X1 g_85_148 (.ZN (n_85_148), .A (n_85_144), .B (n_84_144), .C1 (n_83_143), .C2 (n_88_143) );
AOI211_X1 g_83_147 (.ZN (n_83_147), .A (n_84_146), .B (n_86_143), .C1 (n_82_145), .C2 (n_86_144) );
AOI211_X1 g_85_146 (.ZN (n_85_146), .A (n_85_148), .B (n_87_145), .C1 (n_84_144), .C2 (n_85_142) );
AOI211_X1 g_86_148 (.ZN (n_86_148), .A (n_83_147), .B (n_85_144), .C1 (n_86_143), .C2 (n_83_143) );
AOI211_X1 g_84_149 (.ZN (n_84_149), .A (n_85_146), .B (n_84_146), .C1 (n_87_145), .C2 (n_82_145) );
AOI211_X1 g_86_150 (.ZN (n_86_150), .A (n_86_148), .B (n_85_148), .C1 (n_85_144), .C2 (n_84_144) );
AOI211_X1 g_88_149 (.ZN (n_88_149), .A (n_84_149), .B (n_83_147), .C1 (n_84_146), .C2 (n_86_143) );
AOI211_X1 g_90_150 (.ZN (n_90_150), .A (n_86_150), .B (n_85_146), .C1 (n_85_148), .C2 (n_87_145) );
AOI211_X1 g_91_148 (.ZN (n_91_148), .A (n_88_149), .B (n_86_148), .C1 (n_83_147), .C2 (n_85_144) );
AOI211_X1 g_92_146 (.ZN (n_92_146), .A (n_90_150), .B (n_84_149), .C1 (n_85_146), .C2 (n_84_146) );
AOI211_X1 g_93_148 (.ZN (n_93_148), .A (n_91_148), .B (n_86_150), .C1 (n_86_148), .C2 (n_85_148) );
AOI211_X1 g_94_150 (.ZN (n_94_150), .A (n_92_146), .B (n_88_149), .C1 (n_84_149), .C2 (n_83_147) );
AOI211_X1 g_95_148 (.ZN (n_95_148), .A (n_93_148), .B (n_90_150), .C1 (n_86_150), .C2 (n_85_146) );
AOI211_X1 g_96_146 (.ZN (n_96_146), .A (n_94_150), .B (n_91_148), .C1 (n_88_149), .C2 (n_86_148) );
AOI211_X1 g_97_148 (.ZN (n_97_148), .A (n_95_148), .B (n_92_146), .C1 (n_90_150), .C2 (n_84_149) );
AOI211_X1 g_98_150 (.ZN (n_98_150), .A (n_96_146), .B (n_93_148), .C1 (n_91_148), .C2 (n_86_150) );
AOI211_X1 g_99_148 (.ZN (n_99_148), .A (n_97_148), .B (n_94_150), .C1 (n_92_146), .C2 (n_88_149) );
AOI211_X1 g_100_146 (.ZN (n_100_146), .A (n_98_150), .B (n_95_148), .C1 (n_93_148), .C2 (n_90_150) );
AOI211_X1 g_101_148 (.ZN (n_101_148), .A (n_99_148), .B (n_96_146), .C1 (n_94_150), .C2 (n_91_148) );
AOI211_X1 g_102_150 (.ZN (n_102_150), .A (n_100_146), .B (n_97_148), .C1 (n_95_148), .C2 (n_92_146) );
AOI211_X1 g_103_148 (.ZN (n_103_148), .A (n_101_148), .B (n_98_150), .C1 (n_96_146), .C2 (n_93_148) );
AOI211_X1 g_104_146 (.ZN (n_104_146), .A (n_102_150), .B (n_99_148), .C1 (n_97_148), .C2 (n_94_150) );
AOI211_X1 g_105_148 (.ZN (n_105_148), .A (n_103_148), .B (n_100_146), .C1 (n_98_150), .C2 (n_95_148) );
AOI211_X1 g_106_150 (.ZN (n_106_150), .A (n_104_146), .B (n_101_148), .C1 (n_99_148), .C2 (n_96_146) );
AOI211_X1 g_107_148 (.ZN (n_107_148), .A (n_105_148), .B (n_102_150), .C1 (n_100_146), .C2 (n_97_148) );
AOI211_X1 g_108_146 (.ZN (n_108_146), .A (n_106_150), .B (n_103_148), .C1 (n_101_148), .C2 (n_98_150) );
AOI211_X1 g_109_148 (.ZN (n_109_148), .A (n_107_148), .B (n_104_146), .C1 (n_102_150), .C2 (n_99_148) );
AOI211_X1 g_110_150 (.ZN (n_110_150), .A (n_108_146), .B (n_105_148), .C1 (n_103_148), .C2 (n_100_146) );
AOI211_X1 g_111_148 (.ZN (n_111_148), .A (n_109_148), .B (n_106_150), .C1 (n_104_146), .C2 (n_101_148) );
AOI211_X1 g_112_146 (.ZN (n_112_146), .A (n_110_150), .B (n_107_148), .C1 (n_105_148), .C2 (n_102_150) );
AOI211_X1 g_113_148 (.ZN (n_113_148), .A (n_111_148), .B (n_108_146), .C1 (n_106_150), .C2 (n_103_148) );
AOI211_X1 g_114_150 (.ZN (n_114_150), .A (n_112_146), .B (n_109_148), .C1 (n_107_148), .C2 (n_104_146) );
AOI211_X1 g_115_148 (.ZN (n_115_148), .A (n_113_148), .B (n_110_150), .C1 (n_108_146), .C2 (n_105_148) );
AOI211_X1 g_116_146 (.ZN (n_116_146), .A (n_114_150), .B (n_111_148), .C1 (n_109_148), .C2 (n_106_150) );
AOI211_X1 g_117_148 (.ZN (n_117_148), .A (n_115_148), .B (n_112_146), .C1 (n_110_150), .C2 (n_107_148) );
AOI211_X1 g_118_150 (.ZN (n_118_150), .A (n_116_146), .B (n_113_148), .C1 (n_111_148), .C2 (n_108_146) );
AOI211_X1 g_119_148 (.ZN (n_119_148), .A (n_117_148), .B (n_114_150), .C1 (n_112_146), .C2 (n_109_148) );
AOI211_X1 g_120_146 (.ZN (n_120_146), .A (n_118_150), .B (n_115_148), .C1 (n_113_148), .C2 (n_110_150) );
AOI211_X1 g_121_148 (.ZN (n_121_148), .A (n_119_148), .B (n_116_146), .C1 (n_114_150), .C2 (n_111_148) );
AOI211_X1 g_122_150 (.ZN (n_122_150), .A (n_120_146), .B (n_117_148), .C1 (n_115_148), .C2 (n_112_146) );
AOI211_X1 g_123_148 (.ZN (n_123_148), .A (n_121_148), .B (n_118_150), .C1 (n_116_146), .C2 (n_113_148) );
AOI211_X1 g_124_146 (.ZN (n_124_146), .A (n_122_150), .B (n_119_148), .C1 (n_117_148), .C2 (n_114_150) );
AOI211_X1 g_125_148 (.ZN (n_125_148), .A (n_123_148), .B (n_120_146), .C1 (n_118_150), .C2 (n_115_148) );
AOI211_X1 g_126_150 (.ZN (n_126_150), .A (n_124_146), .B (n_121_148), .C1 (n_119_148), .C2 (n_116_146) );
AOI211_X1 g_127_148 (.ZN (n_127_148), .A (n_125_148), .B (n_122_150), .C1 (n_120_146), .C2 (n_117_148) );
AOI211_X1 g_128_146 (.ZN (n_128_146), .A (n_126_150), .B (n_123_148), .C1 (n_121_148), .C2 (n_118_150) );
AOI211_X1 g_129_148 (.ZN (n_129_148), .A (n_127_148), .B (n_124_146), .C1 (n_122_150), .C2 (n_119_148) );
AOI211_X1 g_130_150 (.ZN (n_130_150), .A (n_128_146), .B (n_125_148), .C1 (n_123_148), .C2 (n_120_146) );
AOI211_X1 g_131_148 (.ZN (n_131_148), .A (n_129_148), .B (n_126_150), .C1 (n_124_146), .C2 (n_121_148) );
AOI211_X1 g_132_146 (.ZN (n_132_146), .A (n_130_150), .B (n_127_148), .C1 (n_125_148), .C2 (n_122_150) );
AOI211_X1 g_133_148 (.ZN (n_133_148), .A (n_131_148), .B (n_128_146), .C1 (n_126_150), .C2 (n_123_148) );
AOI211_X1 g_134_150 (.ZN (n_134_150), .A (n_132_146), .B (n_129_148), .C1 (n_127_148), .C2 (n_124_146) );
AOI211_X1 g_135_148 (.ZN (n_135_148), .A (n_133_148), .B (n_130_150), .C1 (n_128_146), .C2 (n_125_148) );
AOI211_X1 g_136_146 (.ZN (n_136_146), .A (n_134_150), .B (n_131_148), .C1 (n_129_148), .C2 (n_126_150) );
AOI211_X1 g_137_148 (.ZN (n_137_148), .A (n_135_148), .B (n_132_146), .C1 (n_130_150), .C2 (n_127_148) );
AOI211_X1 g_138_150 (.ZN (n_138_150), .A (n_136_146), .B (n_133_148), .C1 (n_131_148), .C2 (n_128_146) );
AOI211_X1 g_139_148 (.ZN (n_139_148), .A (n_137_148), .B (n_134_150), .C1 (n_132_146), .C2 (n_129_148) );
AOI211_X1 g_141_147 (.ZN (n_141_147), .A (n_138_150), .B (n_135_148), .C1 (n_133_148), .C2 (n_130_150) );
AOI211_X1 g_140_149 (.ZN (n_140_149), .A (n_139_148), .B (n_136_146), .C1 (n_134_150), .C2 (n_131_148) );
AOI211_X1 g_142_148 (.ZN (n_142_148), .A (n_141_147), .B (n_137_148), .C1 (n_135_148), .C2 (n_132_146) );
AOI211_X1 g_144_147 (.ZN (n_144_147), .A (n_140_149), .B (n_138_150), .C1 (n_136_146), .C2 (n_133_148) );
AOI211_X1 g_145_145 (.ZN (n_145_145), .A (n_142_148), .B (n_139_148), .C1 (n_137_148), .C2 (n_134_150) );
AOI211_X1 g_143_146 (.ZN (n_143_146), .A (n_144_147), .B (n_141_147), .C1 (n_138_150), .C2 (n_135_148) );
AOI211_X1 g_144_144 (.ZN (n_144_144), .A (n_145_145), .B (n_140_149), .C1 (n_139_148), .C2 (n_136_146) );
AOI211_X1 g_142_145 (.ZN (n_142_145), .A (n_143_146), .B (n_142_148), .C1 (n_141_147), .C2 (n_137_148) );
AOI211_X1 g_143_143 (.ZN (n_143_143), .A (n_144_144), .B (n_144_147), .C1 (n_140_149), .C2 (n_138_150) );
AOI211_X1 g_145_142 (.ZN (n_145_142), .A (n_142_145), .B (n_145_145), .C1 (n_142_148), .C2 (n_139_148) );
AOI211_X1 g_146_144 (.ZN (n_146_144), .A (n_143_143), .B (n_143_146), .C1 (n_144_147), .C2 (n_141_147) );
AOI211_X1 g_147_142 (.ZN (n_147_142), .A (n_145_142), .B (n_144_144), .C1 (n_145_145), .C2 (n_140_149) );
AOI211_X1 g_146_140 (.ZN (n_146_140), .A (n_146_144), .B (n_142_145), .C1 (n_143_146), .C2 (n_142_148) );
AOI211_X1 g_144_141 (.ZN (n_144_141), .A (n_147_142), .B (n_143_143), .C1 (n_144_144), .C2 (n_144_147) );
AOI211_X1 g_145_143 (.ZN (n_145_143), .A (n_146_140), .B (n_145_142), .C1 (n_142_145), .C2 (n_145_145) );
AOI211_X1 g_144_145 (.ZN (n_144_145), .A (n_144_141), .B (n_146_144), .C1 (n_143_143), .C2 (n_143_146) );
AOI211_X1 g_142_146 (.ZN (n_142_146), .A (n_145_143), .B (n_147_142), .C1 (n_145_142), .C2 (n_144_144) );
AOI211_X1 g_143_144 (.ZN (n_143_144), .A (n_144_145), .B (n_146_140), .C1 (n_146_144), .C2 (n_142_145) );
AOI211_X1 g_141_145 (.ZN (n_141_145), .A (n_142_146), .B (n_144_141), .C1 (n_147_142), .C2 (n_143_143) );
AOI211_X1 g_140_147 (.ZN (n_140_147), .A (n_143_144), .B (n_145_143), .C1 (n_146_140), .C2 (n_145_142) );
AOI211_X1 g_138_148 (.ZN (n_138_148), .A (n_141_145), .B (n_144_145), .C1 (n_144_141), .C2 (n_146_144) );
AOI211_X1 g_136_149 (.ZN (n_136_149), .A (n_140_147), .B (n_142_146), .C1 (n_145_143), .C2 (n_147_142) );
AOI211_X1 g_137_147 (.ZN (n_137_147), .A (n_138_148), .B (n_143_144), .C1 (n_144_145), .C2 (n_146_140) );
AOI211_X1 g_139_146 (.ZN (n_139_146), .A (n_136_149), .B (n_141_145), .C1 (n_142_146), .C2 (n_144_141) );
AOI211_X1 g_140_144 (.ZN (n_140_144), .A (n_137_147), .B (n_140_147), .C1 (n_143_144), .C2 (n_145_143) );
AOI211_X1 g_142_143 (.ZN (n_142_143), .A (n_139_146), .B (n_138_148), .C1 (n_141_145), .C2 (n_144_145) );
AOI211_X1 g_143_145 (.ZN (n_143_145), .A (n_140_144), .B (n_136_149), .C1 (n_140_147), .C2 (n_142_146) );
AOI211_X1 g_141_146 (.ZN (n_141_146), .A (n_142_143), .B (n_137_147), .C1 (n_138_148), .C2 (n_143_144) );
AOI211_X1 g_139_147 (.ZN (n_139_147), .A (n_143_145), .B (n_139_146), .C1 (n_136_149), .C2 (n_141_145) );
AOI211_X1 g_138_145 (.ZN (n_138_145), .A (n_141_146), .B (n_140_144), .C1 (n_137_147), .C2 (n_140_147) );
AOI211_X1 g_139_143 (.ZN (n_139_143), .A (n_139_147), .B (n_142_143), .C1 (n_139_146), .C2 (n_138_148) );
AOI211_X1 g_141_144 (.ZN (n_141_144), .A (n_138_145), .B (n_143_145), .C1 (n_140_144), .C2 (n_136_149) );
AOI211_X1 g_139_145 (.ZN (n_139_145), .A (n_139_143), .B (n_141_146), .C1 (n_142_143), .C2 (n_137_147) );
AOI211_X1 g_137_146 (.ZN (n_137_146), .A (n_141_144), .B (n_139_147), .C1 (n_143_145), .C2 (n_139_146) );
AOI211_X1 g_135_147 (.ZN (n_135_147), .A (n_139_145), .B (n_138_145), .C1 (n_141_146), .C2 (n_140_144) );
AOI211_X1 g_134_145 (.ZN (n_134_145), .A (n_137_146), .B (n_139_143), .C1 (n_139_147), .C2 (n_142_143) );
AOI211_X1 g_133_147 (.ZN (n_133_147), .A (n_135_147), .B (n_141_144), .C1 (n_138_145), .C2 (n_143_145) );
AOI211_X1 g_132_149 (.ZN (n_132_149), .A (n_134_145), .B (n_139_145), .C1 (n_139_143), .C2 (n_141_146) );
AOI211_X1 g_134_148 (.ZN (n_134_148), .A (n_133_147), .B (n_137_146), .C1 (n_141_144), .C2 (n_139_147) );
AOI211_X1 g_136_147 (.ZN (n_136_147), .A (n_132_149), .B (n_135_147), .C1 (n_139_145), .C2 (n_138_145) );
AOI211_X1 g_138_146 (.ZN (n_138_146), .A (n_134_148), .B (n_134_145), .C1 (n_137_146), .C2 (n_139_143) );
AOI211_X1 g_140_145 (.ZN (n_140_145), .A (n_136_147), .B (n_133_147), .C1 (n_135_147), .C2 (n_141_144) );
AOI211_X1 g_142_144 (.ZN (n_142_144), .A (n_138_146), .B (n_132_149), .C1 (n_134_145), .C2 (n_139_145) );
AOI211_X1 g_144_143 (.ZN (n_144_143), .A (n_140_145), .B (n_134_148), .C1 (n_133_147), .C2 (n_137_146) );
AOI211_X1 g_145_141 (.ZN (n_145_141), .A (n_142_144), .B (n_136_147), .C1 (n_132_149), .C2 (n_135_147) );
AOI211_X1 g_146_139 (.ZN (n_146_139), .A (n_144_143), .B (n_138_146), .C1 (n_134_148), .C2 (n_134_145) );
AOI211_X1 g_147_137 (.ZN (n_147_137), .A (n_145_141), .B (n_140_145), .C1 (n_136_147), .C2 (n_133_147) );
AOI211_X1 g_148_135 (.ZN (n_148_135), .A (n_146_139), .B (n_142_144), .C1 (n_138_146), .C2 (n_132_149) );
AOI211_X1 g_146_136 (.ZN (n_146_136), .A (n_147_137), .B (n_144_143), .C1 (n_140_145), .C2 (n_134_148) );
AOI211_X1 g_145_138 (.ZN (n_145_138), .A (n_148_135), .B (n_145_141), .C1 (n_142_144), .C2 (n_136_147) );
AOI211_X1 g_143_139 (.ZN (n_143_139), .A (n_146_136), .B (n_146_139), .C1 (n_144_143), .C2 (n_138_146) );
AOI211_X1 g_142_141 (.ZN (n_142_141), .A (n_145_138), .B (n_147_137), .C1 (n_145_141), .C2 (n_140_145) );
AOI211_X1 g_144_140 (.ZN (n_144_140), .A (n_143_139), .B (n_148_135), .C1 (n_146_139), .C2 (n_142_144) );
AOI211_X1 g_143_142 (.ZN (n_143_142), .A (n_142_141), .B (n_146_136), .C1 (n_147_137), .C2 (n_144_143) );
AOI211_X1 g_141_143 (.ZN (n_141_143), .A (n_144_140), .B (n_145_138), .C1 (n_148_135), .C2 (n_145_141) );
AOI211_X1 g_139_144 (.ZN (n_139_144), .A (n_143_142), .B (n_143_139), .C1 (n_146_136), .C2 (n_146_139) );
AOI211_X1 g_140_142 (.ZN (n_140_142), .A (n_141_143), .B (n_142_141), .C1 (n_145_138), .C2 (n_147_137) );
AOI211_X1 g_138_143 (.ZN (n_138_143), .A (n_139_144), .B (n_144_140), .C1 (n_143_139), .C2 (n_148_135) );
AOI211_X1 g_137_145 (.ZN (n_137_145), .A (n_140_142), .B (n_143_142), .C1 (n_142_141), .C2 (n_146_136) );
AOI211_X1 g_135_146 (.ZN (n_135_146), .A (n_138_143), .B (n_141_143), .C1 (n_144_140), .C2 (n_145_138) );
AOI211_X1 g_136_144 (.ZN (n_136_144), .A (n_137_145), .B (n_139_144), .C1 (n_143_142), .C2 (n_143_139) );
AOI211_X1 g_137_142 (.ZN (n_137_142), .A (n_135_146), .B (n_140_142), .C1 (n_141_143), .C2 (n_142_141) );
AOI211_X1 g_138_144 (.ZN (n_138_144), .A (n_136_144), .B (n_138_143), .C1 (n_139_144), .C2 (n_144_140) );
AOI211_X1 g_140_143 (.ZN (n_140_143), .A (n_137_142), .B (n_137_145), .C1 (n_140_142), .C2 (n_143_142) );
AOI211_X1 g_142_142 (.ZN (n_142_142), .A (n_138_144), .B (n_135_146), .C1 (n_138_143), .C2 (n_141_143) );
AOI211_X1 g_143_140 (.ZN (n_143_140), .A (n_140_143), .B (n_136_144), .C1 (n_137_145), .C2 (n_139_144) );
AOI211_X1 g_144_138 (.ZN (n_144_138), .A (n_142_142), .B (n_137_142), .C1 (n_135_146), .C2 (n_140_142) );
AOI211_X1 g_145_136 (.ZN (n_145_136), .A (n_143_140), .B (n_138_144), .C1 (n_136_144), .C2 (n_138_143) );
AOI211_X1 g_146_134 (.ZN (n_146_134), .A (n_144_138), .B (n_140_143), .C1 (n_137_142), .C2 (n_137_145) );
AOI211_X1 g_144_133 (.ZN (n_144_133), .A (n_145_136), .B (n_142_142), .C1 (n_138_144), .C2 (n_135_146) );
AOI211_X1 g_146_132 (.ZN (n_146_132), .A (n_146_134), .B (n_143_140), .C1 (n_140_143), .C2 (n_136_144) );
AOI211_X1 g_148_131 (.ZN (n_148_131), .A (n_144_133), .B (n_144_138), .C1 (n_142_142), .C2 (n_137_142) );
AOI211_X1 g_146_130 (.ZN (n_146_130), .A (n_146_132), .B (n_145_136), .C1 (n_143_140), .C2 (n_138_144) );
AOI211_X1 g_144_129 (.ZN (n_144_129), .A (n_148_131), .B (n_146_134), .C1 (n_144_138), .C2 (n_140_143) );
AOI211_X1 g_146_128 (.ZN (n_146_128), .A (n_146_130), .B (n_144_133), .C1 (n_145_136), .C2 (n_142_142) );
AOI211_X1 g_148_127 (.ZN (n_148_127), .A (n_144_129), .B (n_146_132), .C1 (n_146_134), .C2 (n_143_140) );
AOI211_X1 g_146_126 (.ZN (n_146_126), .A (n_146_128), .B (n_148_131), .C1 (n_144_133), .C2 (n_144_138) );
AOI211_X1 g_144_125 (.ZN (n_144_125), .A (n_148_127), .B (n_146_130), .C1 (n_146_132), .C2 (n_145_136) );
AOI211_X1 g_146_124 (.ZN (n_146_124), .A (n_146_126), .B (n_144_129), .C1 (n_148_131), .C2 (n_146_134) );
AOI211_X1 g_148_123 (.ZN (n_148_123), .A (n_144_125), .B (n_146_128), .C1 (n_146_130), .C2 (n_144_133) );
AOI211_X1 g_147_121 (.ZN (n_147_121), .A (n_146_124), .B (n_148_127), .C1 (n_144_129), .C2 (n_146_132) );
AOI211_X1 g_146_119 (.ZN (n_146_119), .A (n_148_123), .B (n_146_126), .C1 (n_146_128), .C2 (n_148_131) );
AOI211_X1 g_144_118 (.ZN (n_144_118), .A (n_147_121), .B (n_144_125), .C1 (n_148_127), .C2 (n_146_130) );
AOI211_X1 g_143_120 (.ZN (n_143_120), .A (n_146_119), .B (n_146_124), .C1 (n_146_126), .C2 (n_144_129) );
AOI211_X1 g_145_121 (.ZN (n_145_121), .A (n_144_118), .B (n_148_123), .C1 (n_144_125), .C2 (n_146_128) );
AOI211_X1 g_144_119 (.ZN (n_144_119), .A (n_143_120), .B (n_147_121), .C1 (n_146_124), .C2 (n_148_127) );
AOI211_X1 g_143_117 (.ZN (n_143_117), .A (n_145_121), .B (n_146_119), .C1 (n_148_123), .C2 (n_146_126) );
AOI211_X1 g_145_118 (.ZN (n_145_118), .A (n_144_119), .B (n_144_118), .C1 (n_147_121), .C2 (n_144_125) );
AOI211_X1 g_146_120 (.ZN (n_146_120), .A (n_143_117), .B (n_143_120), .C1 (n_146_119), .C2 (n_146_124) );
AOI211_X1 g_145_122 (.ZN (n_145_122), .A (n_145_118), .B (n_145_121), .C1 (n_144_118), .C2 (n_148_123) );
AOI211_X1 g_144_120 (.ZN (n_144_120), .A (n_146_120), .B (n_144_119), .C1 (n_143_120), .C2 (n_147_121) );
AOI211_X1 g_142_119 (.ZN (n_142_119), .A (n_145_122), .B (n_143_117), .C1 (n_145_121), .C2 (n_146_119) );
AOI211_X1 g_140_120 (.ZN (n_140_120), .A (n_144_120), .B (n_145_118), .C1 (n_144_119), .C2 (n_144_118) );
AOI211_X1 g_141_118 (.ZN (n_141_118), .A (n_142_119), .B (n_146_120), .C1 (n_143_117), .C2 (n_143_120) );
AOI211_X1 g_139_119 (.ZN (n_139_119), .A (n_140_120), .B (n_145_122), .C1 (n_145_118), .C2 (n_145_121) );
AOI211_X1 g_138_121 (.ZN (n_138_121), .A (n_141_118), .B (n_144_120), .C1 (n_146_120), .C2 (n_144_119) );
AOI211_X1 g_136_122 (.ZN (n_136_122), .A (n_139_119), .B (n_142_119), .C1 (n_145_122), .C2 (n_143_117) );
AOI211_X1 g_134_123 (.ZN (n_134_123), .A (n_138_121), .B (n_140_120), .C1 (n_144_120), .C2 (n_145_118) );
AOI211_X1 g_132_124 (.ZN (n_132_124), .A (n_136_122), .B (n_141_118), .C1 (n_142_119), .C2 (n_146_120) );
AOI211_X1 g_130_125 (.ZN (n_130_125), .A (n_134_123), .B (n_139_119), .C1 (n_140_120), .C2 (n_145_122) );
AOI211_X1 g_128_126 (.ZN (n_128_126), .A (n_132_124), .B (n_138_121), .C1 (n_141_118), .C2 (n_144_120) );
AOI211_X1 g_129_124 (.ZN (n_129_124), .A (n_130_125), .B (n_136_122), .C1 (n_139_119), .C2 (n_142_119) );
AOI211_X1 g_127_125 (.ZN (n_127_125), .A (n_128_126), .B (n_134_123), .C1 (n_138_121), .C2 (n_140_120) );
AOI211_X1 g_125_126 (.ZN (n_125_126), .A (n_129_124), .B (n_132_124), .C1 (n_136_122), .C2 (n_141_118) );
AOI211_X1 g_123_127 (.ZN (n_123_127), .A (n_127_125), .B (n_130_125), .C1 (n_134_123), .C2 (n_139_119) );
AOI211_X1 g_121_128 (.ZN (n_121_128), .A (n_125_126), .B (n_128_126), .C1 (n_132_124), .C2 (n_138_121) );
AOI211_X1 g_119_129 (.ZN (n_119_129), .A (n_123_127), .B (n_129_124), .C1 (n_130_125), .C2 (n_136_122) );
AOI211_X1 g_117_130 (.ZN (n_117_130), .A (n_121_128), .B (n_127_125), .C1 (n_128_126), .C2 (n_134_123) );
AOI211_X1 g_116_128 (.ZN (n_116_128), .A (n_119_129), .B (n_125_126), .C1 (n_129_124), .C2 (n_132_124) );
AOI211_X1 g_114_129 (.ZN (n_114_129), .A (n_117_130), .B (n_123_127), .C1 (n_127_125), .C2 (n_130_125) );
AOI211_X1 g_112_130 (.ZN (n_112_130), .A (n_116_128), .B (n_121_128), .C1 (n_125_126), .C2 (n_128_126) );
AOI211_X1 g_114_131 (.ZN (n_114_131), .A (n_114_129), .B (n_119_129), .C1 (n_123_127), .C2 (n_129_124) );
AOI211_X1 g_116_130 (.ZN (n_116_130), .A (n_112_130), .B (n_117_130), .C1 (n_121_128), .C2 (n_127_125) );
AOI211_X1 g_118_129 (.ZN (n_118_129), .A (n_114_131), .B (n_116_128), .C1 (n_119_129), .C2 (n_125_126) );
AOI211_X1 g_117_131 (.ZN (n_117_131), .A (n_116_130), .B (n_114_129), .C1 (n_117_130), .C2 (n_123_127) );
AOI211_X1 g_115_130 (.ZN (n_115_130), .A (n_118_129), .B (n_112_130), .C1 (n_116_128), .C2 (n_121_128) );
AOI211_X1 g_117_129 (.ZN (n_117_129), .A (n_117_131), .B (n_114_131), .C1 (n_114_129), .C2 (n_119_129) );
AOI211_X1 g_119_128 (.ZN (n_119_128), .A (n_115_130), .B (n_116_130), .C1 (n_112_130), .C2 (n_117_130) );
AOI211_X1 g_121_127 (.ZN (n_121_127), .A (n_117_129), .B (n_118_129), .C1 (n_114_131), .C2 (n_116_128) );
AOI211_X1 g_120_129 (.ZN (n_120_129), .A (n_119_128), .B (n_117_131), .C1 (n_116_130), .C2 (n_114_129) );
AOI211_X1 g_122_128 (.ZN (n_122_128), .A (n_121_127), .B (n_115_130), .C1 (n_118_129), .C2 (n_112_130) );
AOI211_X1 g_124_127 (.ZN (n_124_127), .A (n_120_129), .B (n_117_129), .C1 (n_117_131), .C2 (n_114_131) );
AOI211_X1 g_126_126 (.ZN (n_126_126), .A (n_122_128), .B (n_119_128), .C1 (n_115_130), .C2 (n_116_130) );
AOI211_X1 g_125_128 (.ZN (n_125_128), .A (n_124_127), .B (n_121_127), .C1 (n_117_129), .C2 (n_118_129) );
AOI211_X1 g_124_126 (.ZN (n_124_126), .A (n_126_126), .B (n_120_129), .C1 (n_119_128), .C2 (n_117_131) );
AOI211_X1 g_122_127 (.ZN (n_122_127), .A (n_125_128), .B (n_122_128), .C1 (n_121_127), .C2 (n_115_130) );
AOI211_X1 g_123_129 (.ZN (n_123_129), .A (n_124_126), .B (n_124_127), .C1 (n_120_129), .C2 (n_117_129) );
AOI211_X1 g_121_130 (.ZN (n_121_130), .A (n_122_127), .B (n_126_126), .C1 (n_122_128), .C2 (n_119_128) );
AOI211_X1 g_119_131 (.ZN (n_119_131), .A (n_123_129), .B (n_125_128), .C1 (n_124_127), .C2 (n_121_127) );
AOI211_X1 g_117_132 (.ZN (n_117_132), .A (n_121_130), .B (n_124_126), .C1 (n_126_126), .C2 (n_120_129) );
AOI211_X1 g_118_130 (.ZN (n_118_130), .A (n_119_131), .B (n_122_127), .C1 (n_125_128), .C2 (n_122_128) );
AOI211_X1 g_116_131 (.ZN (n_116_131), .A (n_117_132), .B (n_123_129), .C1 (n_124_126), .C2 (n_124_127) );
AOI211_X1 g_114_132 (.ZN (n_114_132), .A (n_118_130), .B (n_121_130), .C1 (n_122_127), .C2 (n_126_126) );
AOI211_X1 g_112_133 (.ZN (n_112_133), .A (n_116_131), .B (n_119_131), .C1 (n_123_129), .C2 (n_125_128) );
AOI211_X1 g_113_131 (.ZN (n_113_131), .A (n_114_132), .B (n_117_132), .C1 (n_121_130), .C2 (n_124_126) );
AOI211_X1 g_111_132 (.ZN (n_111_132), .A (n_112_133), .B (n_118_130), .C1 (n_119_131), .C2 (n_122_127) );
AOI211_X1 g_109_133 (.ZN (n_109_133), .A (n_113_131), .B (n_116_131), .C1 (n_117_132), .C2 (n_123_129) );
AOI211_X1 g_111_134 (.ZN (n_111_134), .A (n_111_132), .B (n_114_132), .C1 (n_118_130), .C2 (n_121_130) );
AOI211_X1 g_113_133 (.ZN (n_113_133), .A (n_109_133), .B (n_112_133), .C1 (n_116_131), .C2 (n_119_131) );
AOI211_X1 g_115_132 (.ZN (n_115_132), .A (n_111_134), .B (n_113_131), .C1 (n_114_132), .C2 (n_117_132) );
AOI211_X1 g_114_134 (.ZN (n_114_134), .A (n_113_133), .B (n_111_132), .C1 (n_112_133), .C2 (n_118_130) );
AOI211_X1 g_113_132 (.ZN (n_113_132), .A (n_115_132), .B (n_109_133), .C1 (n_113_131), .C2 (n_116_131) );
AOI211_X1 g_115_131 (.ZN (n_115_131), .A (n_114_134), .B (n_111_134), .C1 (n_111_132), .C2 (n_114_132) );
AOI211_X1 g_116_133 (.ZN (n_116_133), .A (n_113_132), .B (n_113_133), .C1 (n_109_133), .C2 (n_112_133) );
AOI211_X1 g_118_132 (.ZN (n_118_132), .A (n_115_131), .B (n_115_132), .C1 (n_111_134), .C2 (n_113_131) );
AOI211_X1 g_119_130 (.ZN (n_119_130), .A (n_116_133), .B (n_114_134), .C1 (n_113_133), .C2 (n_111_132) );
AOI211_X1 g_121_129 (.ZN (n_121_129), .A (n_118_132), .B (n_113_132), .C1 (n_115_132), .C2 (n_109_133) );
AOI211_X1 g_123_128 (.ZN (n_123_128), .A (n_119_130), .B (n_115_131), .C1 (n_114_134), .C2 (n_111_134) );
AOI211_X1 g_125_127 (.ZN (n_125_127), .A (n_121_129), .B (n_116_133), .C1 (n_113_132), .C2 (n_113_133) );
AOI211_X1 g_127_126 (.ZN (n_127_126), .A (n_123_128), .B (n_118_132), .C1 (n_115_131), .C2 (n_115_132) );
AOI211_X1 g_129_125 (.ZN (n_129_125), .A (n_125_127), .B (n_119_130), .C1 (n_116_133), .C2 (n_114_134) );
AOI211_X1 g_131_124 (.ZN (n_131_124), .A (n_127_126), .B (n_121_129), .C1 (n_118_132), .C2 (n_113_132) );
AOI211_X1 g_133_123 (.ZN (n_133_123), .A (n_129_125), .B (n_123_128), .C1 (n_119_130), .C2 (n_115_131) );
AOI211_X1 g_135_122 (.ZN (n_135_122), .A (n_131_124), .B (n_125_127), .C1 (n_121_129), .C2 (n_116_133) );
AOI211_X1 g_137_121 (.ZN (n_137_121), .A (n_133_123), .B (n_127_126), .C1 (n_123_128), .C2 (n_118_132) );
AOI211_X1 g_139_120 (.ZN (n_139_120), .A (n_135_122), .B (n_129_125), .C1 (n_125_127), .C2 (n_119_130) );
AOI211_X1 g_141_121 (.ZN (n_141_121), .A (n_137_121), .B (n_131_124), .C1 (n_127_126), .C2 (n_121_129) );
AOI211_X1 g_139_122 (.ZN (n_139_122), .A (n_139_120), .B (n_133_123), .C1 (n_129_125), .C2 (n_123_128) );
AOI211_X1 g_137_123 (.ZN (n_137_123), .A (n_141_121), .B (n_135_122), .C1 (n_131_124), .C2 (n_125_127) );
AOI211_X1 g_135_124 (.ZN (n_135_124), .A (n_139_122), .B (n_137_121), .C1 (n_133_123), .C2 (n_127_126) );
AOI211_X1 g_133_125 (.ZN (n_133_125), .A (n_137_123), .B (n_139_120), .C1 (n_135_122), .C2 (n_129_125) );
AOI211_X1 g_131_126 (.ZN (n_131_126), .A (n_135_124), .B (n_141_121), .C1 (n_137_121), .C2 (n_131_124) );
AOI211_X1 g_129_127 (.ZN (n_129_127), .A (n_133_125), .B (n_139_122), .C1 (n_139_120), .C2 (n_133_123) );
AOI211_X1 g_127_128 (.ZN (n_127_128), .A (n_131_126), .B (n_137_123), .C1 (n_141_121), .C2 (n_135_122) );
AOI211_X1 g_125_129 (.ZN (n_125_129), .A (n_129_127), .B (n_135_124), .C1 (n_139_122), .C2 (n_137_121) );
AOI211_X1 g_126_127 (.ZN (n_126_127), .A (n_127_128), .B (n_133_125), .C1 (n_137_123), .C2 (n_139_120) );
AOI211_X1 g_124_128 (.ZN (n_124_128), .A (n_125_129), .B (n_131_126), .C1 (n_135_124), .C2 (n_141_121) );
AOI211_X1 g_122_129 (.ZN (n_122_129), .A (n_126_127), .B (n_129_127), .C1 (n_133_125), .C2 (n_139_122) );
AOI211_X1 g_120_130 (.ZN (n_120_130), .A (n_124_128), .B (n_127_128), .C1 (n_131_126), .C2 (n_137_123) );
AOI211_X1 g_118_131 (.ZN (n_118_131), .A (n_122_129), .B (n_125_129), .C1 (n_129_127), .C2 (n_135_124) );
AOI211_X1 g_116_132 (.ZN (n_116_132), .A (n_120_130), .B (n_126_127), .C1 (n_127_128), .C2 (n_133_125) );
AOI211_X1 g_114_133 (.ZN (n_114_133), .A (n_118_131), .B (n_124_128), .C1 (n_125_129), .C2 (n_131_126) );
AOI211_X1 g_112_134 (.ZN (n_112_134), .A (n_116_132), .B (n_122_129), .C1 (n_126_127), .C2 (n_129_127) );
AOI211_X1 g_110_135 (.ZN (n_110_135), .A (n_114_133), .B (n_120_130), .C1 (n_124_128), .C2 (n_127_128) );
AOI211_X1 g_111_133 (.ZN (n_111_133), .A (n_112_134), .B (n_118_131), .C1 (n_122_129), .C2 (n_125_129) );
AOI211_X1 g_109_134 (.ZN (n_109_134), .A (n_110_135), .B (n_116_132), .C1 (n_120_130), .C2 (n_126_127) );
AOI211_X1 g_107_135 (.ZN (n_107_135), .A (n_111_133), .B (n_114_133), .C1 (n_118_131), .C2 (n_124_128) );
AOI211_X1 g_106_137 (.ZN (n_106_137), .A (n_109_134), .B (n_112_134), .C1 (n_116_132), .C2 (n_122_129) );
AOI211_X1 g_108_136 (.ZN (n_108_136), .A (n_107_135), .B (n_110_135), .C1 (n_114_133), .C2 (n_120_130) );
AOI211_X1 g_107_138 (.ZN (n_107_138), .A (n_106_137), .B (n_111_133), .C1 (n_112_134), .C2 (n_118_131) );
AOI211_X1 g_106_136 (.ZN (n_106_136), .A (n_108_136), .B (n_109_134), .C1 (n_110_135), .C2 (n_116_132) );
AOI211_X1 g_108_135 (.ZN (n_108_135), .A (n_107_138), .B (n_107_135), .C1 (n_111_133), .C2 (n_114_133) );
AOI211_X1 g_110_134 (.ZN (n_110_134), .A (n_106_136), .B (n_106_137), .C1 (n_109_134), .C2 (n_112_134) );
AOI211_X1 g_112_135 (.ZN (n_112_135), .A (n_108_135), .B (n_108_136), .C1 (n_107_135), .C2 (n_110_135) );
AOI211_X1 g_110_136 (.ZN (n_110_136), .A (n_110_134), .B (n_107_138), .C1 (n_106_137), .C2 (n_111_133) );
AOI211_X1 g_108_137 (.ZN (n_108_137), .A (n_112_135), .B (n_106_136), .C1 (n_108_136), .C2 (n_109_134) );
AOI211_X1 g_106_138 (.ZN (n_106_138), .A (n_110_136), .B (n_108_135), .C1 (n_107_138), .C2 (n_107_135) );
AOI211_X1 g_104_137 (.ZN (n_104_137), .A (n_108_137), .B (n_110_134), .C1 (n_106_136), .C2 (n_106_137) );
AOI211_X1 g_102_138 (.ZN (n_102_138), .A (n_106_138), .B (n_112_135), .C1 (n_108_135), .C2 (n_108_136) );
AOI211_X1 g_100_139 (.ZN (n_100_139), .A (n_104_137), .B (n_110_136), .C1 (n_110_134), .C2 (n_107_138) );
AOI211_X1 g_98_140 (.ZN (n_98_140), .A (n_102_138), .B (n_108_137), .C1 (n_112_135), .C2 (n_106_136) );
AOI211_X1 g_96_141 (.ZN (n_96_141), .A (n_100_139), .B (n_106_138), .C1 (n_110_136), .C2 (n_108_135) );
AOI211_X1 g_94_142 (.ZN (n_94_142), .A (n_98_140), .B (n_104_137), .C1 (n_108_137), .C2 (n_110_134) );
AOI211_X1 g_92_143 (.ZN (n_92_143), .A (n_96_141), .B (n_102_138), .C1 (n_106_138), .C2 (n_112_135) );
AOI211_X1 g_90_144 (.ZN (n_90_144), .A (n_94_142), .B (n_100_139), .C1 (n_104_137), .C2 (n_110_136) );
AOI211_X1 g_91_142 (.ZN (n_91_142), .A (n_92_143), .B (n_98_140), .C1 (n_102_138), .C2 (n_108_137) );
AOI211_X1 g_89_143 (.ZN (n_89_143), .A (n_90_144), .B (n_96_141), .C1 (n_100_139), .C2 (n_106_138) );
AOI211_X1 g_87_144 (.ZN (n_87_144), .A (n_91_142), .B (n_94_142), .C1 (n_98_140), .C2 (n_104_137) );
AOI211_X1 g_86_146 (.ZN (n_86_146), .A (n_89_143), .B (n_92_143), .C1 (n_96_141), .C2 (n_102_138) );
AOI211_X1 g_84_145 (.ZN (n_84_145), .A (n_87_144), .B (n_90_144), .C1 (n_94_142), .C2 (n_100_139) );
AOI211_X1 g_85_147 (.ZN (n_85_147), .A (n_86_146), .B (n_91_142), .C1 (n_92_143), .C2 (n_98_140) );
AOI211_X1 g_87_148 (.ZN (n_87_148), .A (n_84_145), .B (n_89_143), .C1 (n_90_144), .C2 (n_96_141) );
AOI211_X1 g_89_147 (.ZN (n_89_147), .A (n_85_147), .B (n_87_144), .C1 (n_91_142), .C2 (n_94_142) );
AOI211_X1 g_87_146 (.ZN (n_87_146), .A (n_87_148), .B (n_86_146), .C1 (n_89_143), .C2 (n_92_143) );
AOI211_X1 g_89_145 (.ZN (n_89_145), .A (n_89_147), .B (n_84_145), .C1 (n_87_144), .C2 (n_90_144) );
AOI211_X1 g_88_147 (.ZN (n_88_147), .A (n_87_146), .B (n_85_147), .C1 (n_86_146), .C2 (n_91_142) );
AOI211_X1 g_90_148 (.ZN (n_90_148), .A (n_89_145), .B (n_87_148), .C1 (n_84_145), .C2 (n_89_143) );
AOI211_X1 g_91_146 (.ZN (n_91_146), .A (n_88_147), .B (n_89_147), .C1 (n_85_147), .C2 (n_87_144) );
AOI211_X1 g_93_147 (.ZN (n_93_147), .A (n_90_148), .B (n_87_146), .C1 (n_87_148), .C2 (n_86_146) );
AOI211_X1 g_92_149 (.ZN (n_92_149), .A (n_91_146), .B (n_89_145), .C1 (n_89_147), .C2 (n_84_145) );
AOI211_X1 g_94_148 (.ZN (n_94_148), .A (n_93_147), .B (n_88_147), .C1 (n_87_146), .C2 (n_85_147) );
AOI211_X1 g_96_149 (.ZN (n_96_149), .A (n_92_149), .B (n_90_148), .C1 (n_89_145), .C2 (n_87_148) );
AOI211_X1 g_97_147 (.ZN (n_97_147), .A (n_94_148), .B (n_91_146), .C1 (n_88_147), .C2 (n_89_147) );
AOI211_X1 g_95_146 (.ZN (n_95_146), .A (n_96_149), .B (n_93_147), .C1 (n_90_148), .C2 (n_87_146) );
AOI211_X1 g_93_145 (.ZN (n_93_145), .A (n_97_147), .B (n_92_149), .C1 (n_91_146), .C2 (n_89_145) );
AOI211_X1 g_91_144 (.ZN (n_91_144), .A (n_95_146), .B (n_94_148), .C1 (n_93_147), .C2 (n_88_147) );
AOI211_X1 g_93_143 (.ZN (n_93_143), .A (n_93_145), .B (n_96_149), .C1 (n_92_149), .C2 (n_90_148) );
AOI211_X1 g_94_145 (.ZN (n_94_145), .A (n_91_144), .B (n_97_147), .C1 (n_94_148), .C2 (n_91_146) );
AOI211_X1 g_95_147 (.ZN (n_95_147), .A (n_93_143), .B (n_95_146), .C1 (n_96_149), .C2 (n_93_147) );
AOI211_X1 g_93_146 (.ZN (n_93_146), .A (n_94_145), .B (n_93_145), .C1 (n_97_147), .C2 (n_92_149) );
AOI211_X1 g_94_144 (.ZN (n_94_144), .A (n_95_147), .B (n_91_144), .C1 (n_95_146), .C2 (n_94_148) );
AOI211_X1 g_93_142 (.ZN (n_93_142), .A (n_93_146), .B (n_93_143), .C1 (n_93_145), .C2 (n_96_149) );
AOI211_X1 g_92_144 (.ZN (n_92_144), .A (n_94_144), .B (n_94_145), .C1 (n_91_144), .C2 (n_97_147) );
AOI211_X1 g_90_143 (.ZN (n_90_143), .A (n_93_142), .B (n_95_147), .C1 (n_93_143), .C2 (n_95_146) );
AOI211_X1 g_88_144 (.ZN (n_88_144), .A (n_92_144), .B (n_93_146), .C1 (n_94_145), .C2 (n_93_145) );
AOI211_X1 g_86_145 (.ZN (n_86_145), .A (n_90_143), .B (n_94_144), .C1 (n_95_147), .C2 (n_91_144) );
AOI211_X1 g_87_143 (.ZN (n_87_143), .A (n_88_144), .B (n_93_142), .C1 (n_93_146), .C2 (n_93_143) );
AOI211_X1 g_88_145 (.ZN (n_88_145), .A (n_86_145), .B (n_92_144), .C1 (n_94_144), .C2 (n_94_145) );
AOI211_X1 g_87_147 (.ZN (n_87_147), .A (n_87_143), .B (n_90_143), .C1 (n_93_142), .C2 (n_95_147) );
AOI211_X1 g_89_146 (.ZN (n_89_146), .A (n_88_145), .B (n_88_144), .C1 (n_92_144), .C2 (n_93_146) );
AOI211_X1 g_91_145 (.ZN (n_91_145), .A (n_87_147), .B (n_86_145), .C1 (n_90_143), .C2 (n_94_144) );
AOI211_X1 g_92_147 (.ZN (n_92_147), .A (n_89_146), .B (n_87_143), .C1 (n_88_144), .C2 (n_93_142) );
AOI211_X1 g_90_146 (.ZN (n_90_146), .A (n_91_145), .B (n_88_145), .C1 (n_86_145), .C2 (n_92_144) );
AOI211_X1 g_89_144 (.ZN (n_89_144), .A (n_92_147), .B (n_87_147), .C1 (n_87_143), .C2 (n_90_143) );
AOI211_X1 g_88_146 (.ZN (n_88_146), .A (n_90_146), .B (n_89_146), .C1 (n_88_145), .C2 (n_88_144) );
AOI211_X1 g_89_148 (.ZN (n_89_148), .A (n_89_144), .B (n_91_145), .C1 (n_87_147), .C2 (n_86_145) );
AOI211_X1 g_91_147 (.ZN (n_91_147), .A (n_88_146), .B (n_92_147), .C1 (n_89_146), .C2 (n_87_143) );
AOI211_X1 g_90_145 (.ZN (n_90_145), .A (n_89_148), .B (n_90_146), .C1 (n_91_145), .C2 (n_88_145) );
AOI211_X1 g_91_143 (.ZN (n_91_143), .A (n_91_147), .B (n_89_144), .C1 (n_92_147), .C2 (n_87_147) );
AOI211_X1 g_92_145 (.ZN (n_92_145), .A (n_90_145), .B (n_88_146), .C1 (n_90_146), .C2 (n_89_146) );
AOI211_X1 g_94_146 (.ZN (n_94_146), .A (n_91_143), .B (n_89_148), .C1 (n_89_144), .C2 (n_91_145) );
AOI211_X1 g_93_144 (.ZN (n_93_144), .A (n_92_145), .B (n_91_147), .C1 (n_88_146), .C2 (n_92_147) );
AOI211_X1 g_95_143 (.ZN (n_95_143), .A (n_94_146), .B (n_90_145), .C1 (n_89_148), .C2 (n_90_146) );
AOI211_X1 g_96_145 (.ZN (n_96_145), .A (n_93_144), .B (n_91_143), .C1 (n_91_147), .C2 (n_89_144) );
AOI211_X1 g_97_143 (.ZN (n_97_143), .A (n_95_143), .B (n_92_145), .C1 (n_90_145), .C2 (n_88_146) );
AOI211_X1 g_95_144 (.ZN (n_95_144), .A (n_96_145), .B (n_94_146), .C1 (n_91_143), .C2 (n_89_148) );
AOI211_X1 g_96_142 (.ZN (n_96_142), .A (n_97_143), .B (n_93_144), .C1 (n_92_145), .C2 (n_91_147) );
AOI211_X1 g_94_143 (.ZN (n_94_143), .A (n_95_144), .B (n_95_143), .C1 (n_94_146), .C2 (n_90_145) );
AOI211_X1 g_95_141 (.ZN (n_95_141), .A (n_96_142), .B (n_96_145), .C1 (n_93_144), .C2 (n_91_143) );
AOI211_X1 g_97_140 (.ZN (n_97_140), .A (n_94_143), .B (n_97_143), .C1 (n_95_143), .C2 (n_92_145) );
AOI211_X1 g_99_139 (.ZN (n_99_139), .A (n_95_141), .B (n_95_144), .C1 (n_96_145), .C2 (n_94_146) );
AOI211_X1 g_98_141 (.ZN (n_98_141), .A (n_97_140), .B (n_96_142), .C1 (n_97_143), .C2 (n_93_144) );
AOI211_X1 g_100_140 (.ZN (n_100_140), .A (n_99_139), .B (n_94_143), .C1 (n_95_144), .C2 (n_95_143) );
AOI211_X1 g_101_138 (.ZN (n_101_138), .A (n_98_141), .B (n_95_141), .C1 (n_96_142), .C2 (n_96_145) );
AOI211_X1 g_103_137 (.ZN (n_103_137), .A (n_100_140), .B (n_97_140), .C1 (n_94_143), .C2 (n_97_143) );
AOI211_X1 g_102_139 (.ZN (n_102_139), .A (n_101_138), .B (n_99_139), .C1 (n_95_141), .C2 (n_95_144) );
AOI211_X1 g_104_138 (.ZN (n_104_138), .A (n_103_137), .B (n_98_141), .C1 (n_97_140), .C2 (n_96_142) );
AOI211_X1 g_103_140 (.ZN (n_103_140), .A (n_102_139), .B (n_100_140), .C1 (n_99_139), .C2 (n_94_143) );
AOI211_X1 g_105_139 (.ZN (n_105_139), .A (n_104_138), .B (n_101_138), .C1 (n_98_141), .C2 (n_95_141) );
AOI211_X1 g_107_140 (.ZN (n_107_140), .A (n_103_140), .B (n_103_137), .C1 (n_100_140), .C2 (n_97_140) );
AOI211_X1 g_109_139 (.ZN (n_109_139), .A (n_105_139), .B (n_102_139), .C1 (n_101_138), .C2 (n_99_139) );
AOI211_X1 g_110_137 (.ZN (n_110_137), .A (n_107_140), .B (n_104_138), .C1 (n_103_137), .C2 (n_98_141) );
AOI211_X1 g_111_135 (.ZN (n_111_135), .A (n_109_139), .B (n_103_140), .C1 (n_102_139), .C2 (n_100_140) );
AOI211_X1 g_113_134 (.ZN (n_113_134), .A (n_110_137), .B (n_105_139), .C1 (n_104_138), .C2 (n_101_138) );
AOI211_X1 g_115_133 (.ZN (n_115_133), .A (n_111_135), .B (n_107_140), .C1 (n_103_140), .C2 (n_103_137) );
AOI211_X1 g_114_135 (.ZN (n_114_135), .A (n_113_134), .B (n_109_139), .C1 (n_105_139), .C2 (n_102_139) );
AOI211_X1 g_112_136 (.ZN (n_112_136), .A (n_115_133), .B (n_110_137), .C1 (n_107_140), .C2 (n_104_138) );
AOI211_X1 g_111_138 (.ZN (n_111_138), .A (n_114_135), .B (n_111_135), .C1 (n_109_139), .C2 (n_103_140) );
AOI211_X1 g_109_137 (.ZN (n_109_137), .A (n_112_136), .B (n_113_134), .C1 (n_110_137), .C2 (n_105_139) );
AOI211_X1 g_111_136 (.ZN (n_111_136), .A (n_111_138), .B (n_115_133), .C1 (n_111_135), .C2 (n_107_140) );
AOI211_X1 g_113_135 (.ZN (n_113_135), .A (n_109_137), .B (n_114_135), .C1 (n_113_134), .C2 (n_109_139) );
AOI211_X1 g_115_134 (.ZN (n_115_134), .A (n_111_136), .B (n_112_136), .C1 (n_115_133), .C2 (n_110_137) );
AOI211_X1 g_117_133 (.ZN (n_117_133), .A (n_113_135), .B (n_111_138), .C1 (n_114_135), .C2 (n_111_135) );
AOI211_X1 g_119_132 (.ZN (n_119_132), .A (n_115_134), .B (n_109_137), .C1 (n_112_136), .C2 (n_113_134) );
AOI211_X1 g_121_131 (.ZN (n_121_131), .A (n_117_133), .B (n_111_136), .C1 (n_111_138), .C2 (n_115_133) );
AOI211_X1 g_123_130 (.ZN (n_123_130), .A (n_119_132), .B (n_113_135), .C1 (n_109_137), .C2 (n_114_135) );
AOI211_X1 g_122_132 (.ZN (n_122_132), .A (n_121_131), .B (n_115_134), .C1 (n_111_136), .C2 (n_112_136) );
AOI211_X1 g_120_131 (.ZN (n_120_131), .A (n_123_130), .B (n_117_133), .C1 (n_113_135), .C2 (n_111_138) );
AOI211_X1 g_122_130 (.ZN (n_122_130), .A (n_122_132), .B (n_119_132), .C1 (n_115_134), .C2 (n_109_137) );
AOI211_X1 g_124_129 (.ZN (n_124_129), .A (n_120_131), .B (n_121_131), .C1 (n_117_133), .C2 (n_111_136) );
AOI211_X1 g_126_128 (.ZN (n_126_128), .A (n_122_130), .B (n_123_130), .C1 (n_119_132), .C2 (n_113_135) );
AOI211_X1 g_128_127 (.ZN (n_128_127), .A (n_124_129), .B (n_122_132), .C1 (n_121_131), .C2 (n_115_134) );
AOI211_X1 g_130_126 (.ZN (n_130_126), .A (n_126_128), .B (n_120_131), .C1 (n_123_130), .C2 (n_117_133) );
AOI211_X1 g_132_125 (.ZN (n_132_125), .A (n_128_127), .B (n_122_130), .C1 (n_122_132), .C2 (n_119_132) );
AOI211_X1 g_134_124 (.ZN (n_134_124), .A (n_130_126), .B (n_124_129), .C1 (n_120_131), .C2 (n_121_131) );
AOI211_X1 g_136_123 (.ZN (n_136_123), .A (n_132_125), .B (n_126_128), .C1 (n_122_130), .C2 (n_123_130) );
AOI211_X1 g_138_122 (.ZN (n_138_122), .A (n_134_124), .B (n_128_127), .C1 (n_124_129), .C2 (n_122_132) );
AOI211_X1 g_140_121 (.ZN (n_140_121), .A (n_136_123), .B (n_130_126), .C1 (n_126_128), .C2 (n_120_131) );
AOI211_X1 g_142_120 (.ZN (n_142_120), .A (n_138_122), .B (n_132_125), .C1 (n_128_127), .C2 (n_122_130) );
AOI211_X1 g_143_122 (.ZN (n_143_122), .A (n_140_121), .B (n_134_124), .C1 (n_130_126), .C2 (n_124_129) );
AOI211_X1 g_141_123 (.ZN (n_141_123), .A (n_142_120), .B (n_136_123), .C1 (n_132_125), .C2 (n_126_128) );
AOI211_X1 g_142_121 (.ZN (n_142_121), .A (n_143_122), .B (n_138_122), .C1 (n_134_124), .C2 (n_128_127) );
AOI211_X1 g_143_119 (.ZN (n_143_119), .A (n_141_123), .B (n_140_121), .C1 (n_136_123), .C2 (n_130_126) );
AOI211_X1 g_141_120 (.ZN (n_141_120), .A (n_142_121), .B (n_142_120), .C1 (n_138_122), .C2 (n_132_125) );
AOI211_X1 g_140_122 (.ZN (n_140_122), .A (n_143_119), .B (n_143_122), .C1 (n_140_121), .C2 (n_134_124) );
AOI211_X1 g_138_123 (.ZN (n_138_123), .A (n_141_120), .B (n_141_123), .C1 (n_142_120), .C2 (n_136_123) );
AOI211_X1 g_136_124 (.ZN (n_136_124), .A (n_140_122), .B (n_142_121), .C1 (n_143_122), .C2 (n_138_122) );
AOI211_X1 g_134_125 (.ZN (n_134_125), .A (n_138_123), .B (n_143_119), .C1 (n_141_123), .C2 (n_140_121) );
AOI211_X1 g_132_126 (.ZN (n_132_126), .A (n_136_124), .B (n_141_120), .C1 (n_142_121), .C2 (n_142_120) );
AOI211_X1 g_130_127 (.ZN (n_130_127), .A (n_134_125), .B (n_140_122), .C1 (n_143_119), .C2 (n_143_122) );
AOI211_X1 g_128_128 (.ZN (n_128_128), .A (n_132_126), .B (n_138_123), .C1 (n_141_120), .C2 (n_141_123) );
AOI211_X1 g_129_126 (.ZN (n_129_126), .A (n_130_127), .B (n_136_124), .C1 (n_140_122), .C2 (n_142_121) );
AOI211_X1 g_127_127 (.ZN (n_127_127), .A (n_128_128), .B (n_134_125), .C1 (n_138_123), .C2 (n_143_119) );
AOI211_X1 g_126_129 (.ZN (n_126_129), .A (n_129_126), .B (n_132_126), .C1 (n_136_124), .C2 (n_141_120) );
AOI211_X1 g_124_130 (.ZN (n_124_130), .A (n_127_127), .B (n_130_127), .C1 (n_134_125), .C2 (n_140_122) );
AOI211_X1 g_122_131 (.ZN (n_122_131), .A (n_126_129), .B (n_128_128), .C1 (n_132_126), .C2 (n_138_123) );
AOI211_X1 g_120_132 (.ZN (n_120_132), .A (n_124_130), .B (n_129_126), .C1 (n_130_127), .C2 (n_136_124) );
AOI211_X1 g_118_133 (.ZN (n_118_133), .A (n_122_131), .B (n_127_127), .C1 (n_128_128), .C2 (n_134_125) );
AOI211_X1 g_116_134 (.ZN (n_116_134), .A (n_120_132), .B (n_126_129), .C1 (n_129_126), .C2 (n_132_126) );
AOI211_X1 g_115_136 (.ZN (n_115_136), .A (n_118_133), .B (n_124_130), .C1 (n_127_127), .C2 (n_130_127) );
AOI211_X1 g_113_137 (.ZN (n_113_137), .A (n_116_134), .B (n_122_131), .C1 (n_126_129), .C2 (n_128_128) );
AOI211_X1 g_112_139 (.ZN (n_112_139), .A (n_115_136), .B (n_120_132), .C1 (n_124_130), .C2 (n_129_126) );
AOI211_X1 g_111_137 (.ZN (n_111_137), .A (n_113_137), .B (n_118_133), .C1 (n_122_131), .C2 (n_127_127) );
AOI211_X1 g_109_136 (.ZN (n_109_136), .A (n_112_139), .B (n_116_134), .C1 (n_120_132), .C2 (n_126_129) );
AOI211_X1 g_108_138 (.ZN (n_108_138), .A (n_111_137), .B (n_115_136), .C1 (n_118_133), .C2 (n_124_130) );
AOI211_X1 g_106_139 (.ZN (n_106_139), .A (n_109_136), .B (n_113_137), .C1 (n_116_134), .C2 (n_122_131) );
AOI211_X1 g_107_137 (.ZN (n_107_137), .A (n_108_138), .B (n_112_139), .C1 (n_115_136), .C2 (n_120_132) );
AOI211_X1 g_105_138 (.ZN (n_105_138), .A (n_106_139), .B (n_111_137), .C1 (n_113_137), .C2 (n_118_133) );
AOI211_X1 g_103_139 (.ZN (n_103_139), .A (n_107_137), .B (n_109_136), .C1 (n_112_139), .C2 (n_116_134) );
AOI211_X1 g_101_140 (.ZN (n_101_140), .A (n_105_138), .B (n_108_138), .C1 (n_111_137), .C2 (n_115_136) );
AOI211_X1 g_99_141 (.ZN (n_99_141), .A (n_103_139), .B (n_106_139), .C1 (n_109_136), .C2 (n_113_137) );
AOI211_X1 g_97_142 (.ZN (n_97_142), .A (n_101_140), .B (n_107_137), .C1 (n_108_138), .C2 (n_112_139) );
AOI211_X1 g_96_144 (.ZN (n_96_144), .A (n_99_141), .B (n_105_138), .C1 (n_106_139), .C2 (n_111_137) );
AOI211_X1 g_98_145 (.ZN (n_98_145), .A (n_97_142), .B (n_103_139), .C1 (n_107_137), .C2 (n_109_136) );
AOI211_X1 g_99_147 (.ZN (n_99_147), .A (n_96_144), .B (n_101_140), .C1 (n_105_138), .C2 (n_108_138) );
AOI211_X1 g_100_149 (.ZN (n_100_149), .A (n_98_145), .B (n_99_141), .C1 (n_103_139), .C2 (n_106_139) );
AOI211_X1 g_101_147 (.ZN (n_101_147), .A (n_99_147), .B (n_97_142), .C1 (n_101_140), .C2 (n_107_137) );
AOI211_X1 g_102_145 (.ZN (n_102_145), .A (n_100_149), .B (n_96_144), .C1 (n_99_141), .C2 (n_105_138) );
AOI211_X1 g_103_147 (.ZN (n_103_147), .A (n_101_147), .B (n_98_145), .C1 (n_97_142), .C2 (n_103_139) );
AOI211_X1 g_104_149 (.ZN (n_104_149), .A (n_102_145), .B (n_99_147), .C1 (n_96_144), .C2 (n_101_140) );
AOI211_X1 g_105_147 (.ZN (n_105_147), .A (n_103_147), .B (n_100_149), .C1 (n_98_145), .C2 (n_99_141) );
AOI211_X1 g_106_145 (.ZN (n_106_145), .A (n_104_149), .B (n_101_147), .C1 (n_99_147), .C2 (n_97_142) );
AOI211_X1 g_107_147 (.ZN (n_107_147), .A (n_105_147), .B (n_102_145), .C1 (n_100_149), .C2 (n_96_144) );
AOI211_X1 g_108_149 (.ZN (n_108_149), .A (n_106_145), .B (n_103_147), .C1 (n_101_147), .C2 (n_98_145) );
AOI211_X1 g_109_147 (.ZN (n_109_147), .A (n_107_147), .B (n_104_149), .C1 (n_102_145), .C2 (n_99_147) );
AOI211_X1 g_110_145 (.ZN (n_110_145), .A (n_108_149), .B (n_105_147), .C1 (n_103_147), .C2 (n_100_149) );
AOI211_X1 g_111_147 (.ZN (n_111_147), .A (n_109_147), .B (n_106_145), .C1 (n_104_149), .C2 (n_101_147) );
AOI211_X1 g_112_149 (.ZN (n_112_149), .A (n_110_145), .B (n_107_147), .C1 (n_105_147), .C2 (n_102_145) );
AOI211_X1 g_113_147 (.ZN (n_113_147), .A (n_111_147), .B (n_108_149), .C1 (n_106_145), .C2 (n_103_147) );
AOI211_X1 g_114_145 (.ZN (n_114_145), .A (n_112_149), .B (n_109_147), .C1 (n_107_147), .C2 (n_104_149) );
AOI211_X1 g_115_147 (.ZN (n_115_147), .A (n_113_147), .B (n_110_145), .C1 (n_108_149), .C2 (n_105_147) );
AOI211_X1 g_116_149 (.ZN (n_116_149), .A (n_114_145), .B (n_111_147), .C1 (n_109_147), .C2 (n_106_145) );
AOI211_X1 g_117_147 (.ZN (n_117_147), .A (n_115_147), .B (n_112_149), .C1 (n_110_145), .C2 (n_107_147) );
AOI211_X1 g_118_145 (.ZN (n_118_145), .A (n_116_149), .B (n_113_147), .C1 (n_111_147), .C2 (n_108_149) );
AOI211_X1 g_119_147 (.ZN (n_119_147), .A (n_117_147), .B (n_114_145), .C1 (n_112_149), .C2 (n_109_147) );
AOI211_X1 g_120_149 (.ZN (n_120_149), .A (n_118_145), .B (n_115_147), .C1 (n_113_147), .C2 (n_110_145) );
AOI211_X1 g_121_147 (.ZN (n_121_147), .A (n_119_147), .B (n_116_149), .C1 (n_114_145), .C2 (n_111_147) );
AOI211_X1 g_122_145 (.ZN (n_122_145), .A (n_120_149), .B (n_117_147), .C1 (n_115_147), .C2 (n_112_149) );
AOI211_X1 g_123_147 (.ZN (n_123_147), .A (n_121_147), .B (n_118_145), .C1 (n_116_149), .C2 (n_113_147) );
AOI211_X1 g_124_149 (.ZN (n_124_149), .A (n_122_145), .B (n_119_147), .C1 (n_117_147), .C2 (n_114_145) );
AOI211_X1 g_125_147 (.ZN (n_125_147), .A (n_123_147), .B (n_120_149), .C1 (n_118_145), .C2 (n_115_147) );
AOI211_X1 g_126_145 (.ZN (n_126_145), .A (n_124_149), .B (n_121_147), .C1 (n_119_147), .C2 (n_116_149) );
AOI211_X1 g_127_147 (.ZN (n_127_147), .A (n_125_147), .B (n_122_145), .C1 (n_120_149), .C2 (n_117_147) );
AOI211_X1 g_128_149 (.ZN (n_128_149), .A (n_126_145), .B (n_123_147), .C1 (n_121_147), .C2 (n_118_145) );
AOI211_X1 g_130_148 (.ZN (n_130_148), .A (n_127_147), .B (n_124_149), .C1 (n_122_145), .C2 (n_119_147) );
AOI211_X1 g_132_147 (.ZN (n_132_147), .A (n_128_149), .B (n_125_147), .C1 (n_123_147), .C2 (n_120_149) );
AOI211_X1 g_134_146 (.ZN (n_134_146), .A (n_130_148), .B (n_126_145), .C1 (n_124_149), .C2 (n_121_147) );
AOI211_X1 g_136_145 (.ZN (n_136_145), .A (n_132_147), .B (n_127_147), .C1 (n_125_147), .C2 (n_122_145) );
AOI211_X1 g_137_143 (.ZN (n_137_143), .A (n_134_146), .B (n_128_149), .C1 (n_126_145), .C2 (n_123_147) );
AOI211_X1 g_139_142 (.ZN (n_139_142), .A (n_136_145), .B (n_130_148), .C1 (n_127_147), .C2 (n_124_149) );
AOI211_X1 g_141_141 (.ZN (n_141_141), .A (n_137_143), .B (n_132_147), .C1 (n_128_149), .C2 (n_125_147) );
AOI211_X1 g_142_139 (.ZN (n_142_139), .A (n_139_142), .B (n_134_146), .C1 (n_130_148), .C2 (n_126_145) );
AOI211_X1 g_143_141 (.ZN (n_143_141), .A (n_141_141), .B (n_136_145), .C1 (n_132_147), .C2 (n_127_147) );
AOI211_X1 g_141_142 (.ZN (n_141_142), .A (n_142_139), .B (n_137_143), .C1 (n_134_146), .C2 (n_128_149) );
AOI211_X1 g_140_140 (.ZN (n_140_140), .A (n_143_141), .B (n_139_142), .C1 (n_136_145), .C2 (n_130_148) );
AOI211_X1 g_138_141 (.ZN (n_138_141), .A (n_141_142), .B (n_141_141), .C1 (n_137_143), .C2 (n_132_147) );
AOI211_X1 g_136_140 (.ZN (n_136_140), .A (n_140_140), .B (n_142_139), .C1 (n_139_142), .C2 (n_134_146) );
AOI211_X1 g_135_142 (.ZN (n_135_142), .A (n_138_141), .B (n_143_141), .C1 (n_141_141), .C2 (n_136_145) );
AOI211_X1 g_137_141 (.ZN (n_137_141), .A (n_136_140), .B (n_141_142), .C1 (n_142_139), .C2 (n_137_143) );
AOI211_X1 g_139_140 (.ZN (n_139_140), .A (n_135_142), .B (n_140_140), .C1 (n_143_141), .C2 (n_139_142) );
AOI211_X1 g_141_139 (.ZN (n_141_139), .A (n_137_141), .B (n_138_141), .C1 (n_141_142), .C2 (n_141_141) );
AOI211_X1 g_140_141 (.ZN (n_140_141), .A (n_139_140), .B (n_136_140), .C1 (n_140_140), .C2 (n_142_139) );
AOI211_X1 g_142_140 (.ZN (n_142_140), .A (n_141_139), .B (n_135_142), .C1 (n_138_141), .C2 (n_143_141) );
AOI211_X1 g_144_139 (.ZN (n_144_139), .A (n_140_141), .B (n_137_141), .C1 (n_136_140), .C2 (n_141_142) );
AOI211_X1 g_145_137 (.ZN (n_145_137), .A (n_142_140), .B (n_139_140), .C1 (n_135_142), .C2 (n_140_140) );
AOI211_X1 g_143_138 (.ZN (n_143_138), .A (n_144_139), .B (n_141_139), .C1 (n_137_141), .C2 (n_138_141) );
AOI211_X1 g_144_136 (.ZN (n_144_136), .A (n_145_137), .B (n_140_141), .C1 (n_139_140), .C2 (n_136_140) );
AOI211_X1 g_146_135 (.ZN (n_146_135), .A (n_143_138), .B (n_142_140), .C1 (n_141_139), .C2 (n_135_142) );
AOI211_X1 g_147_133 (.ZN (n_147_133), .A (n_144_136), .B (n_144_139), .C1 (n_140_141), .C2 (n_137_141) );
AOI211_X1 g_145_134 (.ZN (n_145_134), .A (n_146_135), .B (n_145_137), .C1 (n_142_140), .C2 (n_139_140) );
AOI211_X1 g_143_135 (.ZN (n_143_135), .A (n_147_133), .B (n_143_138), .C1 (n_144_139), .C2 (n_141_139) );
AOI211_X1 g_142_137 (.ZN (n_142_137), .A (n_145_134), .B (n_144_136), .C1 (n_145_137), .C2 (n_140_141) );
AOI211_X1 g_140_138 (.ZN (n_140_138), .A (n_143_135), .B (n_146_135), .C1 (n_143_138), .C2 (n_142_140) );
AOI211_X1 g_141_140 (.ZN (n_141_140), .A (n_142_137), .B (n_147_133), .C1 (n_144_136), .C2 (n_144_139) );
AOI211_X1 g_139_141 (.ZN (n_139_141), .A (n_140_138), .B (n_145_134), .C1 (n_146_135), .C2 (n_145_137) );
AOI211_X1 g_138_139 (.ZN (n_138_139), .A (n_141_140), .B (n_143_135), .C1 (n_147_133), .C2 (n_143_138) );
AOI211_X1 g_139_137 (.ZN (n_139_137), .A (n_139_141), .B (n_142_137), .C1 (n_145_134), .C2 (n_144_136) );
AOI211_X1 g_140_139 (.ZN (n_140_139), .A (n_138_139), .B (n_140_138), .C1 (n_143_135), .C2 (n_146_135) );
AOI211_X1 g_142_138 (.ZN (n_142_138), .A (n_139_137), .B (n_141_140), .C1 (n_142_137), .C2 (n_147_133) );
AOI211_X1 g_143_136 (.ZN (n_143_136), .A (n_140_139), .B (n_139_141), .C1 (n_140_138), .C2 (n_145_134) );
AOI211_X1 g_144_134 (.ZN (n_144_134), .A (n_142_138), .B (n_138_139), .C1 (n_141_140), .C2 (n_143_135) );
AOI211_X1 g_145_132 (.ZN (n_145_132), .A (n_143_136), .B (n_139_137), .C1 (n_139_141), .C2 (n_142_137) );
AOI211_X1 g_143_131 (.ZN (n_143_131), .A (n_144_134), .B (n_140_139), .C1 (n_138_139), .C2 (n_140_138) );
AOI211_X1 g_145_130 (.ZN (n_145_130), .A (n_145_132), .B (n_142_138), .C1 (n_139_137), .C2 (n_141_140) );
AOI211_X1 g_147_129 (.ZN (n_147_129), .A (n_143_131), .B (n_143_136), .C1 (n_140_139), .C2 (n_139_141) );
AOI211_X1 g_145_128 (.ZN (n_145_128), .A (n_145_130), .B (n_144_134), .C1 (n_142_138), .C2 (n_138_139) );
AOI211_X1 g_143_127 (.ZN (n_143_127), .A (n_147_129), .B (n_145_132), .C1 (n_143_136), .C2 (n_139_137) );
AOI211_X1 g_145_126 (.ZN (n_145_126), .A (n_145_128), .B (n_143_131), .C1 (n_144_134), .C2 (n_140_139) );
AOI211_X1 g_147_125 (.ZN (n_147_125), .A (n_143_127), .B (n_145_130), .C1 (n_145_132), .C2 (n_142_138) );
AOI211_X1 g_146_123 (.ZN (n_146_123), .A (n_145_126), .B (n_147_129), .C1 (n_143_131), .C2 (n_143_136) );
AOI211_X1 g_144_124 (.ZN (n_144_124), .A (n_147_125), .B (n_145_128), .C1 (n_145_130), .C2 (n_144_134) );
AOI211_X1 g_142_123 (.ZN (n_142_123), .A (n_146_123), .B (n_143_127), .C1 (n_147_129), .C2 (n_145_132) );
AOI211_X1 g_144_122 (.ZN (n_144_122), .A (n_144_124), .B (n_145_126), .C1 (n_145_128), .C2 (n_143_131) );
AOI211_X1 g_145_120 (.ZN (n_145_120), .A (n_142_123), .B (n_147_125), .C1 (n_143_127), .C2 (n_145_130) );
AOI211_X1 g_143_121 (.ZN (n_143_121), .A (n_144_122), .B (n_146_123), .C1 (n_145_126), .C2 (n_147_129) );
AOI211_X1 g_141_122 (.ZN (n_141_122), .A (n_145_120), .B (n_144_124), .C1 (n_147_125), .C2 (n_145_128) );
AOI211_X1 g_139_123 (.ZN (n_139_123), .A (n_143_121), .B (n_142_123), .C1 (n_146_123), .C2 (n_143_127) );
AOI211_X1 g_137_124 (.ZN (n_137_124), .A (n_141_122), .B (n_144_122), .C1 (n_144_124), .C2 (n_145_126) );
AOI211_X1 g_135_125 (.ZN (n_135_125), .A (n_139_123), .B (n_145_120), .C1 (n_142_123), .C2 (n_147_125) );
AOI211_X1 g_133_126 (.ZN (n_133_126), .A (n_137_124), .B (n_143_121), .C1 (n_144_122), .C2 (n_146_123) );
AOI211_X1 g_131_127 (.ZN (n_131_127), .A (n_135_125), .B (n_141_122), .C1 (n_145_120), .C2 (n_144_124) );
AOI211_X1 g_129_128 (.ZN (n_129_128), .A (n_133_126), .B (n_139_123), .C1 (n_143_121), .C2 (n_142_123) );
AOI211_X1 g_127_129 (.ZN (n_127_129), .A (n_131_127), .B (n_137_124), .C1 (n_141_122), .C2 (n_144_122) );
AOI211_X1 g_125_130 (.ZN (n_125_130), .A (n_129_128), .B (n_135_125), .C1 (n_139_123), .C2 (n_145_120) );
AOI211_X1 g_123_131 (.ZN (n_123_131), .A (n_127_129), .B (n_133_126), .C1 (n_137_124), .C2 (n_143_121) );
AOI211_X1 g_121_132 (.ZN (n_121_132), .A (n_125_130), .B (n_131_127), .C1 (n_135_125), .C2 (n_141_122) );
AOI211_X1 g_119_133 (.ZN (n_119_133), .A (n_123_131), .B (n_129_128), .C1 (n_133_126), .C2 (n_139_123) );
AOI211_X1 g_117_134 (.ZN (n_117_134), .A (n_121_132), .B (n_127_129), .C1 (n_131_127), .C2 (n_137_124) );
AOI211_X1 g_115_135 (.ZN (n_115_135), .A (n_119_133), .B (n_125_130), .C1 (n_129_128), .C2 (n_135_125) );
AOI211_X1 g_113_136 (.ZN (n_113_136), .A (n_117_134), .B (n_123_131), .C1 (n_127_129), .C2 (n_133_126) );
AOI211_X1 g_112_138 (.ZN (n_112_138), .A (n_115_135), .B (n_121_132), .C1 (n_125_130), .C2 (n_131_127) );
AOI211_X1 g_114_137 (.ZN (n_114_137), .A (n_113_136), .B (n_119_133), .C1 (n_123_131), .C2 (n_129_128) );
AOI211_X1 g_116_136 (.ZN (n_116_136), .A (n_112_138), .B (n_117_134), .C1 (n_121_132), .C2 (n_127_129) );
AOI211_X1 g_118_135 (.ZN (n_118_135), .A (n_114_137), .B (n_115_135), .C1 (n_119_133), .C2 (n_125_130) );
AOI211_X1 g_120_134 (.ZN (n_120_134), .A (n_116_136), .B (n_113_136), .C1 (n_117_134), .C2 (n_123_131) );
AOI211_X1 g_122_133 (.ZN (n_122_133), .A (n_118_135), .B (n_112_138), .C1 (n_115_135), .C2 (n_121_132) );
AOI211_X1 g_124_132 (.ZN (n_124_132), .A (n_120_134), .B (n_114_137), .C1 (n_113_136), .C2 (n_119_133) );
AOI211_X1 g_126_131 (.ZN (n_126_131), .A (n_122_133), .B (n_116_136), .C1 (n_112_138), .C2 (n_117_134) );
AOI211_X1 g_128_130 (.ZN (n_128_130), .A (n_124_132), .B (n_118_135), .C1 (n_114_137), .C2 (n_115_135) );
AOI211_X1 g_130_129 (.ZN (n_130_129), .A (n_126_131), .B (n_120_134), .C1 (n_116_136), .C2 (n_113_136) );
AOI211_X1 g_132_128 (.ZN (n_132_128), .A (n_128_130), .B (n_122_133), .C1 (n_118_135), .C2 (n_112_138) );
AOI211_X1 g_134_127 (.ZN (n_134_127), .A (n_130_129), .B (n_124_132), .C1 (n_120_134), .C2 (n_114_137) );
AOI211_X1 g_136_126 (.ZN (n_136_126), .A (n_132_128), .B (n_126_131), .C1 (n_122_133), .C2 (n_116_136) );
AOI211_X1 g_138_125 (.ZN (n_138_125), .A (n_134_127), .B (n_128_130), .C1 (n_124_132), .C2 (n_118_135) );
AOI211_X1 g_140_124 (.ZN (n_140_124), .A (n_136_126), .B (n_130_129), .C1 (n_126_131), .C2 (n_120_134) );
AOI211_X1 g_142_125 (.ZN (n_142_125), .A (n_138_125), .B (n_132_128), .C1 (n_128_130), .C2 (n_122_133) );
AOI211_X1 g_143_123 (.ZN (n_143_123), .A (n_140_124), .B (n_134_127), .C1 (n_130_129), .C2 (n_124_132) );
AOI211_X1 g_144_121 (.ZN (n_144_121), .A (n_142_125), .B (n_136_126), .C1 (n_132_128), .C2 (n_126_131) );
AOI211_X1 g_146_122 (.ZN (n_146_122), .A (n_143_123), .B (n_138_125), .C1 (n_134_127), .C2 (n_128_130) );
AOI211_X1 g_145_124 (.ZN (n_145_124), .A (n_144_121), .B (n_140_124), .C1 (n_136_126), .C2 (n_130_129) );
AOI211_X1 g_144_126 (.ZN (n_144_126), .A (n_146_122), .B (n_142_125), .C1 (n_138_125), .C2 (n_132_128) );
AOI211_X1 g_146_127 (.ZN (n_146_127), .A (n_145_124), .B (n_143_123), .C1 (n_140_124), .C2 (n_134_127) );
AOI211_X1 g_145_125 (.ZN (n_145_125), .A (n_144_126), .B (n_144_121), .C1 (n_142_125), .C2 (n_136_126) );
AOI211_X1 g_144_123 (.ZN (n_144_123), .A (n_146_127), .B (n_146_122), .C1 (n_143_123), .C2 (n_138_125) );
AOI211_X1 g_142_122 (.ZN (n_142_122), .A (n_145_125), .B (n_145_124), .C1 (n_144_121), .C2 (n_140_124) );
AOI211_X1 g_143_124 (.ZN (n_143_124), .A (n_144_123), .B (n_144_126), .C1 (n_146_122), .C2 (n_142_125) );
AOI211_X1 g_141_125 (.ZN (n_141_125), .A (n_142_122), .B (n_146_127), .C1 (n_145_124), .C2 (n_143_123) );
AOI211_X1 g_140_123 (.ZN (n_140_123), .A (n_143_124), .B (n_145_125), .C1 (n_144_126), .C2 (n_144_121) );
AOI211_X1 g_142_124 (.ZN (n_142_124), .A (n_141_125), .B (n_144_123), .C1 (n_146_127), .C2 (n_146_122) );
AOI211_X1 g_143_126 (.ZN (n_143_126), .A (n_140_123), .B (n_142_122), .C1 (n_145_125), .C2 (n_145_124) );
AOI211_X1 g_144_128 (.ZN (n_144_128), .A (n_142_124), .B (n_143_124), .C1 (n_144_123), .C2 (n_144_126) );
AOI211_X1 g_142_127 (.ZN (n_142_127), .A (n_143_126), .B (n_141_125), .C1 (n_142_122), .C2 (n_146_127) );
AOI211_X1 g_143_125 (.ZN (n_143_125), .A (n_144_128), .B (n_140_123), .C1 (n_143_124), .C2 (n_145_125) );
AOI211_X1 g_141_124 (.ZN (n_141_124), .A (n_142_127), .B (n_142_124), .C1 (n_141_125), .C2 (n_144_123) );
AOI211_X1 g_139_125 (.ZN (n_139_125), .A (n_143_125), .B (n_143_126), .C1 (n_140_123), .C2 (n_142_122) );
AOI211_X1 g_141_126 (.ZN (n_141_126), .A (n_141_124), .B (n_144_128), .C1 (n_142_124), .C2 (n_143_124) );
AOI211_X1 g_142_128 (.ZN (n_142_128), .A (n_139_125), .B (n_142_127), .C1 (n_143_126), .C2 (n_141_125) );
AOI211_X1 g_144_127 (.ZN (n_144_127), .A (n_141_126), .B (n_143_125), .C1 (n_144_128), .C2 (n_140_123) );
AOI211_X1 g_142_126 (.ZN (n_142_126), .A (n_142_128), .B (n_141_124), .C1 (n_142_127), .C2 (n_142_124) );
AOI211_X1 g_140_125 (.ZN (n_140_125), .A (n_144_127), .B (n_139_125), .C1 (n_143_125), .C2 (n_143_126) );
AOI211_X1 g_138_124 (.ZN (n_138_124), .A (n_142_126), .B (n_141_126), .C1 (n_141_124), .C2 (n_144_128) );
AOI211_X1 g_136_125 (.ZN (n_136_125), .A (n_140_125), .B (n_142_128), .C1 (n_139_125), .C2 (n_142_127) );
AOI211_X1 g_134_126 (.ZN (n_134_126), .A (n_138_124), .B (n_144_127), .C1 (n_141_126), .C2 (n_143_125) );
AOI211_X1 g_132_127 (.ZN (n_132_127), .A (n_136_125), .B (n_142_126), .C1 (n_142_128), .C2 (n_141_124) );
AOI211_X1 g_130_128 (.ZN (n_130_128), .A (n_134_126), .B (n_140_125), .C1 (n_144_127), .C2 (n_139_125) );
AOI211_X1 g_128_129 (.ZN (n_128_129), .A (n_132_127), .B (n_138_124), .C1 (n_142_126), .C2 (n_141_126) );
AOI211_X1 g_126_130 (.ZN (n_126_130), .A (n_130_128), .B (n_136_125), .C1 (n_140_125), .C2 (n_142_128) );
AOI211_X1 g_124_131 (.ZN (n_124_131), .A (n_128_129), .B (n_134_126), .C1 (n_138_124), .C2 (n_144_127) );
AOI211_X1 g_123_133 (.ZN (n_123_133), .A (n_126_130), .B (n_132_127), .C1 (n_136_125), .C2 (n_142_126) );
AOI211_X1 g_125_132 (.ZN (n_125_132), .A (n_124_131), .B (n_130_128), .C1 (n_134_126), .C2 (n_140_125) );
AOI211_X1 g_127_131 (.ZN (n_127_131), .A (n_123_133), .B (n_128_129), .C1 (n_132_127), .C2 (n_138_124) );
AOI211_X1 g_129_130 (.ZN (n_129_130), .A (n_125_132), .B (n_126_130), .C1 (n_130_128), .C2 (n_136_125) );
AOI211_X1 g_131_129 (.ZN (n_131_129), .A (n_127_131), .B (n_124_131), .C1 (n_128_129), .C2 (n_134_126) );
AOI211_X1 g_133_128 (.ZN (n_133_128), .A (n_129_130), .B (n_123_133), .C1 (n_126_130), .C2 (n_132_127) );
AOI211_X1 g_135_127 (.ZN (n_135_127), .A (n_131_129), .B (n_125_132), .C1 (n_124_131), .C2 (n_130_128) );
AOI211_X1 g_137_126 (.ZN (n_137_126), .A (n_133_128), .B (n_127_131), .C1 (n_123_133), .C2 (n_128_129) );
AOI211_X1 g_139_127 (.ZN (n_139_127), .A (n_135_127), .B (n_129_130), .C1 (n_125_132), .C2 (n_126_130) );
AOI211_X1 g_137_128 (.ZN (n_137_128), .A (n_137_126), .B (n_131_129), .C1 (n_127_131), .C2 (n_124_131) );
AOI211_X1 g_138_126 (.ZN (n_138_126), .A (n_139_127), .B (n_133_128), .C1 (n_129_130), .C2 (n_123_133) );
AOI211_X1 g_139_124 (.ZN (n_139_124), .A (n_137_128), .B (n_135_127), .C1 (n_131_129), .C2 (n_125_132) );
AOI211_X1 g_140_126 (.ZN (n_140_126), .A (n_138_126), .B (n_137_126), .C1 (n_133_128), .C2 (n_127_131) );
AOI211_X1 g_141_128 (.ZN (n_141_128), .A (n_139_124), .B (n_139_127), .C1 (n_135_127), .C2 (n_129_130) );
AOI211_X1 g_143_129 (.ZN (n_143_129), .A (n_140_126), .B (n_137_128), .C1 (n_137_126), .C2 (n_131_129) );
AOI211_X1 g_141_130 (.ZN (n_141_130), .A (n_141_128), .B (n_138_126), .C1 (n_139_127), .C2 (n_133_128) );
AOI211_X1 g_140_128 (.ZN (n_140_128), .A (n_143_129), .B (n_139_124), .C1 (n_137_128), .C2 (n_135_127) );
AOI211_X1 g_139_126 (.ZN (n_139_126), .A (n_141_130), .B (n_140_126), .C1 (n_138_126), .C2 (n_137_126) );
AOI211_X1 g_137_125 (.ZN (n_137_125), .A (n_140_128), .B (n_141_128), .C1 (n_139_124), .C2 (n_139_127) );
AOI211_X1 g_138_127 (.ZN (n_138_127), .A (n_139_126), .B (n_143_129), .C1 (n_140_126), .C2 (n_137_128) );
AOI211_X1 g_139_129 (.ZN (n_139_129), .A (n_137_125), .B (n_141_130), .C1 (n_141_128), .C2 (n_138_126) );
AOI211_X1 g_140_127 (.ZN (n_140_127), .A (n_138_127), .B (n_140_128), .C1 (n_143_129), .C2 (n_139_124) );
AOI211_X1 g_138_128 (.ZN (n_138_128), .A (n_139_129), .B (n_139_126), .C1 (n_141_130), .C2 (n_140_126) );
AOI211_X1 g_136_127 (.ZN (n_136_127), .A (n_140_127), .B (n_137_125), .C1 (n_140_128), .C2 (n_141_128) );
AOI211_X1 g_135_129 (.ZN (n_135_129), .A (n_138_128), .B (n_138_127), .C1 (n_139_126), .C2 (n_143_129) );
AOI211_X1 g_133_130 (.ZN (n_133_130), .A (n_136_127), .B (n_139_129), .C1 (n_137_125), .C2 (n_141_130) );
AOI211_X1 g_134_128 (.ZN (n_134_128), .A (n_135_129), .B (n_140_127), .C1 (n_138_127), .C2 (n_140_128) );
AOI211_X1 g_135_126 (.ZN (n_135_126), .A (n_133_130), .B (n_138_128), .C1 (n_139_129), .C2 (n_139_126) );
AOI211_X1 g_133_127 (.ZN (n_133_127), .A (n_134_128), .B (n_136_127), .C1 (n_140_127), .C2 (n_137_125) );
AOI211_X1 g_131_128 (.ZN (n_131_128), .A (n_135_126), .B (n_135_129), .C1 (n_138_128), .C2 (n_138_127) );
AOI211_X1 g_129_129 (.ZN (n_129_129), .A (n_133_127), .B (n_133_130), .C1 (n_136_127), .C2 (n_139_129) );
AOI211_X1 g_127_130 (.ZN (n_127_130), .A (n_131_128), .B (n_134_128), .C1 (n_135_129), .C2 (n_140_127) );
AOI211_X1 g_125_131 (.ZN (n_125_131), .A (n_129_129), .B (n_135_126), .C1 (n_133_130), .C2 (n_138_128) );
AOI211_X1 g_123_132 (.ZN (n_123_132), .A (n_127_130), .B (n_133_127), .C1 (n_134_128), .C2 (n_136_127) );
AOI211_X1 g_121_133 (.ZN (n_121_133), .A (n_125_131), .B (n_131_128), .C1 (n_135_126), .C2 (n_135_129) );
AOI211_X1 g_119_134 (.ZN (n_119_134), .A (n_123_132), .B (n_129_129), .C1 (n_133_127), .C2 (n_133_130) );
AOI211_X1 g_117_135 (.ZN (n_117_135), .A (n_121_133), .B (n_127_130), .C1 (n_131_128), .C2 (n_134_128) );
AOI211_X1 g_116_137 (.ZN (n_116_137), .A (n_119_134), .B (n_125_131), .C1 (n_129_129), .C2 (n_135_126) );
AOI211_X1 g_114_136 (.ZN (n_114_136), .A (n_117_135), .B (n_123_132), .C1 (n_127_130), .C2 (n_133_127) );
AOI211_X1 g_116_135 (.ZN (n_116_135), .A (n_116_137), .B (n_121_133), .C1 (n_125_131), .C2 (n_131_128) );
AOI211_X1 g_118_134 (.ZN (n_118_134), .A (n_114_136), .B (n_119_134), .C1 (n_123_132), .C2 (n_129_129) );
AOI211_X1 g_120_133 (.ZN (n_120_133), .A (n_116_135), .B (n_117_135), .C1 (n_121_133), .C2 (n_127_130) );
AOI211_X1 g_119_135 (.ZN (n_119_135), .A (n_118_134), .B (n_116_137), .C1 (n_119_134), .C2 (n_125_131) );
AOI211_X1 g_121_134 (.ZN (n_121_134), .A (n_120_133), .B (n_114_136), .C1 (n_117_135), .C2 (n_123_132) );
AOI211_X1 g_120_136 (.ZN (n_120_136), .A (n_119_135), .B (n_116_135), .C1 (n_116_137), .C2 (n_121_133) );
AOI211_X1 g_122_135 (.ZN (n_122_135), .A (n_121_134), .B (n_118_134), .C1 (n_114_136), .C2 (n_119_134) );
AOI211_X1 g_124_134 (.ZN (n_124_134), .A (n_120_136), .B (n_120_133), .C1 (n_116_135), .C2 (n_117_135) );
AOI211_X1 g_126_133 (.ZN (n_126_133), .A (n_122_135), .B (n_119_135), .C1 (n_118_134), .C2 (n_116_137) );
AOI211_X1 g_128_132 (.ZN (n_128_132), .A (n_124_134), .B (n_121_134), .C1 (n_120_133), .C2 (n_114_136) );
AOI211_X1 g_130_131 (.ZN (n_130_131), .A (n_126_133), .B (n_120_136), .C1 (n_119_135), .C2 (n_116_135) );
AOI211_X1 g_132_130 (.ZN (n_132_130), .A (n_128_132), .B (n_122_135), .C1 (n_121_134), .C2 (n_118_134) );
AOI211_X1 g_134_129 (.ZN (n_134_129), .A (n_130_131), .B (n_124_134), .C1 (n_120_136), .C2 (n_120_133) );
AOI211_X1 g_136_128 (.ZN (n_136_128), .A (n_132_130), .B (n_126_133), .C1 (n_122_135), .C2 (n_119_135) );
AOI211_X1 g_137_130 (.ZN (n_137_130), .A (n_134_129), .B (n_128_132), .C1 (n_124_134), .C2 (n_121_134) );
AOI211_X1 g_135_131 (.ZN (n_135_131), .A (n_136_128), .B (n_130_131), .C1 (n_126_133), .C2 (n_120_136) );
AOI211_X1 g_136_129 (.ZN (n_136_129), .A (n_137_130), .B (n_132_130), .C1 (n_128_132), .C2 (n_122_135) );
AOI211_X1 g_137_127 (.ZN (n_137_127), .A (n_135_131), .B (n_134_129), .C1 (n_130_131), .C2 (n_124_134) );
AOI211_X1 g_135_128 (.ZN (n_135_128), .A (n_136_129), .B (n_136_128), .C1 (n_132_130), .C2 (n_126_133) );
AOI211_X1 g_133_129 (.ZN (n_133_129), .A (n_137_127), .B (n_137_130), .C1 (n_134_129), .C2 (n_128_132) );
AOI211_X1 g_131_130 (.ZN (n_131_130), .A (n_135_128), .B (n_135_131), .C1 (n_136_128), .C2 (n_130_131) );
AOI211_X1 g_129_131 (.ZN (n_129_131), .A (n_133_129), .B (n_136_129), .C1 (n_137_130), .C2 (n_132_130) );
AOI211_X1 g_127_132 (.ZN (n_127_132), .A (n_131_130), .B (n_137_127), .C1 (n_135_131), .C2 (n_134_129) );
AOI211_X1 g_125_133 (.ZN (n_125_133), .A (n_129_131), .B (n_135_128), .C1 (n_136_129), .C2 (n_136_128) );
AOI211_X1 g_123_134 (.ZN (n_123_134), .A (n_127_132), .B (n_133_129), .C1 (n_137_127), .C2 (n_137_130) );
AOI211_X1 g_121_135 (.ZN (n_121_135), .A (n_125_133), .B (n_131_130), .C1 (n_135_128), .C2 (n_135_131) );
AOI211_X1 g_119_136 (.ZN (n_119_136), .A (n_123_134), .B (n_129_131), .C1 (n_133_129), .C2 (n_136_129) );
AOI211_X1 g_117_137 (.ZN (n_117_137), .A (n_121_135), .B (n_127_132), .C1 (n_131_130), .C2 (n_137_127) );
AOI211_X1 g_115_138 (.ZN (n_115_138), .A (n_119_136), .B (n_125_133), .C1 (n_129_131), .C2 (n_135_128) );
AOI211_X1 g_113_139 (.ZN (n_113_139), .A (n_117_137), .B (n_123_134), .C1 (n_127_132), .C2 (n_133_129) );
AOI211_X1 g_112_137 (.ZN (n_112_137), .A (n_115_138), .B (n_121_135), .C1 (n_125_133), .C2 (n_131_130) );
AOI211_X1 g_110_138 (.ZN (n_110_138), .A (n_113_139), .B (n_119_136), .C1 (n_123_134), .C2 (n_129_131) );
AOI211_X1 g_108_139 (.ZN (n_108_139), .A (n_112_137), .B (n_117_137), .C1 (n_121_135), .C2 (n_127_132) );
AOI211_X1 g_106_140 (.ZN (n_106_140), .A (n_110_138), .B (n_115_138), .C1 (n_119_136), .C2 (n_125_133) );
AOI211_X1 g_104_139 (.ZN (n_104_139), .A (n_108_139), .B (n_113_139), .C1 (n_117_137), .C2 (n_123_134) );
AOI211_X1 g_102_140 (.ZN (n_102_140), .A (n_106_140), .B (n_112_137), .C1 (n_115_138), .C2 (n_121_135) );
AOI211_X1 g_100_141 (.ZN (n_100_141), .A (n_104_139), .B (n_110_138), .C1 (n_113_139), .C2 (n_119_136) );
AOI211_X1 g_98_142 (.ZN (n_98_142), .A (n_102_140), .B (n_108_139), .C1 (n_112_137), .C2 (n_117_137) );
AOI211_X1 g_96_143 (.ZN (n_96_143), .A (n_100_141), .B (n_106_140), .C1 (n_110_138), .C2 (n_115_138) );
AOI211_X1 g_95_145 (.ZN (n_95_145), .A (n_98_142), .B (n_104_139), .C1 (n_108_139), .C2 (n_113_139) );
AOI211_X1 g_97_144 (.ZN (n_97_144), .A (n_96_143), .B (n_102_140), .C1 (n_106_140), .C2 (n_112_137) );
AOI211_X1 g_99_143 (.ZN (n_99_143), .A (n_95_145), .B (n_100_141), .C1 (n_104_139), .C2 (n_110_138) );
AOI211_X1 g_101_142 (.ZN (n_101_142), .A (n_97_144), .B (n_98_142), .C1 (n_102_140), .C2 (n_108_139) );
AOI211_X1 g_103_141 (.ZN (n_103_141), .A (n_99_143), .B (n_96_143), .C1 (n_100_141), .C2 (n_106_140) );
AOI211_X1 g_105_140 (.ZN (n_105_140), .A (n_101_142), .B (n_95_145), .C1 (n_98_142), .C2 (n_104_139) );
AOI211_X1 g_107_139 (.ZN (n_107_139), .A (n_103_141), .B (n_97_144), .C1 (n_96_143), .C2 (n_102_140) );
AOI211_X1 g_109_138 (.ZN (n_109_138), .A (n_105_140), .B (n_99_143), .C1 (n_95_145), .C2 (n_100_141) );
AOI211_X1 g_110_140 (.ZN (n_110_140), .A (n_107_139), .B (n_101_142), .C1 (n_97_144), .C2 (n_98_142) );
AOI211_X1 g_108_141 (.ZN (n_108_141), .A (n_109_138), .B (n_103_141), .C1 (n_99_143), .C2 (n_96_143) );
AOI211_X1 g_106_142 (.ZN (n_106_142), .A (n_110_140), .B (n_105_140), .C1 (n_101_142), .C2 (n_95_145) );
AOI211_X1 g_104_141 (.ZN (n_104_141), .A (n_108_141), .B (n_107_139), .C1 (n_103_141), .C2 (n_97_144) );
AOI211_X1 g_102_142 (.ZN (n_102_142), .A (n_106_142), .B (n_109_138), .C1 (n_105_140), .C2 (n_99_143) );
AOI211_X1 g_100_143 (.ZN (n_100_143), .A (n_104_141), .B (n_110_140), .C1 (n_107_139), .C2 (n_101_142) );
AOI211_X1 g_101_141 (.ZN (n_101_141), .A (n_102_142), .B (n_108_141), .C1 (n_109_138), .C2 (n_103_141) );
AOI211_X1 g_99_142 (.ZN (n_99_142), .A (n_100_143), .B (n_106_142), .C1 (n_110_140), .C2 (n_105_140) );
AOI211_X1 g_98_144 (.ZN (n_98_144), .A (n_101_141), .B (n_104_141), .C1 (n_108_141), .C2 (n_107_139) );
AOI211_X1 g_97_146 (.ZN (n_97_146), .A (n_99_142), .B (n_102_142), .C1 (n_106_142), .C2 (n_109_138) );
AOI211_X1 g_98_148 (.ZN (n_98_148), .A (n_98_144), .B (n_100_143), .C1 (n_104_141), .C2 (n_110_140) );
AOI211_X1 g_96_147 (.ZN (n_96_147), .A (n_97_146), .B (n_101_141), .C1 (n_102_142), .C2 (n_108_141) );
AOI211_X1 g_98_146 (.ZN (n_98_146), .A (n_98_148), .B (n_99_142), .C1 (n_100_143), .C2 (n_106_142) );
AOI211_X1 g_100_145 (.ZN (n_100_145), .A (n_96_147), .B (n_98_144), .C1 (n_101_141), .C2 (n_104_141) );
AOI211_X1 g_101_143 (.ZN (n_101_143), .A (n_98_146), .B (n_97_146), .C1 (n_99_142), .C2 (n_102_142) );
AOI211_X1 g_99_144 (.ZN (n_99_144), .A (n_100_145), .B (n_98_148), .C1 (n_98_144), .C2 (n_100_143) );
AOI211_X1 g_97_145 (.ZN (n_97_145), .A (n_101_143), .B (n_96_147), .C1 (n_97_146), .C2 (n_101_141) );
AOI211_X1 g_99_146 (.ZN (n_99_146), .A (n_99_144), .B (n_98_146), .C1 (n_98_148), .C2 (n_99_142) );
AOI211_X1 g_100_144 (.ZN (n_100_144), .A (n_97_145), .B (n_100_145), .C1 (n_96_147), .C2 (n_98_144) );
AOI211_X1 g_98_143 (.ZN (n_98_143), .A (n_99_146), .B (n_101_143), .C1 (n_98_146), .C2 (n_97_146) );
AOI211_X1 g_100_142 (.ZN (n_100_142), .A (n_100_144), .B (n_99_144), .C1 (n_100_145), .C2 (n_98_148) );
AOI211_X1 g_102_141 (.ZN (n_102_141), .A (n_98_143), .B (n_97_145), .C1 (n_101_143), .C2 (n_96_147) );
AOI211_X1 g_104_140 (.ZN (n_104_140), .A (n_100_142), .B (n_99_146), .C1 (n_99_144), .C2 (n_98_146) );
AOI211_X1 g_103_142 (.ZN (n_103_142), .A (n_102_141), .B (n_100_144), .C1 (n_97_145), .C2 (n_100_145) );
AOI211_X1 g_105_141 (.ZN (n_105_141), .A (n_104_140), .B (n_98_143), .C1 (n_99_146), .C2 (n_101_143) );
AOI211_X1 g_104_143 (.ZN (n_104_143), .A (n_103_142), .B (n_100_142), .C1 (n_100_144), .C2 (n_99_144) );
AOI211_X1 g_102_144 (.ZN (n_102_144), .A (n_105_141), .B (n_102_141), .C1 (n_98_143), .C2 (n_97_145) );
AOI211_X1 g_101_146 (.ZN (n_101_146), .A (n_104_143), .B (n_104_140), .C1 (n_100_142), .C2 (n_99_146) );
AOI211_X1 g_99_145 (.ZN (n_99_145), .A (n_102_144), .B (n_103_142), .C1 (n_102_141), .C2 (n_100_144) );
AOI211_X1 g_101_144 (.ZN (n_101_144), .A (n_101_146), .B (n_105_141), .C1 (n_104_140), .C2 (n_98_143) );
AOI211_X1 g_103_143 (.ZN (n_103_143), .A (n_99_145), .B (n_104_143), .C1 (n_103_142), .C2 (n_100_142) );
AOI211_X1 g_105_142 (.ZN (n_105_142), .A (n_101_144), .B (n_102_144), .C1 (n_105_141), .C2 (n_102_141) );
AOI211_X1 g_107_141 (.ZN (n_107_141), .A (n_103_143), .B (n_101_146), .C1 (n_104_143), .C2 (n_104_140) );
AOI211_X1 g_109_140 (.ZN (n_109_140), .A (n_105_142), .B (n_99_145), .C1 (n_102_144), .C2 (n_103_142) );
AOI211_X1 g_111_139 (.ZN (n_111_139), .A (n_107_141), .B (n_101_144), .C1 (n_101_146), .C2 (n_105_141) );
AOI211_X1 g_113_138 (.ZN (n_113_138), .A (n_109_140), .B (n_103_143), .C1 (n_99_145), .C2 (n_104_143) );
AOI211_X1 g_115_137 (.ZN (n_115_137), .A (n_111_139), .B (n_105_142), .C1 (n_101_144), .C2 (n_102_144) );
AOI211_X1 g_117_136 (.ZN (n_117_136), .A (n_113_138), .B (n_107_141), .C1 (n_103_143), .C2 (n_101_146) );
AOI211_X1 g_116_138 (.ZN (n_116_138), .A (n_115_137), .B (n_109_140), .C1 (n_105_142), .C2 (n_99_145) );
AOI211_X1 g_118_137 (.ZN (n_118_137), .A (n_117_136), .B (n_111_139), .C1 (n_107_141), .C2 (n_101_144) );
AOI211_X1 g_117_139 (.ZN (n_117_139), .A (n_116_138), .B (n_113_138), .C1 (n_109_140), .C2 (n_103_143) );
AOI211_X1 g_119_138 (.ZN (n_119_138), .A (n_118_137), .B (n_115_137), .C1 (n_111_139), .C2 (n_105_142) );
AOI211_X1 g_118_136 (.ZN (n_118_136), .A (n_117_139), .B (n_117_136), .C1 (n_113_138), .C2 (n_107_141) );
AOI211_X1 g_120_135 (.ZN (n_120_135), .A (n_119_138), .B (n_116_138), .C1 (n_115_137), .C2 (n_109_140) );
AOI211_X1 g_122_134 (.ZN (n_122_134), .A (n_118_136), .B (n_118_137), .C1 (n_117_136), .C2 (n_111_139) );
AOI211_X1 g_124_133 (.ZN (n_124_133), .A (n_120_135), .B (n_117_139), .C1 (n_116_138), .C2 (n_113_138) );
AOI211_X1 g_126_132 (.ZN (n_126_132), .A (n_122_134), .B (n_119_138), .C1 (n_118_137), .C2 (n_115_137) );
AOI211_X1 g_128_131 (.ZN (n_128_131), .A (n_124_133), .B (n_118_136), .C1 (n_117_139), .C2 (n_117_136) );
AOI211_X1 g_130_130 (.ZN (n_130_130), .A (n_126_132), .B (n_120_135), .C1 (n_119_138), .C2 (n_116_138) );
AOI211_X1 g_132_129 (.ZN (n_132_129), .A (n_128_131), .B (n_122_134), .C1 (n_118_136), .C2 (n_118_137) );
AOI211_X1 g_131_131 (.ZN (n_131_131), .A (n_130_130), .B (n_124_133), .C1 (n_120_135), .C2 (n_117_139) );
AOI211_X1 g_129_132 (.ZN (n_129_132), .A (n_132_129), .B (n_126_132), .C1 (n_122_134), .C2 (n_119_138) );
AOI211_X1 g_127_133 (.ZN (n_127_133), .A (n_131_131), .B (n_128_131), .C1 (n_124_133), .C2 (n_118_136) );
AOI211_X1 g_125_134 (.ZN (n_125_134), .A (n_129_132), .B (n_130_130), .C1 (n_126_132), .C2 (n_120_135) );
AOI211_X1 g_123_135 (.ZN (n_123_135), .A (n_127_133), .B (n_132_129), .C1 (n_128_131), .C2 (n_122_134) );
AOI211_X1 g_121_136 (.ZN (n_121_136), .A (n_125_134), .B (n_131_131), .C1 (n_130_130), .C2 (n_124_133) );
AOI211_X1 g_119_137 (.ZN (n_119_137), .A (n_123_135), .B (n_129_132), .C1 (n_132_129), .C2 (n_126_132) );
AOI211_X1 g_117_138 (.ZN (n_117_138), .A (n_121_136), .B (n_127_133), .C1 (n_131_131), .C2 (n_128_131) );
AOI211_X1 g_115_139 (.ZN (n_115_139), .A (n_119_137), .B (n_125_134), .C1 (n_129_132), .C2 (n_130_130) );
AOI211_X1 g_113_140 (.ZN (n_113_140), .A (n_117_138), .B (n_123_135), .C1 (n_127_133), .C2 (n_132_129) );
AOI211_X1 g_114_138 (.ZN (n_114_138), .A (n_115_139), .B (n_121_136), .C1 (n_125_134), .C2 (n_131_131) );
AOI211_X1 g_115_140 (.ZN (n_115_140), .A (n_113_140), .B (n_119_137), .C1 (n_123_135), .C2 (n_129_132) );
AOI211_X1 g_113_141 (.ZN (n_113_141), .A (n_114_138), .B (n_117_138), .C1 (n_121_136), .C2 (n_127_133) );
AOI211_X1 g_114_139 (.ZN (n_114_139), .A (n_115_140), .B (n_115_139), .C1 (n_119_137), .C2 (n_125_134) );
AOI211_X1 g_112_140 (.ZN (n_112_140), .A (n_113_141), .B (n_113_140), .C1 (n_117_138), .C2 (n_123_135) );
AOI211_X1 g_110_139 (.ZN (n_110_139), .A (n_114_139), .B (n_114_138), .C1 (n_115_139), .C2 (n_121_136) );
AOI211_X1 g_108_140 (.ZN (n_108_140), .A (n_112_140), .B (n_115_140), .C1 (n_113_140), .C2 (n_119_137) );
AOI211_X1 g_106_141 (.ZN (n_106_141), .A (n_110_139), .B (n_113_141), .C1 (n_114_138), .C2 (n_117_138) );
AOI211_X1 g_104_142 (.ZN (n_104_142), .A (n_108_140), .B (n_114_139), .C1 (n_115_140), .C2 (n_115_139) );
AOI211_X1 g_102_143 (.ZN (n_102_143), .A (n_106_141), .B (n_112_140), .C1 (n_113_141), .C2 (n_113_140) );
AOI211_X1 g_101_145 (.ZN (n_101_145), .A (n_104_142), .B (n_110_139), .C1 (n_114_139), .C2 (n_114_138) );
AOI211_X1 g_100_147 (.ZN (n_100_147), .A (n_102_143), .B (n_108_140), .C1 (n_112_140), .C2 (n_115_140) );
AOI211_X1 g_102_148 (.ZN (n_102_148), .A (n_101_145), .B (n_106_141), .C1 (n_110_139), .C2 (n_113_141) );
AOI211_X1 g_103_146 (.ZN (n_103_146), .A (n_100_147), .B (n_104_142), .C1 (n_108_140), .C2 (n_114_139) );
AOI211_X1 g_104_144 (.ZN (n_104_144), .A (n_102_148), .B (n_102_143), .C1 (n_106_141), .C2 (n_112_140) );
AOI211_X1 g_106_143 (.ZN (n_106_143), .A (n_103_146), .B (n_101_145), .C1 (n_104_142), .C2 (n_110_139) );
AOI211_X1 g_108_142 (.ZN (n_108_142), .A (n_104_144), .B (n_100_147), .C1 (n_102_143), .C2 (n_108_140) );
AOI211_X1 g_110_141 (.ZN (n_110_141), .A (n_106_143), .B (n_102_148), .C1 (n_101_145), .C2 (n_106_141) );
AOI211_X1 g_109_143 (.ZN (n_109_143), .A (n_108_142), .B (n_103_146), .C1 (n_100_147), .C2 (n_104_142) );
AOI211_X1 g_111_142 (.ZN (n_111_142), .A (n_110_141), .B (n_104_144), .C1 (n_102_148), .C2 (n_102_143) );
AOI211_X1 g_109_141 (.ZN (n_109_141), .A (n_109_143), .B (n_106_143), .C1 (n_103_146), .C2 (n_101_145) );
AOI211_X1 g_111_140 (.ZN (n_111_140), .A (n_111_142), .B (n_108_142), .C1 (n_104_144), .C2 (n_100_147) );
AOI211_X1 g_110_142 (.ZN (n_110_142), .A (n_109_141), .B (n_110_141), .C1 (n_106_143), .C2 (n_102_148) );
AOI211_X1 g_112_141 (.ZN (n_112_141), .A (n_111_140), .B (n_109_143), .C1 (n_108_142), .C2 (n_103_146) );
AOI211_X1 g_114_140 (.ZN (n_114_140), .A (n_110_142), .B (n_111_142), .C1 (n_110_141), .C2 (n_104_144) );
AOI211_X1 g_116_139 (.ZN (n_116_139), .A (n_112_141), .B (n_109_141), .C1 (n_109_143), .C2 (n_106_143) );
AOI211_X1 g_118_138 (.ZN (n_118_138), .A (n_114_140), .B (n_111_140), .C1 (n_111_142), .C2 (n_108_142) );
AOI211_X1 g_120_137 (.ZN (n_120_137), .A (n_116_139), .B (n_110_142), .C1 (n_109_141), .C2 (n_110_141) );
AOI211_X1 g_122_136 (.ZN (n_122_136), .A (n_118_138), .B (n_112_141), .C1 (n_111_140), .C2 (n_109_143) );
AOI211_X1 g_124_135 (.ZN (n_124_135), .A (n_120_137), .B (n_114_140), .C1 (n_110_142), .C2 (n_111_142) );
AOI211_X1 g_126_134 (.ZN (n_126_134), .A (n_122_136), .B (n_116_139), .C1 (n_112_141), .C2 (n_109_141) );
AOI211_X1 g_128_133 (.ZN (n_128_133), .A (n_124_135), .B (n_118_138), .C1 (n_114_140), .C2 (n_111_140) );
AOI211_X1 g_130_132 (.ZN (n_130_132), .A (n_126_134), .B (n_120_137), .C1 (n_116_139), .C2 (n_110_142) );
AOI211_X1 g_132_131 (.ZN (n_132_131), .A (n_128_133), .B (n_122_136), .C1 (n_118_138), .C2 (n_112_141) );
AOI211_X1 g_134_130 (.ZN (n_134_130), .A (n_130_132), .B (n_124_135), .C1 (n_120_137), .C2 (n_114_140) );
AOI211_X1 g_133_132 (.ZN (n_133_132), .A (n_132_131), .B (n_126_134), .C1 (n_122_136), .C2 (n_116_139) );
AOI211_X1 g_131_133 (.ZN (n_131_133), .A (n_134_130), .B (n_128_133), .C1 (n_124_135), .C2 (n_118_138) );
AOI211_X1 g_129_134 (.ZN (n_129_134), .A (n_133_132), .B (n_130_132), .C1 (n_126_134), .C2 (n_120_137) );
AOI211_X1 g_127_135 (.ZN (n_127_135), .A (n_131_133), .B (n_132_131), .C1 (n_128_133), .C2 (n_122_136) );
AOI211_X1 g_125_136 (.ZN (n_125_136), .A (n_129_134), .B (n_134_130), .C1 (n_130_132), .C2 (n_124_135) );
AOI211_X1 g_123_137 (.ZN (n_123_137), .A (n_127_135), .B (n_133_132), .C1 (n_132_131), .C2 (n_126_134) );
AOI211_X1 g_121_138 (.ZN (n_121_138), .A (n_125_136), .B (n_131_133), .C1 (n_134_130), .C2 (n_128_133) );
AOI211_X1 g_119_139 (.ZN (n_119_139), .A (n_123_137), .B (n_129_134), .C1 (n_133_132), .C2 (n_130_132) );
AOI211_X1 g_117_140 (.ZN (n_117_140), .A (n_121_138), .B (n_127_135), .C1 (n_131_133), .C2 (n_132_131) );
AOI211_X1 g_115_141 (.ZN (n_115_141), .A (n_119_139), .B (n_125_136), .C1 (n_129_134), .C2 (n_134_130) );
AOI211_X1 g_113_142 (.ZN (n_113_142), .A (n_117_140), .B (n_123_137), .C1 (n_127_135), .C2 (n_133_132) );
AOI211_X1 g_111_141 (.ZN (n_111_141), .A (n_115_141), .B (n_121_138), .C1 (n_125_136), .C2 (n_131_133) );
AOI211_X1 g_109_142 (.ZN (n_109_142), .A (n_113_142), .B (n_119_139), .C1 (n_123_137), .C2 (n_129_134) );
AOI211_X1 g_107_143 (.ZN (n_107_143), .A (n_111_141), .B (n_117_140), .C1 (n_121_138), .C2 (n_127_135) );
AOI211_X1 g_105_144 (.ZN (n_105_144), .A (n_109_142), .B (n_115_141), .C1 (n_119_139), .C2 (n_125_136) );
AOI211_X1 g_103_145 (.ZN (n_103_145), .A (n_107_143), .B (n_113_142), .C1 (n_117_140), .C2 (n_123_137) );
AOI211_X1 g_105_146 (.ZN (n_105_146), .A (n_105_144), .B (n_111_141), .C1 (n_115_141), .C2 (n_121_138) );
AOI211_X1 g_106_148 (.ZN (n_106_148), .A (n_103_145), .B (n_109_142), .C1 (n_113_142), .C2 (n_119_139) );
AOI211_X1 g_104_147 (.ZN (n_104_147), .A (n_105_146), .B (n_107_143), .C1 (n_111_141), .C2 (n_117_140) );
AOI211_X1 g_102_146 (.ZN (n_102_146), .A (n_106_148), .B (n_105_144), .C1 (n_109_142), .C2 (n_115_141) );
AOI211_X1 g_103_144 (.ZN (n_103_144), .A (n_104_147), .B (n_103_145), .C1 (n_107_143), .C2 (n_113_142) );
AOI211_X1 g_105_145 (.ZN (n_105_145), .A (n_102_146), .B (n_105_146), .C1 (n_105_144), .C2 (n_111_141) );
AOI211_X1 g_107_144 (.ZN (n_107_144), .A (n_103_144), .B (n_106_148), .C1 (n_103_145), .C2 (n_109_142) );
AOI211_X1 g_105_143 (.ZN (n_105_143), .A (n_105_145), .B (n_104_147), .C1 (n_105_146), .C2 (n_107_143) );
AOI211_X1 g_107_142 (.ZN (n_107_142), .A (n_107_144), .B (n_102_146), .C1 (n_106_148), .C2 (n_105_144) );
AOI211_X1 g_108_144 (.ZN (n_108_144), .A (n_105_143), .B (n_103_144), .C1 (n_104_147), .C2 (n_103_145) );
AOI211_X1 g_107_146 (.ZN (n_107_146), .A (n_107_142), .B (n_105_145), .C1 (n_102_146), .C2 (n_105_146) );
AOI211_X1 g_106_144 (.ZN (n_106_144), .A (n_108_144), .B (n_107_144), .C1 (n_103_144), .C2 (n_106_148) );
AOI211_X1 g_104_145 (.ZN (n_104_145), .A (n_107_146), .B (n_105_143), .C1 (n_105_145), .C2 (n_104_147) );
AOI211_X1 g_106_146 (.ZN (n_106_146), .A (n_106_144), .B (n_107_142), .C1 (n_107_144), .C2 (n_102_146) );
AOI211_X1 g_108_145 (.ZN (n_108_145), .A (n_104_145), .B (n_108_144), .C1 (n_105_143), .C2 (n_103_144) );
AOI211_X1 g_110_144 (.ZN (n_110_144), .A (n_106_146), .B (n_107_146), .C1 (n_107_142), .C2 (n_105_145) );
AOI211_X1 g_108_143 (.ZN (n_108_143), .A (n_108_145), .B (n_106_144), .C1 (n_108_144), .C2 (n_107_144) );
AOI211_X1 g_107_145 (.ZN (n_107_145), .A (n_110_144), .B (n_104_145), .C1 (n_107_146), .C2 (n_105_143) );
AOI211_X1 g_109_146 (.ZN (n_109_146), .A (n_108_143), .B (n_106_146), .C1 (n_106_144), .C2 (n_107_142) );
AOI211_X1 g_110_148 (.ZN (n_110_148), .A (n_107_145), .B (n_108_145), .C1 (n_104_145), .C2 (n_108_144) );
AOI211_X1 g_108_147 (.ZN (n_108_147), .A (n_109_146), .B (n_110_144), .C1 (n_106_146), .C2 (n_107_146) );
AOI211_X1 g_109_145 (.ZN (n_109_145), .A (n_110_148), .B (n_108_143), .C1 (n_108_145), .C2 (n_106_144) );
AOI211_X1 g_111_146 (.ZN (n_111_146), .A (n_108_147), .B (n_107_145), .C1 (n_110_144), .C2 (n_104_145) );
AOI211_X1 g_112_144 (.ZN (n_112_144), .A (n_109_145), .B (n_109_146), .C1 (n_108_143), .C2 (n_106_146) );
AOI211_X1 g_110_143 (.ZN (n_110_143), .A (n_111_146), .B (n_110_148), .C1 (n_107_145), .C2 (n_108_145) );
AOI211_X1 g_112_142 (.ZN (n_112_142), .A (n_112_144), .B (n_108_147), .C1 (n_109_146), .C2 (n_110_144) );
AOI211_X1 g_111_144 (.ZN (n_111_144), .A (n_110_143), .B (n_109_145), .C1 (n_110_148), .C2 (n_108_143) );
AOI211_X1 g_110_146 (.ZN (n_110_146), .A (n_112_142), .B (n_111_146), .C1 (n_108_147), .C2 (n_107_145) );
AOI211_X1 g_109_144 (.ZN (n_109_144), .A (n_111_144), .B (n_112_144), .C1 (n_109_145), .C2 (n_109_146) );
AOI211_X1 g_111_143 (.ZN (n_111_143), .A (n_110_146), .B (n_110_143), .C1 (n_111_146), .C2 (n_110_148) );
AOI211_X1 g_112_145 (.ZN (n_112_145), .A (n_109_144), .B (n_112_142), .C1 (n_112_144), .C2 (n_108_147) );
AOI211_X1 g_113_143 (.ZN (n_113_143), .A (n_111_143), .B (n_111_144), .C1 (n_110_143), .C2 (n_109_145) );
AOI211_X1 g_114_141 (.ZN (n_114_141), .A (n_112_145), .B (n_110_146), .C1 (n_112_142), .C2 (n_111_146) );
AOI211_X1 g_116_140 (.ZN (n_116_140), .A (n_113_143), .B (n_109_144), .C1 (n_111_144), .C2 (n_112_144) );
AOI211_X1 g_118_139 (.ZN (n_118_139), .A (n_114_141), .B (n_111_143), .C1 (n_110_146), .C2 (n_110_143) );
AOI211_X1 g_120_138 (.ZN (n_120_138), .A (n_116_140), .B (n_112_145), .C1 (n_109_144), .C2 (n_112_142) );
AOI211_X1 g_122_137 (.ZN (n_122_137), .A (n_118_139), .B (n_113_143), .C1 (n_111_143), .C2 (n_111_144) );
AOI211_X1 g_124_136 (.ZN (n_124_136), .A (n_120_138), .B (n_114_141), .C1 (n_112_145), .C2 (n_110_146) );
AOI211_X1 g_126_135 (.ZN (n_126_135), .A (n_122_137), .B (n_116_140), .C1 (n_113_143), .C2 (n_109_144) );
AOI211_X1 g_128_134 (.ZN (n_128_134), .A (n_124_136), .B (n_118_139), .C1 (n_114_141), .C2 (n_111_143) );
AOI211_X1 g_130_133 (.ZN (n_130_133), .A (n_126_135), .B (n_120_138), .C1 (n_116_140), .C2 (n_112_145) );
AOI211_X1 g_132_132 (.ZN (n_132_132), .A (n_128_134), .B (n_122_137), .C1 (n_118_139), .C2 (n_113_143) );
AOI211_X1 g_134_131 (.ZN (n_134_131), .A (n_130_133), .B (n_124_136), .C1 (n_120_138), .C2 (n_114_141) );
AOI211_X1 g_136_130 (.ZN (n_136_130), .A (n_132_132), .B (n_126_135), .C1 (n_122_137), .C2 (n_116_140) );
AOI211_X1 g_138_129 (.ZN (n_138_129), .A (n_134_131), .B (n_128_134), .C1 (n_124_136), .C2 (n_118_139) );
AOI211_X1 g_139_131 (.ZN (n_139_131), .A (n_136_130), .B (n_130_133), .C1 (n_126_135), .C2 (n_120_138) );
AOI211_X1 g_140_129 (.ZN (n_140_129), .A (n_138_129), .B (n_132_132), .C1 (n_128_134), .C2 (n_122_137) );
AOI211_X1 g_141_127 (.ZN (n_141_127), .A (n_139_131), .B (n_134_131), .C1 (n_130_133), .C2 (n_124_136) );
AOI211_X1 g_142_129 (.ZN (n_142_129), .A (n_140_129), .B (n_136_130), .C1 (n_132_132), .C2 (n_126_135) );
AOI211_X1 g_144_130 (.ZN (n_144_130), .A (n_141_127), .B (n_138_129), .C1 (n_134_131), .C2 (n_128_134) );
AOI211_X1 g_143_128 (.ZN (n_143_128), .A (n_142_129), .B (n_139_131), .C1 (n_136_130), .C2 (n_130_133) );
AOI211_X1 g_145_129 (.ZN (n_145_129), .A (n_144_130), .B (n_140_129), .C1 (n_138_129), .C2 (n_132_132) );
AOI211_X1 g_146_131 (.ZN (n_146_131), .A (n_143_128), .B (n_141_127), .C1 (n_139_131), .C2 (n_134_131) );
AOI211_X1 g_144_132 (.ZN (n_144_132), .A (n_145_129), .B (n_142_129), .C1 (n_140_129), .C2 (n_136_130) );
AOI211_X1 g_143_130 (.ZN (n_143_130), .A (n_146_131), .B (n_144_130), .C1 (n_141_127), .C2 (n_138_129) );
AOI211_X1 g_141_129 (.ZN (n_141_129), .A (n_144_132), .B (n_143_128), .C1 (n_142_129), .C2 (n_139_131) );
AOI211_X1 g_139_128 (.ZN (n_139_128), .A (n_143_130), .B (n_145_129), .C1 (n_144_130), .C2 (n_140_129) );
AOI211_X1 g_137_129 (.ZN (n_137_129), .A (n_141_129), .B (n_146_131), .C1 (n_143_128), .C2 (n_141_127) );
AOI211_X1 g_135_130 (.ZN (n_135_130), .A (n_139_128), .B (n_144_132), .C1 (n_145_129), .C2 (n_142_129) );
AOI211_X1 g_133_131 (.ZN (n_133_131), .A (n_137_129), .B (n_143_130), .C1 (n_146_131), .C2 (n_144_130) );
AOI211_X1 g_131_132 (.ZN (n_131_132), .A (n_135_130), .B (n_141_129), .C1 (n_144_132), .C2 (n_143_128) );
AOI211_X1 g_129_133 (.ZN (n_129_133), .A (n_133_131), .B (n_139_128), .C1 (n_143_130), .C2 (n_145_129) );
AOI211_X1 g_127_134 (.ZN (n_127_134), .A (n_131_132), .B (n_137_129), .C1 (n_141_129), .C2 (n_146_131) );
AOI211_X1 g_125_135 (.ZN (n_125_135), .A (n_129_133), .B (n_135_130), .C1 (n_139_128), .C2 (n_144_132) );
AOI211_X1 g_123_136 (.ZN (n_123_136), .A (n_127_134), .B (n_133_131), .C1 (n_137_129), .C2 (n_143_130) );
AOI211_X1 g_121_137 (.ZN (n_121_137), .A (n_125_135), .B (n_131_132), .C1 (n_135_130), .C2 (n_141_129) );
AOI211_X1 g_120_139 (.ZN (n_120_139), .A (n_123_136), .B (n_129_133), .C1 (n_133_131), .C2 (n_139_128) );
AOI211_X1 g_122_138 (.ZN (n_122_138), .A (n_121_137), .B (n_127_134), .C1 (n_131_132), .C2 (n_137_129) );
AOI211_X1 g_124_137 (.ZN (n_124_137), .A (n_120_139), .B (n_125_135), .C1 (n_129_133), .C2 (n_135_130) );
AOI211_X1 g_126_136 (.ZN (n_126_136), .A (n_122_138), .B (n_123_136), .C1 (n_127_134), .C2 (n_133_131) );
AOI211_X1 g_128_135 (.ZN (n_128_135), .A (n_124_137), .B (n_121_137), .C1 (n_125_135), .C2 (n_131_132) );
AOI211_X1 g_130_134 (.ZN (n_130_134), .A (n_126_136), .B (n_120_139), .C1 (n_123_136), .C2 (n_129_133) );
AOI211_X1 g_132_133 (.ZN (n_132_133), .A (n_128_135), .B (n_122_138), .C1 (n_121_137), .C2 (n_127_134) );
AOI211_X1 g_134_132 (.ZN (n_134_132), .A (n_130_134), .B (n_124_137), .C1 (n_120_139), .C2 (n_125_135) );
AOI211_X1 g_136_131 (.ZN (n_136_131), .A (n_132_133), .B (n_126_136), .C1 (n_122_138), .C2 (n_123_136) );
AOI211_X1 g_138_130 (.ZN (n_138_130), .A (n_134_132), .B (n_128_135), .C1 (n_124_137), .C2 (n_121_137) );
AOI211_X1 g_137_132 (.ZN (n_137_132), .A (n_136_131), .B (n_130_134), .C1 (n_126_136), .C2 (n_120_139) );
AOI211_X1 g_135_133 (.ZN (n_135_133), .A (n_138_130), .B (n_132_133), .C1 (n_128_135), .C2 (n_122_138) );
AOI211_X1 g_133_134 (.ZN (n_133_134), .A (n_137_132), .B (n_134_132), .C1 (n_130_134), .C2 (n_124_137) );
AOI211_X1 g_131_135 (.ZN (n_131_135), .A (n_135_133), .B (n_136_131), .C1 (n_132_133), .C2 (n_126_136) );
AOI211_X1 g_129_136 (.ZN (n_129_136), .A (n_133_134), .B (n_138_130), .C1 (n_134_132), .C2 (n_128_135) );
AOI211_X1 g_127_137 (.ZN (n_127_137), .A (n_131_135), .B (n_137_132), .C1 (n_136_131), .C2 (n_130_134) );
AOI211_X1 g_125_138 (.ZN (n_125_138), .A (n_129_136), .B (n_135_133), .C1 (n_138_130), .C2 (n_132_133) );
AOI211_X1 g_123_139 (.ZN (n_123_139), .A (n_127_137), .B (n_133_134), .C1 (n_137_132), .C2 (n_134_132) );
AOI211_X1 g_121_140 (.ZN (n_121_140), .A (n_125_138), .B (n_131_135), .C1 (n_135_133), .C2 (n_136_131) );
AOI211_X1 g_119_141 (.ZN (n_119_141), .A (n_123_139), .B (n_129_136), .C1 (n_133_134), .C2 (n_138_130) );
AOI211_X1 g_117_142 (.ZN (n_117_142), .A (n_121_140), .B (n_127_137), .C1 (n_131_135), .C2 (n_137_132) );
AOI211_X1 g_118_140 (.ZN (n_118_140), .A (n_119_141), .B (n_125_138), .C1 (n_129_136), .C2 (n_135_133) );
AOI211_X1 g_116_141 (.ZN (n_116_141), .A (n_117_142), .B (n_123_139), .C1 (n_127_137), .C2 (n_133_134) );
AOI211_X1 g_115_143 (.ZN (n_115_143), .A (n_118_140), .B (n_121_140), .C1 (n_125_138), .C2 (n_131_135) );
AOI211_X1 g_113_144 (.ZN (n_113_144), .A (n_116_141), .B (n_119_141), .C1 (n_123_139), .C2 (n_129_136) );
AOI211_X1 g_114_142 (.ZN (n_114_142), .A (n_115_143), .B (n_117_142), .C1 (n_121_140), .C2 (n_127_137) );
AOI211_X1 g_112_143 (.ZN (n_112_143), .A (n_113_144), .B (n_118_140), .C1 (n_119_141), .C2 (n_125_138) );
AOI211_X1 g_111_145 (.ZN (n_111_145), .A (n_114_142), .B (n_116_141), .C1 (n_117_142), .C2 (n_123_139) );
AOI211_X1 g_112_147 (.ZN (n_112_147), .A (n_112_143), .B (n_115_143), .C1 (n_118_140), .C2 (n_121_140) );
AOI211_X1 g_114_146 (.ZN (n_114_146), .A (n_111_145), .B (n_113_144), .C1 (n_116_141), .C2 (n_119_141) );
AOI211_X1 g_116_145 (.ZN (n_116_145), .A (n_112_147), .B (n_114_142), .C1 (n_115_143), .C2 (n_117_142) );
AOI211_X1 g_114_144 (.ZN (n_114_144), .A (n_114_146), .B (n_112_143), .C1 (n_113_144), .C2 (n_118_140) );
AOI211_X1 g_113_146 (.ZN (n_113_146), .A (n_116_145), .B (n_111_145), .C1 (n_114_142), .C2 (n_116_141) );
AOI211_X1 g_114_148 (.ZN (n_114_148), .A (n_114_144), .B (n_112_147), .C1 (n_112_143), .C2 (n_115_143) );
AOI211_X1 g_115_146 (.ZN (n_115_146), .A (n_113_146), .B (n_114_146), .C1 (n_111_145), .C2 (n_113_144) );
AOI211_X1 g_113_145 (.ZN (n_113_145), .A (n_114_148), .B (n_116_145), .C1 (n_112_147), .C2 (n_114_142) );
AOI211_X1 g_115_144 (.ZN (n_115_144), .A (n_115_146), .B (n_114_144), .C1 (n_114_146), .C2 (n_112_143) );
AOI211_X1 g_117_143 (.ZN (n_117_143), .A (n_113_145), .B (n_113_146), .C1 (n_116_145), .C2 (n_111_145) );
AOI211_X1 g_115_142 (.ZN (n_115_142), .A (n_115_144), .B (n_114_148), .C1 (n_114_144), .C2 (n_112_147) );
AOI211_X1 g_116_144 (.ZN (n_116_144), .A (n_117_143), .B (n_115_146), .C1 (n_113_146), .C2 (n_114_146) );
AOI211_X1 g_114_143 (.ZN (n_114_143), .A (n_115_142), .B (n_113_145), .C1 (n_114_148), .C2 (n_116_145) );
AOI211_X1 g_116_142 (.ZN (n_116_142), .A (n_116_144), .B (n_115_144), .C1 (n_115_146), .C2 (n_114_144) );
AOI211_X1 g_118_141 (.ZN (n_118_141), .A (n_114_143), .B (n_117_143), .C1 (n_113_145), .C2 (n_113_146) );
AOI211_X1 g_120_140 (.ZN (n_120_140), .A (n_116_142), .B (n_115_142), .C1 (n_115_144), .C2 (n_114_148) );
AOI211_X1 g_122_139 (.ZN (n_122_139), .A (n_118_141), .B (n_116_144), .C1 (n_117_143), .C2 (n_115_146) );
AOI211_X1 g_124_138 (.ZN (n_124_138), .A (n_120_140), .B (n_114_143), .C1 (n_115_142), .C2 (n_113_145) );
AOI211_X1 g_126_137 (.ZN (n_126_137), .A (n_122_139), .B (n_116_142), .C1 (n_116_144), .C2 (n_115_144) );
AOI211_X1 g_128_136 (.ZN (n_128_136), .A (n_124_138), .B (n_118_141), .C1 (n_114_143), .C2 (n_117_143) );
AOI211_X1 g_130_135 (.ZN (n_130_135), .A (n_126_137), .B (n_120_140), .C1 (n_116_142), .C2 (n_115_142) );
AOI211_X1 g_132_134 (.ZN (n_132_134), .A (n_128_136), .B (n_122_139), .C1 (n_118_141), .C2 (n_116_144) );
AOI211_X1 g_134_133 (.ZN (n_134_133), .A (n_130_135), .B (n_124_138), .C1 (n_120_140), .C2 (n_114_143) );
AOI211_X1 g_136_132 (.ZN (n_136_132), .A (n_132_134), .B (n_126_137), .C1 (n_122_139), .C2 (n_116_142) );
AOI211_X1 g_138_131 (.ZN (n_138_131), .A (n_134_133), .B (n_128_136), .C1 (n_124_138), .C2 (n_118_141) );
AOI211_X1 g_140_130 (.ZN (n_140_130), .A (n_136_132), .B (n_130_135), .C1 (n_126_137), .C2 (n_120_140) );
AOI211_X1 g_142_131 (.ZN (n_142_131), .A (n_138_131), .B (n_132_134), .C1 (n_128_136), .C2 (n_122_139) );
AOI211_X1 g_140_132 (.ZN (n_140_132), .A (n_140_130), .B (n_134_133), .C1 (n_130_135), .C2 (n_124_138) );
AOI211_X1 g_139_130 (.ZN (n_139_130), .A (n_142_131), .B (n_136_132), .C1 (n_132_134), .C2 (n_126_137) );
AOI211_X1 g_137_131 (.ZN (n_137_131), .A (n_140_132), .B (n_138_131), .C1 (n_134_133), .C2 (n_128_136) );
AOI211_X1 g_135_132 (.ZN (n_135_132), .A (n_139_130), .B (n_140_130), .C1 (n_136_132), .C2 (n_130_135) );
AOI211_X1 g_133_133 (.ZN (n_133_133), .A (n_137_131), .B (n_142_131), .C1 (n_138_131), .C2 (n_132_134) );
AOI211_X1 g_131_134 (.ZN (n_131_134), .A (n_135_132), .B (n_140_132), .C1 (n_140_130), .C2 (n_134_133) );
AOI211_X1 g_129_135 (.ZN (n_129_135), .A (n_133_133), .B (n_139_130), .C1 (n_142_131), .C2 (n_136_132) );
AOI211_X1 g_127_136 (.ZN (n_127_136), .A (n_131_134), .B (n_137_131), .C1 (n_140_132), .C2 (n_138_131) );
AOI211_X1 g_125_137 (.ZN (n_125_137), .A (n_129_135), .B (n_135_132), .C1 (n_139_130), .C2 (n_140_130) );
AOI211_X1 g_123_138 (.ZN (n_123_138), .A (n_127_136), .B (n_133_133), .C1 (n_137_131), .C2 (n_142_131) );
AOI211_X1 g_121_139 (.ZN (n_121_139), .A (n_125_137), .B (n_131_134), .C1 (n_135_132), .C2 (n_140_132) );
AOI211_X1 g_119_140 (.ZN (n_119_140), .A (n_123_138), .B (n_129_135), .C1 (n_133_133), .C2 (n_139_130) );
AOI211_X1 g_117_141 (.ZN (n_117_141), .A (n_121_139), .B (n_127_136), .C1 (n_131_134), .C2 (n_137_131) );
AOI211_X1 g_116_143 (.ZN (n_116_143), .A (n_119_140), .B (n_125_137), .C1 (n_129_135), .C2 (n_135_132) );
AOI211_X1 g_115_145 (.ZN (n_115_145), .A (n_117_141), .B (n_123_138), .C1 (n_127_136), .C2 (n_133_133) );
AOI211_X1 g_116_147 (.ZN (n_116_147), .A (n_116_143), .B (n_121_139), .C1 (n_125_137), .C2 (n_131_134) );
AOI211_X1 g_117_145 (.ZN (n_117_145), .A (n_115_145), .B (n_119_140), .C1 (n_123_138), .C2 (n_129_135) );
AOI211_X1 g_118_143 (.ZN (n_118_143), .A (n_116_147), .B (n_117_141), .C1 (n_121_139), .C2 (n_127_136) );
AOI211_X1 g_120_142 (.ZN (n_120_142), .A (n_117_145), .B (n_116_143), .C1 (n_119_140), .C2 (n_125_137) );
AOI211_X1 g_122_141 (.ZN (n_122_141), .A (n_118_143), .B (n_115_145), .C1 (n_117_141), .C2 (n_123_138) );
AOI211_X1 g_124_140 (.ZN (n_124_140), .A (n_120_142), .B (n_116_147), .C1 (n_116_143), .C2 (n_121_139) );
AOI211_X1 g_126_139 (.ZN (n_126_139), .A (n_122_141), .B (n_117_145), .C1 (n_115_145), .C2 (n_119_140) );
AOI211_X1 g_128_138 (.ZN (n_128_138), .A (n_124_140), .B (n_118_143), .C1 (n_116_147), .C2 (n_117_141) );
AOI211_X1 g_130_137 (.ZN (n_130_137), .A (n_126_139), .B (n_120_142), .C1 (n_117_145), .C2 (n_116_143) );
AOI211_X1 g_132_136 (.ZN (n_132_136), .A (n_128_138), .B (n_122_141), .C1 (n_118_143), .C2 (n_115_145) );
AOI211_X1 g_134_135 (.ZN (n_134_135), .A (n_130_137), .B (n_124_140), .C1 (n_120_142), .C2 (n_116_147) );
AOI211_X1 g_136_134 (.ZN (n_136_134), .A (n_132_136), .B (n_126_139), .C1 (n_122_141), .C2 (n_117_145) );
AOI211_X1 g_138_133 (.ZN (n_138_133), .A (n_134_135), .B (n_128_138), .C1 (n_124_140), .C2 (n_118_143) );
AOI211_X1 g_137_135 (.ZN (n_137_135), .A (n_136_134), .B (n_130_137), .C1 (n_126_139), .C2 (n_120_142) );
AOI211_X1 g_136_133 (.ZN (n_136_133), .A (n_138_133), .B (n_132_136), .C1 (n_128_138), .C2 (n_122_141) );
AOI211_X1 g_138_132 (.ZN (n_138_132), .A (n_137_135), .B (n_134_135), .C1 (n_130_137), .C2 (n_124_140) );
AOI211_X1 g_140_131 (.ZN (n_140_131), .A (n_136_133), .B (n_136_134), .C1 (n_132_136), .C2 (n_126_139) );
AOI211_X1 g_142_130 (.ZN (n_142_130), .A (n_138_132), .B (n_138_133), .C1 (n_134_135), .C2 (n_128_138) );
AOI211_X1 g_144_131 (.ZN (n_144_131), .A (n_140_131), .B (n_137_135), .C1 (n_136_134), .C2 (n_130_137) );
AOI211_X1 g_142_132 (.ZN (n_142_132), .A (n_142_130), .B (n_136_133), .C1 (n_138_133), .C2 (n_132_136) );
AOI211_X1 g_143_134 (.ZN (n_143_134), .A (n_144_131), .B (n_138_132), .C1 (n_137_135), .C2 (n_134_135) );
AOI211_X1 g_145_133 (.ZN (n_145_133), .A (n_142_132), .B (n_140_131), .C1 (n_136_133), .C2 (n_136_134) );
AOI211_X1 g_143_132 (.ZN (n_143_132), .A (n_143_134), .B (n_142_130), .C1 (n_138_132), .C2 (n_138_133) );
AOI211_X1 g_141_131 (.ZN (n_141_131), .A (n_145_133), .B (n_144_131), .C1 (n_140_131), .C2 (n_137_135) );
AOI211_X1 g_142_133 (.ZN (n_142_133), .A (n_143_132), .B (n_142_132), .C1 (n_142_130), .C2 (n_136_133) );
AOI211_X1 g_141_135 (.ZN (n_141_135), .A (n_141_131), .B (n_143_134), .C1 (n_144_131), .C2 (n_138_132) );
AOI211_X1 g_140_133 (.ZN (n_140_133), .A (n_142_133), .B (n_145_133), .C1 (n_142_132), .C2 (n_140_131) );
AOI211_X1 g_142_134 (.ZN (n_142_134), .A (n_141_135), .B (n_143_132), .C1 (n_143_134), .C2 (n_142_130) );
AOI211_X1 g_141_132 (.ZN (n_141_132), .A (n_140_133), .B (n_141_131), .C1 (n_145_133), .C2 (n_144_131) );
AOI211_X1 g_143_133 (.ZN (n_143_133), .A (n_142_134), .B (n_142_133), .C1 (n_143_132), .C2 (n_142_132) );
AOI211_X1 g_144_135 (.ZN (n_144_135), .A (n_141_132), .B (n_141_135), .C1 (n_141_131), .C2 (n_143_134) );
AOI211_X1 g_143_137 (.ZN (n_143_137), .A (n_143_133), .B (n_140_133), .C1 (n_142_133), .C2 (n_145_133) );
AOI211_X1 g_141_136 (.ZN (n_141_136), .A (n_144_135), .B (n_142_134), .C1 (n_141_135), .C2 (n_143_132) );
AOI211_X1 g_140_134 (.ZN (n_140_134), .A (n_143_137), .B (n_141_132), .C1 (n_140_133), .C2 (n_141_131) );
AOI211_X1 g_139_132 (.ZN (n_139_132), .A (n_141_136), .B (n_143_133), .C1 (n_142_134), .C2 (n_142_133) );
AOI211_X1 g_141_133 (.ZN (n_141_133), .A (n_140_134), .B (n_144_135), .C1 (n_141_132), .C2 (n_141_135) );
AOI211_X1 g_142_135 (.ZN (n_142_135), .A (n_139_132), .B (n_143_137), .C1 (n_143_133), .C2 (n_140_133) );
AOI211_X1 g_141_137 (.ZN (n_141_137), .A (n_141_133), .B (n_141_136), .C1 (n_144_135), .C2 (n_142_134) );
AOI211_X1 g_139_136 (.ZN (n_139_136), .A (n_142_135), .B (n_140_134), .C1 (n_143_137), .C2 (n_141_132) );
AOI211_X1 g_138_134 (.ZN (n_138_134), .A (n_141_137), .B (n_139_132), .C1 (n_141_136), .C2 (n_143_133) );
AOI211_X1 g_140_135 (.ZN (n_140_135), .A (n_139_136), .B (n_141_133), .C1 (n_140_134), .C2 (n_144_135) );
AOI211_X1 g_139_133 (.ZN (n_139_133), .A (n_138_134), .B (n_142_135), .C1 (n_139_132), .C2 (n_143_137) );
AOI211_X1 g_141_134 (.ZN (n_141_134), .A (n_140_135), .B (n_141_137), .C1 (n_141_133), .C2 (n_141_136) );
AOI211_X1 g_142_136 (.ZN (n_142_136), .A (n_139_133), .B (n_139_136), .C1 (n_142_135), .C2 (n_140_134) );
AOI211_X1 g_141_138 (.ZN (n_141_138), .A (n_141_134), .B (n_138_134), .C1 (n_141_137), .C2 (n_139_132) );
AOI211_X1 g_140_136 (.ZN (n_140_136), .A (n_142_136), .B (n_140_135), .C1 (n_139_136), .C2 (n_141_133) );
AOI211_X1 g_139_134 (.ZN (n_139_134), .A (n_141_138), .B (n_139_133), .C1 (n_138_134), .C2 (n_142_135) );
AOI211_X1 g_137_133 (.ZN (n_137_133), .A (n_140_136), .B (n_141_134), .C1 (n_140_135), .C2 (n_141_137) );
AOI211_X1 g_138_135 (.ZN (n_138_135), .A (n_139_134), .B (n_142_136), .C1 (n_139_133), .C2 (n_139_136) );
AOI211_X1 g_137_137 (.ZN (n_137_137), .A (n_137_133), .B (n_141_138), .C1 (n_141_134), .C2 (n_138_134) );
AOI211_X1 g_139_138 (.ZN (n_139_138), .A (n_138_135), .B (n_140_136), .C1 (n_142_136), .C2 (n_140_135) );
AOI211_X1 g_138_140 (.ZN (n_138_140), .A (n_137_137), .B (n_139_134), .C1 (n_141_138), .C2 (n_139_133) );
AOI211_X1 g_137_138 (.ZN (n_137_138), .A (n_139_138), .B (n_137_133), .C1 (n_140_136), .C2 (n_141_134) );
AOI211_X1 g_139_139 (.ZN (n_139_139), .A (n_138_140), .B (n_138_135), .C1 (n_139_134), .C2 (n_142_136) );
AOI211_X1 g_140_137 (.ZN (n_140_137), .A (n_137_138), .B (n_137_137), .C1 (n_137_133), .C2 (n_141_138) );
AOI211_X1 g_139_135 (.ZN (n_139_135), .A (n_139_139), .B (n_139_138), .C1 (n_138_135), .C2 (n_140_136) );
AOI211_X1 g_137_134 (.ZN (n_137_134), .A (n_140_137), .B (n_138_140), .C1 (n_137_137), .C2 (n_139_134) );
AOI211_X1 g_138_136 (.ZN (n_138_136), .A (n_139_135), .B (n_137_138), .C1 (n_139_138), .C2 (n_137_133) );
AOI211_X1 g_136_135 (.ZN (n_136_135), .A (n_137_134), .B (n_139_139), .C1 (n_138_140), .C2 (n_138_135) );
AOI211_X1 g_134_134 (.ZN (n_134_134), .A (n_138_136), .B (n_140_137), .C1 (n_137_138), .C2 (n_137_137) );
AOI211_X1 g_132_135 (.ZN (n_132_135), .A (n_136_135), .B (n_139_135), .C1 (n_139_139), .C2 (n_139_138) );
AOI211_X1 g_130_136 (.ZN (n_130_136), .A (n_134_134), .B (n_137_134), .C1 (n_140_137), .C2 (n_138_140) );
AOI211_X1 g_128_137 (.ZN (n_128_137), .A (n_132_135), .B (n_138_136), .C1 (n_139_135), .C2 (n_137_138) );
AOI211_X1 g_126_138 (.ZN (n_126_138), .A (n_130_136), .B (n_136_135), .C1 (n_137_134), .C2 (n_139_139) );
AOI211_X1 g_124_139 (.ZN (n_124_139), .A (n_128_137), .B (n_134_134), .C1 (n_138_136), .C2 (n_140_137) );
AOI211_X1 g_122_140 (.ZN (n_122_140), .A (n_126_138), .B (n_132_135), .C1 (n_136_135), .C2 (n_139_135) );
AOI211_X1 g_120_141 (.ZN (n_120_141), .A (n_124_139), .B (n_130_136), .C1 (n_134_134), .C2 (n_137_134) );
AOI211_X1 g_118_142 (.ZN (n_118_142), .A (n_122_140), .B (n_128_137), .C1 (n_132_135), .C2 (n_138_136) );
AOI211_X1 g_117_144 (.ZN (n_117_144), .A (n_120_141), .B (n_126_138), .C1 (n_130_136), .C2 (n_136_135) );
AOI211_X1 g_119_143 (.ZN (n_119_143), .A (n_118_142), .B (n_124_139), .C1 (n_128_137), .C2 (n_134_134) );
AOI211_X1 g_121_142 (.ZN (n_121_142), .A (n_117_144), .B (n_122_140), .C1 (n_126_138), .C2 (n_132_135) );
AOI211_X1 g_123_141 (.ZN (n_123_141), .A (n_119_143), .B (n_120_141), .C1 (n_124_139), .C2 (n_130_136) );
AOI211_X1 g_125_140 (.ZN (n_125_140), .A (n_121_142), .B (n_118_142), .C1 (n_122_140), .C2 (n_128_137) );
AOI211_X1 g_127_139 (.ZN (n_127_139), .A (n_123_141), .B (n_117_144), .C1 (n_120_141), .C2 (n_126_138) );
AOI211_X1 g_129_138 (.ZN (n_129_138), .A (n_125_140), .B (n_119_143), .C1 (n_118_142), .C2 (n_124_139) );
AOI211_X1 g_131_137 (.ZN (n_131_137), .A (n_127_139), .B (n_121_142), .C1 (n_117_144), .C2 (n_122_140) );
AOI211_X1 g_133_136 (.ZN (n_133_136), .A (n_129_138), .B (n_123_141), .C1 (n_119_143), .C2 (n_120_141) );
AOI211_X1 g_135_135 (.ZN (n_135_135), .A (n_131_137), .B (n_125_140), .C1 (n_121_142), .C2 (n_118_142) );
AOI211_X1 g_137_136 (.ZN (n_137_136), .A (n_133_136), .B (n_127_139), .C1 (n_123_141), .C2 (n_117_144) );
AOI211_X1 g_135_137 (.ZN (n_135_137), .A (n_135_135), .B (n_129_138), .C1 (n_125_140), .C2 (n_119_143) );
AOI211_X1 g_136_139 (.ZN (n_136_139), .A (n_137_136), .B (n_131_137), .C1 (n_127_139), .C2 (n_121_142) );
AOI211_X1 g_138_138 (.ZN (n_138_138), .A (n_135_137), .B (n_133_136), .C1 (n_129_138), .C2 (n_123_141) );
AOI211_X1 g_136_137 (.ZN (n_136_137), .A (n_136_139), .B (n_135_135), .C1 (n_131_137), .C2 (n_125_140) );
AOI211_X1 g_134_136 (.ZN (n_134_136), .A (n_138_138), .B (n_137_136), .C1 (n_133_136), .C2 (n_127_139) );
AOI211_X1 g_135_134 (.ZN (n_135_134), .A (n_136_137), .B (n_135_137), .C1 (n_135_135), .C2 (n_129_138) );
AOI211_X1 g_136_136 (.ZN (n_136_136), .A (n_134_136), .B (n_136_139), .C1 (n_137_136), .C2 (n_131_137) );
AOI211_X1 g_138_137 (.ZN (n_138_137), .A (n_135_134), .B (n_138_138), .C1 (n_135_137), .C2 (n_133_136) );
AOI211_X1 g_137_139 (.ZN (n_137_139), .A (n_136_136), .B (n_136_137), .C1 (n_136_139), .C2 (n_135_135) );
AOI211_X1 g_135_138 (.ZN (n_135_138), .A (n_138_137), .B (n_134_136), .C1 (n_138_138), .C2 (n_137_136) );
AOI211_X1 g_133_137 (.ZN (n_133_137), .A (n_137_139), .B (n_135_134), .C1 (n_136_137), .C2 (n_135_137) );
AOI211_X1 g_135_136 (.ZN (n_135_136), .A (n_135_138), .B (n_136_136), .C1 (n_134_136), .C2 (n_136_139) );
AOI211_X1 g_133_135 (.ZN (n_133_135), .A (n_133_137), .B (n_138_137), .C1 (n_135_134), .C2 (n_138_138) );
AOI211_X1 g_131_136 (.ZN (n_131_136), .A (n_135_136), .B (n_137_139), .C1 (n_136_136), .C2 (n_136_137) );
AOI211_X1 g_129_137 (.ZN (n_129_137), .A (n_133_135), .B (n_135_138), .C1 (n_138_137), .C2 (n_134_136) );
AOI211_X1 g_127_138 (.ZN (n_127_138), .A (n_131_136), .B (n_133_137), .C1 (n_137_139), .C2 (n_135_134) );
AOI211_X1 g_125_139 (.ZN (n_125_139), .A (n_129_137), .B (n_135_136), .C1 (n_135_138), .C2 (n_136_136) );
AOI211_X1 g_123_140 (.ZN (n_123_140), .A (n_127_138), .B (n_133_135), .C1 (n_133_137), .C2 (n_138_137) );
AOI211_X1 g_121_141 (.ZN (n_121_141), .A (n_125_139), .B (n_131_136), .C1 (n_135_136), .C2 (n_137_139) );
AOI211_X1 g_119_142 (.ZN (n_119_142), .A (n_123_140), .B (n_129_137), .C1 (n_133_135), .C2 (n_135_138) );
AOI211_X1 g_120_144 (.ZN (n_120_144), .A (n_121_141), .B (n_127_138), .C1 (n_131_136), .C2 (n_133_137) );
AOI211_X1 g_119_146 (.ZN (n_119_146), .A (n_119_142), .B (n_125_139), .C1 (n_129_137), .C2 (n_135_136) );
AOI211_X1 g_118_148 (.ZN (n_118_148), .A (n_120_144), .B (n_123_140), .C1 (n_127_138), .C2 (n_133_135) );
AOI211_X1 g_117_146 (.ZN (n_117_146), .A (n_119_146), .B (n_121_141), .C1 (n_125_139), .C2 (n_131_136) );
AOI211_X1 g_118_144 (.ZN (n_118_144), .A (n_118_148), .B (n_119_142), .C1 (n_123_140), .C2 (n_129_137) );
AOI211_X1 g_120_143 (.ZN (n_120_143), .A (n_117_146), .B (n_120_144), .C1 (n_121_141), .C2 (n_127_138) );
AOI211_X1 g_119_145 (.ZN (n_119_145), .A (n_118_144), .B (n_119_146), .C1 (n_119_142), .C2 (n_125_139) );
AOI211_X1 g_121_146 (.ZN (n_121_146), .A (n_120_143), .B (n_118_148), .C1 (n_120_144), .C2 (n_123_140) );
AOI211_X1 g_122_148 (.ZN (n_122_148), .A (n_119_145), .B (n_117_146), .C1 (n_119_146), .C2 (n_121_141) );
AOI211_X1 g_120_147 (.ZN (n_120_147), .A (n_121_146), .B (n_118_144), .C1 (n_118_148), .C2 (n_119_142) );
AOI211_X1 g_118_146 (.ZN (n_118_146), .A (n_122_148), .B (n_120_143), .C1 (n_117_146), .C2 (n_120_144) );
AOI211_X1 g_119_144 (.ZN (n_119_144), .A (n_120_147), .B (n_119_145), .C1 (n_118_144), .C2 (n_119_146) );
AOI211_X1 g_121_143 (.ZN (n_121_143), .A (n_118_146), .B (n_121_146), .C1 (n_120_143), .C2 (n_118_148) );
AOI211_X1 g_120_145 (.ZN (n_120_145), .A (n_119_144), .B (n_122_148), .C1 (n_119_145), .C2 (n_117_146) );
AOI211_X1 g_122_144 (.ZN (n_122_144), .A (n_121_143), .B (n_120_147), .C1 (n_121_146), .C2 (n_118_144) );
AOI211_X1 g_123_142 (.ZN (n_123_142), .A (n_120_145), .B (n_118_146), .C1 (n_122_148), .C2 (n_120_143) );
AOI211_X1 g_125_141 (.ZN (n_125_141), .A (n_122_144), .B (n_119_144), .C1 (n_120_147), .C2 (n_119_145) );
AOI211_X1 g_127_140 (.ZN (n_127_140), .A (n_123_142), .B (n_121_143), .C1 (n_118_146), .C2 (n_121_146) );
AOI211_X1 g_129_139 (.ZN (n_129_139), .A (n_125_141), .B (n_120_145), .C1 (n_119_144), .C2 (n_122_148) );
AOI211_X1 g_131_138 (.ZN (n_131_138), .A (n_127_140), .B (n_122_144), .C1 (n_121_143), .C2 (n_120_147) );
AOI211_X1 g_130_140 (.ZN (n_130_140), .A (n_129_139), .B (n_123_142), .C1 (n_120_145), .C2 (n_118_146) );
AOI211_X1 g_128_139 (.ZN (n_128_139), .A (n_131_138), .B (n_125_141), .C1 (n_122_144), .C2 (n_119_144) );
AOI211_X1 g_130_138 (.ZN (n_130_138), .A (n_130_140), .B (n_127_140), .C1 (n_123_142), .C2 (n_121_143) );
AOI211_X1 g_132_137 (.ZN (n_132_137), .A (n_128_139), .B (n_129_139), .C1 (n_125_141), .C2 (n_120_145) );
AOI211_X1 g_134_138 (.ZN (n_134_138), .A (n_130_138), .B (n_131_138), .C1 (n_127_140), .C2 (n_122_144) );
AOI211_X1 g_132_139 (.ZN (n_132_139), .A (n_132_137), .B (n_130_140), .C1 (n_129_139), .C2 (n_123_142) );
AOI211_X1 g_134_140 (.ZN (n_134_140), .A (n_134_138), .B (n_128_139), .C1 (n_131_138), .C2 (n_125_141) );
AOI211_X1 g_133_138 (.ZN (n_133_138), .A (n_132_139), .B (n_130_138), .C1 (n_130_140), .C2 (n_127_140) );
AOI211_X1 g_131_139 (.ZN (n_131_139), .A (n_134_140), .B (n_132_137), .C1 (n_128_139), .C2 (n_129_139) );
AOI211_X1 g_129_140 (.ZN (n_129_140), .A (n_133_138), .B (n_134_138), .C1 (n_130_138), .C2 (n_131_138) );
AOI211_X1 g_127_141 (.ZN (n_127_141), .A (n_131_139), .B (n_132_139), .C1 (n_132_137), .C2 (n_130_140) );
AOI211_X1 g_125_142 (.ZN (n_125_142), .A (n_129_140), .B (n_134_140), .C1 (n_134_138), .C2 (n_128_139) );
AOI211_X1 g_126_140 (.ZN (n_126_140), .A (n_127_141), .B (n_133_138), .C1 (n_132_139), .C2 (n_130_138) );
AOI211_X1 g_124_141 (.ZN (n_124_141), .A (n_125_142), .B (n_131_139), .C1 (n_134_140), .C2 (n_132_137) );
AOI211_X1 g_122_142 (.ZN (n_122_142), .A (n_126_140), .B (n_129_140), .C1 (n_133_138), .C2 (n_134_138) );
AOI211_X1 g_121_144 (.ZN (n_121_144), .A (n_124_141), .B (n_127_141), .C1 (n_131_139), .C2 (n_132_139) );
AOI211_X1 g_123_143 (.ZN (n_123_143), .A (n_122_142), .B (n_125_142), .C1 (n_129_140), .C2 (n_134_140) );
AOI211_X1 g_124_145 (.ZN (n_124_145), .A (n_121_144), .B (n_126_140), .C1 (n_127_141), .C2 (n_133_138) );
AOI211_X1 g_122_146 (.ZN (n_122_146), .A (n_123_143), .B (n_124_141), .C1 (n_125_142), .C2 (n_131_139) );
AOI211_X1 g_123_144 (.ZN (n_123_144), .A (n_124_145), .B (n_122_142), .C1 (n_126_140), .C2 (n_129_140) );
AOI211_X1 g_121_145 (.ZN (n_121_145), .A (n_122_146), .B (n_121_144), .C1 (n_124_141), .C2 (n_127_141) );
AOI211_X1 g_123_146 (.ZN (n_123_146), .A (n_123_144), .B (n_123_143), .C1 (n_122_142), .C2 (n_125_142) );
AOI211_X1 g_124_144 (.ZN (n_124_144), .A (n_121_145), .B (n_124_145), .C1 (n_121_144), .C2 (n_126_140) );
AOI211_X1 g_122_143 (.ZN (n_122_143), .A (n_123_146), .B (n_122_146), .C1 (n_123_143), .C2 (n_124_141) );
AOI211_X1 g_124_142 (.ZN (n_124_142), .A (n_124_144), .B (n_123_144), .C1 (n_124_145), .C2 (n_122_142) );
AOI211_X1 g_126_141 (.ZN (n_126_141), .A (n_122_143), .B (n_121_145), .C1 (n_122_146), .C2 (n_121_144) );
AOI211_X1 g_125_143 (.ZN (n_125_143), .A (n_124_142), .B (n_123_146), .C1 (n_123_144), .C2 (n_123_143) );
AOI211_X1 g_127_142 (.ZN (n_127_142), .A (n_126_141), .B (n_124_144), .C1 (n_121_145), .C2 (n_124_145) );
AOI211_X1 g_128_140 (.ZN (n_128_140), .A (n_125_143), .B (n_122_143), .C1 (n_123_146), .C2 (n_122_146) );
AOI211_X1 g_130_139 (.ZN (n_130_139), .A (n_127_142), .B (n_124_142), .C1 (n_124_144), .C2 (n_123_144) );
AOI211_X1 g_132_138 (.ZN (n_132_138), .A (n_128_140), .B (n_126_141), .C1 (n_122_143), .C2 (n_121_145) );
AOI211_X1 g_134_137 (.ZN (n_134_137), .A (n_130_139), .B (n_125_143), .C1 (n_124_142), .C2 (n_123_146) );
AOI211_X1 g_136_138 (.ZN (n_136_138), .A (n_132_138), .B (n_127_142), .C1 (n_126_141), .C2 (n_124_144) );
AOI211_X1 g_134_139 (.ZN (n_134_139), .A (n_134_137), .B (n_128_140), .C1 (n_125_143), .C2 (n_122_143) );
AOI211_X1 g_132_140 (.ZN (n_132_140), .A (n_136_138), .B (n_130_139), .C1 (n_127_142), .C2 (n_124_142) );
AOI211_X1 g_130_141 (.ZN (n_130_141), .A (n_134_139), .B (n_132_138), .C1 (n_128_140), .C2 (n_126_141) );
AOI211_X1 g_128_142 (.ZN (n_128_142), .A (n_132_140), .B (n_134_137), .C1 (n_130_139), .C2 (n_125_143) );
AOI211_X1 g_126_143 (.ZN (n_126_143), .A (n_130_141), .B (n_136_138), .C1 (n_132_138), .C2 (n_127_142) );
AOI211_X1 g_125_145 (.ZN (n_125_145), .A (n_128_142), .B (n_134_139), .C1 (n_134_137), .C2 (n_128_140) );
AOI211_X1 g_124_143 (.ZN (n_124_143), .A (n_126_143), .B (n_132_140), .C1 (n_136_138), .C2 (n_130_139) );
AOI211_X1 g_123_145 (.ZN (n_123_145), .A (n_125_145), .B (n_130_141), .C1 (n_134_139), .C2 (n_132_138) );
AOI211_X1 g_124_147 (.ZN (n_124_147), .A (n_124_143), .B (n_128_142), .C1 (n_132_140), .C2 (n_134_137) );
AOI211_X1 g_126_148 (.ZN (n_126_148), .A (n_123_145), .B (n_126_143), .C1 (n_130_141), .C2 (n_136_138) );
AOI211_X1 g_125_146 (.ZN (n_125_146), .A (n_124_147), .B (n_125_145), .C1 (n_128_142), .C2 (n_134_139) );
AOI211_X1 g_126_144 (.ZN (n_126_144), .A (n_126_148), .B (n_124_143), .C1 (n_126_143), .C2 (n_132_140) );
AOI211_X1 g_127_146 (.ZN (n_127_146), .A (n_125_146), .B (n_123_145), .C1 (n_125_145), .C2 (n_130_141) );
AOI211_X1 g_129_147 (.ZN (n_129_147), .A (n_126_144), .B (n_124_147), .C1 (n_124_143), .C2 (n_128_142) );
AOI211_X1 g_131_146 (.ZN (n_131_146), .A (n_127_146), .B (n_126_148), .C1 (n_123_145), .C2 (n_126_143) );
AOI211_X1 g_133_145 (.ZN (n_133_145), .A (n_129_147), .B (n_125_146), .C1 (n_124_147), .C2 (n_125_145) );
AOI211_X1 g_135_144 (.ZN (n_135_144), .A (n_131_146), .B (n_126_144), .C1 (n_126_148), .C2 (n_124_143) );
AOI211_X1 g_136_142 (.ZN (n_136_142), .A (n_133_145), .B (n_127_146), .C1 (n_125_146), .C2 (n_123_145) );
AOI211_X1 g_137_140 (.ZN (n_137_140), .A (n_135_144), .B (n_129_147), .C1 (n_126_144), .C2 (n_124_147) );
AOI211_X1 g_135_139 (.ZN (n_135_139), .A (n_136_142), .B (n_131_146), .C1 (n_127_146), .C2 (n_126_148) );
AOI211_X1 g_136_141 (.ZN (n_136_141), .A (n_137_140), .B (n_133_145), .C1 (n_129_147), .C2 (n_125_146) );
AOI211_X1 g_138_142 (.ZN (n_138_142), .A (n_135_139), .B (n_135_144), .C1 (n_131_146), .C2 (n_126_144) );
AOI211_X1 g_137_144 (.ZN (n_137_144), .A (n_136_141), .B (n_136_142), .C1 (n_133_145), .C2 (n_127_146) );
AOI211_X1 g_135_143 (.ZN (n_135_143), .A (n_138_142), .B (n_137_140), .C1 (n_135_144), .C2 (n_129_147) );
AOI211_X1 g_134_141 (.ZN (n_134_141), .A (n_137_144), .B (n_135_139), .C1 (n_136_142), .C2 (n_131_146) );
AOI211_X1 g_133_139 (.ZN (n_133_139), .A (n_135_143), .B (n_136_141), .C1 (n_137_140), .C2 (n_133_145) );
AOI211_X1 g_135_140 (.ZN (n_135_140), .A (n_134_141), .B (n_138_142), .C1 (n_135_139), .C2 (n_135_144) );
AOI211_X1 g_133_141 (.ZN (n_133_141), .A (n_133_139), .B (n_137_144), .C1 (n_136_141), .C2 (n_136_142) );
AOI211_X1 g_131_140 (.ZN (n_131_140), .A (n_135_140), .B (n_135_143), .C1 (n_138_142), .C2 (n_137_140) );
AOI211_X1 g_129_141 (.ZN (n_129_141), .A (n_133_141), .B (n_134_141), .C1 (n_137_144), .C2 (n_135_139) );
AOI211_X1 g_131_142 (.ZN (n_131_142), .A (n_131_140), .B (n_133_139), .C1 (n_135_143), .C2 (n_136_141) );
AOI211_X1 g_133_143 (.ZN (n_133_143), .A (n_129_141), .B (n_135_140), .C1 (n_134_141), .C2 (n_138_142) );
AOI211_X1 g_132_141 (.ZN (n_132_141), .A (n_131_142), .B (n_133_141), .C1 (n_133_139), .C2 (n_137_144) );
AOI211_X1 g_134_142 (.ZN (n_134_142), .A (n_133_143), .B (n_131_140), .C1 (n_135_140), .C2 (n_135_143) );
AOI211_X1 g_133_140 (.ZN (n_133_140), .A (n_132_141), .B (n_129_141), .C1 (n_133_141), .C2 (n_134_141) );
AOI211_X1 g_135_141 (.ZN (n_135_141), .A (n_134_142), .B (n_131_142), .C1 (n_131_140), .C2 (n_133_139) );
AOI211_X1 g_136_143 (.ZN (n_136_143), .A (n_133_140), .B (n_133_143), .C1 (n_129_141), .C2 (n_135_140) );
AOI211_X1 g_135_145 (.ZN (n_135_145), .A (n_135_141), .B (n_132_141), .C1 (n_131_142), .C2 (n_133_141) );
AOI211_X1 g_134_143 (.ZN (n_134_143), .A (n_136_143), .B (n_134_142), .C1 (n_133_143), .C2 (n_131_140) );
AOI211_X1 g_132_142 (.ZN (n_132_142), .A (n_135_145), .B (n_133_140), .C1 (n_132_141), .C2 (n_129_141) );
AOI211_X1 g_133_144 (.ZN (n_133_144), .A (n_134_143), .B (n_135_141), .C1 (n_134_142), .C2 (n_131_142) );
AOI211_X1 g_131_143 (.ZN (n_131_143), .A (n_132_142), .B (n_136_143), .C1 (n_133_140), .C2 (n_133_143) );
AOI211_X1 g_133_142 (.ZN (n_133_142), .A (n_133_144), .B (n_135_145), .C1 (n_135_141), .C2 (n_132_141) );
AOI211_X1 g_131_141 (.ZN (n_131_141), .A (n_131_143), .B (n_134_143), .C1 (n_136_143), .C2 (n_134_142) );
AOI211_X1 g_129_142 (.ZN (n_129_142), .A (n_133_142), .B (n_132_142), .C1 (n_135_145), .C2 (n_133_140) );
AOI211_X1 g_128_144 (.ZN (n_128_144), .A (n_131_141), .B (n_133_144), .C1 (n_134_143), .C2 (n_135_141) );
AOI211_X1 g_130_143 (.ZN (n_130_143), .A (n_129_142), .B (n_131_143), .C1 (n_132_142), .C2 (n_136_143) );
AOI211_X1 g_132_144 (.ZN (n_132_144), .A (n_128_144), .B (n_133_142), .C1 (n_133_144), .C2 (n_135_145) );
AOI211_X1 g_130_145 (.ZN (n_130_145), .A (n_130_143), .B (n_131_141), .C1 (n_131_143), .C2 (n_134_143) );
AOI211_X1 g_131_147 (.ZN (n_131_147), .A (n_132_144), .B (n_129_142), .C1 (n_133_142), .C2 (n_132_142) );
AOI211_X1 g_133_146 (.ZN (n_133_146), .A (n_130_145), .B (n_128_144), .C1 (n_131_141), .C2 (n_133_144) );
AOI211_X1 g_134_144 (.ZN (n_134_144), .A (n_131_147), .B (n_130_143), .C1 (n_129_142), .C2 (n_131_143) );
AOI211_X1 g_132_145 (.ZN (n_132_145), .A (n_133_146), .B (n_132_144), .C1 (n_128_144), .C2 (n_133_142) );
AOI211_X1 g_130_144 (.ZN (n_130_144), .A (n_134_144), .B (n_130_145), .C1 (n_130_143), .C2 (n_131_141) );
AOI211_X1 g_132_143 (.ZN (n_132_143), .A (n_132_145), .B (n_131_147), .C1 (n_132_144), .C2 (n_129_142) );
AOI211_X1 g_131_145 (.ZN (n_131_145), .A (n_130_144), .B (n_133_146), .C1 (n_130_145), .C2 (n_128_144) );
AOI211_X1 g_129_146 (.ZN (n_129_146), .A (n_132_143), .B (n_134_144), .C1 (n_131_147), .C2 (n_130_143) );
AOI211_X1 g_127_145 (.ZN (n_127_145), .A (n_131_145), .B (n_132_145), .C1 (n_133_146), .C2 (n_132_144) );
AOI211_X1 g_129_144 (.ZN (n_129_144), .A (n_129_146), .B (n_130_144), .C1 (n_134_144), .C2 (n_130_145) );
AOI211_X1 g_130_142 (.ZN (n_130_142), .A (n_127_145), .B (n_132_143), .C1 (n_132_145), .C2 (n_131_147) );
AOI211_X1 g_128_143 (.ZN (n_128_143), .A (n_129_144), .B (n_131_145), .C1 (n_130_144), .C2 (n_133_146) );
AOI211_X1 g_126_142 (.ZN (n_126_142), .A (n_130_142), .B (n_129_146), .C1 (n_132_143), .C2 (n_134_144) );
AOI211_X1 g_128_141 (.ZN (n_128_141), .A (n_128_143), .B (n_127_145), .C1 (n_131_145), .C2 (n_132_145) );
AOI211_X1 g_127_143 (.ZN (n_127_143), .A (n_126_142), .B (n_129_144), .C1 (n_129_146), .C2 (n_130_144) );
AOI211_X1 g_125_144 (.ZN (n_125_144), .A (n_128_141), .B (n_130_142), .C1 (n_127_145), .C2 (n_132_143) );
AOI211_X1 g_126_146 (.ZN (n_126_146), .A (n_127_143), .B (n_128_143), .C1 (n_129_144), .C2 (n_131_145) );
AOI211_X1 g_128_145 (.ZN (n_128_145), .A (n_125_144), .B (n_126_142), .C1 (n_130_142), .C2 (n_129_146) );
AOI211_X1 g_129_143 (.ZN (n_129_143), .A (n_126_146), .B (n_128_141), .C1 (n_128_143), .C2 (n_127_145) );
AOI211_X1 g_127_144 (.ZN (n_127_144), .A (n_128_145), .B (n_127_143), .C1 (n_126_142), .C2 (n_129_144) );
AOI211_X1 g_129_145 (.ZN (n_129_145), .A (n_129_143), .B (n_125_144), .C1 (n_128_141), .C2 (n_130_142) );
AOI211_X1 g_131_144 (.ZN (n_131_144), .A (n_127_144), .B (n_126_146), .C1 (n_127_143), .C2 (n_128_143) );
AOI211_X1 g_130_146 (.ZN (n_130_146), .A (n_129_145), .B (n_128_145), .C1 (n_125_144), .C2 (n_126_142) );
AOI211_X1 g_128_147 (.ZN (n_128_147), .A (n_131_144), .B (n_129_143), .C1 (n_126_146), .C2 (n_128_141) );
endmodule
