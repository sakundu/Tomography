module mesh(clk, in, out);
input clk, in;
output out;
AOI211_X1 g_4_4 (.ZN (n_4_4) );
AOI211_X1 g_5_2 (.ZN (n_5_2) );
AOI211_X1 g_7_1 (.ZN (n_7_1), .A (n_4_4) );
AOI211_X1 g_9_2 (.ZN (n_9_2), .A (n_5_2) );
AOI211_X1 g_11_1 (.ZN (n_11_1), .A (n_7_1) );
AOI211_X1 g_13_2 (.ZN (n_13_2), .A (n_9_2), .B (n_4_4) );
AOI211_X1 g_15_1 (.ZN (n_15_1), .A (n_11_1), .B (n_5_2) );
AOI211_X1 g_17_2 (.ZN (n_17_2), .A (n_13_2), .B (n_7_1), .C1 (n_4_4) );
AOI211_X1 g_19_1 (.ZN (n_19_1), .A (n_15_1), .B (n_9_2), .C1 (n_5_2) );
AOI211_X1 g_21_2 (.ZN (n_21_2), .A (n_17_2), .B (n_11_1), .C1 (n_7_1) );
AOI211_X1 g_23_1 (.ZN (n_23_1), .A (n_19_1), .B (n_13_2), .C1 (n_9_2), .C2 (n_4_4) );
AOI211_X1 g_25_2 (.ZN (n_25_2), .A (n_21_2), .B (n_15_1), .C1 (n_11_1), .C2 (n_5_2) );
AOI211_X1 g_27_1 (.ZN (n_27_1), .A (n_23_1), .B (n_17_2), .C1 (n_13_2), .C2 (n_7_1) );
AOI211_X1 g_29_2 (.ZN (n_29_2), .A (n_25_2), .B (n_19_1), .C1 (n_15_1), .C2 (n_9_2) );
AOI211_X1 g_31_1 (.ZN (n_31_1), .A (n_27_1), .B (n_21_2), .C1 (n_17_2), .C2 (n_11_1) );
AOI211_X1 g_33_2 (.ZN (n_33_2), .A (n_29_2), .B (n_23_1), .C1 (n_19_1), .C2 (n_13_2) );
AOI211_X1 g_35_1 (.ZN (n_35_1), .A (n_31_1), .B (n_25_2), .C1 (n_21_2), .C2 (n_15_1) );
AOI211_X1 g_37_2 (.ZN (n_37_2), .A (n_33_2), .B (n_27_1), .C1 (n_23_1), .C2 (n_17_2) );
AOI211_X1 g_39_1 (.ZN (n_39_1), .A (n_35_1), .B (n_29_2), .C1 (n_25_2), .C2 (n_19_1) );
AOI211_X1 g_41_2 (.ZN (n_41_2), .A (n_37_2), .B (n_31_1), .C1 (n_27_1), .C2 (n_21_2) );
AOI211_X1 g_43_1 (.ZN (n_43_1), .A (n_39_1), .B (n_33_2), .C1 (n_29_2), .C2 (n_23_1) );
AOI211_X1 g_45_2 (.ZN (n_45_2), .A (n_41_2), .B (n_35_1), .C1 (n_31_1), .C2 (n_25_2) );
AOI211_X1 g_47_1 (.ZN (n_47_1), .A (n_43_1), .B (n_37_2), .C1 (n_33_2), .C2 (n_27_1) );
AOI211_X1 g_49_2 (.ZN (n_49_2), .A (n_45_2), .B (n_39_1), .C1 (n_35_1), .C2 (n_29_2) );
AOI211_X1 g_51_1 (.ZN (n_51_1), .A (n_47_1), .B (n_41_2), .C1 (n_37_2), .C2 (n_31_1) );
AOI211_X1 g_53_2 (.ZN (n_53_2), .A (n_49_2), .B (n_43_1), .C1 (n_39_1), .C2 (n_33_2) );
AOI211_X1 g_55_1 (.ZN (n_55_1), .A (n_51_1), .B (n_45_2), .C1 (n_41_2), .C2 (n_35_1) );
AOI211_X1 g_57_2 (.ZN (n_57_2), .A (n_53_2), .B (n_47_1), .C1 (n_43_1), .C2 (n_37_2) );
AOI211_X1 g_59_1 (.ZN (n_59_1), .A (n_55_1), .B (n_49_2), .C1 (n_45_2), .C2 (n_39_1) );
AOI211_X1 g_61_2 (.ZN (n_61_2), .A (n_57_2), .B (n_51_1), .C1 (n_47_1), .C2 (n_41_2) );
AOI211_X1 g_63_1 (.ZN (n_63_1), .A (n_59_1), .B (n_53_2), .C1 (n_49_2), .C2 (n_43_1) );
AOI211_X1 g_65_2 (.ZN (n_65_2), .A (n_61_2), .B (n_55_1), .C1 (n_51_1), .C2 (n_45_2) );
AOI211_X1 g_67_1 (.ZN (n_67_1), .A (n_63_1), .B (n_57_2), .C1 (n_53_2), .C2 (n_47_1) );
AOI211_X1 g_69_2 (.ZN (n_69_2), .A (n_65_2), .B (n_59_1), .C1 (n_55_1), .C2 (n_49_2) );
AOI211_X1 g_71_1 (.ZN (n_71_1), .A (n_67_1), .B (n_61_2), .C1 (n_57_2), .C2 (n_51_1) );
AOI211_X1 g_73_2 (.ZN (n_73_2), .A (n_69_2), .B (n_63_1), .C1 (n_59_1), .C2 (n_53_2) );
AOI211_X1 g_75_1 (.ZN (n_75_1), .A (n_71_1), .B (n_65_2), .C1 (n_61_2), .C2 (n_55_1) );
AOI211_X1 g_77_2 (.ZN (n_77_2), .A (n_73_2), .B (n_67_1), .C1 (n_63_1), .C2 (n_57_2) );
AOI211_X1 g_79_1 (.ZN (n_79_1), .A (n_75_1), .B (n_69_2), .C1 (n_65_2), .C2 (n_59_1) );
AOI211_X1 g_81_2 (.ZN (n_81_2), .A (n_77_2), .B (n_71_1), .C1 (n_67_1), .C2 (n_61_2) );
AOI211_X1 g_83_1 (.ZN (n_83_1), .A (n_79_1), .B (n_73_2), .C1 (n_69_2), .C2 (n_63_1) );
AOI211_X1 g_85_2 (.ZN (n_85_2), .A (n_81_2), .B (n_75_1), .C1 (n_71_1), .C2 (n_65_2) );
AOI211_X1 g_87_1 (.ZN (n_87_1), .A (n_83_1), .B (n_77_2), .C1 (n_73_2), .C2 (n_67_1) );
AOI211_X1 g_89_2 (.ZN (n_89_2), .A (n_85_2), .B (n_79_1), .C1 (n_75_1), .C2 (n_69_2) );
AOI211_X1 g_91_1 (.ZN (n_91_1), .A (n_87_1), .B (n_81_2), .C1 (n_77_2), .C2 (n_71_1) );
AOI211_X1 g_93_2 (.ZN (n_93_2), .A (n_89_2), .B (n_83_1), .C1 (n_79_1), .C2 (n_73_2) );
AOI211_X1 g_95_1 (.ZN (n_95_1), .A (n_91_1), .B (n_85_2), .C1 (n_81_2), .C2 (n_75_1) );
AOI211_X1 g_97_2 (.ZN (n_97_2), .A (n_93_2), .B (n_87_1), .C1 (n_83_1), .C2 (n_77_2) );
AOI211_X1 g_99_1 (.ZN (n_99_1), .A (n_95_1), .B (n_89_2), .C1 (n_85_2), .C2 (n_79_1) );
AOI211_X1 g_100_3 (.ZN (n_100_3), .A (n_97_2), .B (n_91_1), .C1 (n_87_1), .C2 (n_81_2) );
AOI211_X1 g_98_2 (.ZN (n_98_2), .A (n_99_1), .B (n_93_2), .C1 (n_89_2), .C2 (n_83_1) );
AOI211_X1 g_100_1 (.ZN (n_100_1), .A (n_100_3), .B (n_95_1), .C1 (n_91_1), .C2 (n_85_2) );
AOI211_X1 g_99_3 (.ZN (n_99_3), .A (n_98_2), .B (n_97_2), .C1 (n_93_2), .C2 (n_87_1) );
AOI211_X1 g_98_1 (.ZN (n_98_1), .A (n_100_1), .B (n_99_1), .C1 (n_95_1), .C2 (n_89_2) );
AOI211_X1 g_100_2 (.ZN (n_100_2), .A (n_99_3), .B (n_100_3), .C1 (n_97_2), .C2 (n_91_1) );
AOI211_X1 g_99_4 (.ZN (n_99_4), .A (n_98_1), .B (n_98_2), .C1 (n_99_1), .C2 (n_93_2) );
AOI211_X1 g_100_6 (.ZN (n_100_6), .A (n_100_2), .B (n_100_1), .C1 (n_100_3), .C2 (n_95_1) );
AOI211_X1 g_99_8 (.ZN (n_99_8), .A (n_99_4), .B (n_99_3), .C1 (n_98_2), .C2 (n_97_2) );
AOI211_X1 g_100_10 (.ZN (n_100_10), .A (n_100_6), .B (n_98_1), .C1 (n_100_1), .C2 (n_99_1) );
AOI211_X1 g_99_12 (.ZN (n_99_12), .A (n_99_8), .B (n_100_2), .C1 (n_99_3), .C2 (n_100_3) );
AOI211_X1 g_100_14 (.ZN (n_100_14), .A (n_100_10), .B (n_99_4), .C1 (n_98_1), .C2 (n_98_2) );
AOI211_X1 g_99_16 (.ZN (n_99_16), .A (n_99_12), .B (n_100_6), .C1 (n_100_2), .C2 (n_100_1) );
AOI211_X1 g_100_18 (.ZN (n_100_18), .A (n_100_14), .B (n_99_8), .C1 (n_99_4), .C2 (n_99_3) );
AOI211_X1 g_99_20 (.ZN (n_99_20), .A (n_99_16), .B (n_100_10), .C1 (n_100_6), .C2 (n_98_1) );
AOI211_X1 g_100_22 (.ZN (n_100_22), .A (n_100_18), .B (n_99_12), .C1 (n_99_8), .C2 (n_100_2) );
AOI211_X1 g_99_24 (.ZN (n_99_24), .A (n_99_20), .B (n_100_14), .C1 (n_100_10), .C2 (n_99_4) );
AOI211_X1 g_100_26 (.ZN (n_100_26), .A (n_100_22), .B (n_99_16), .C1 (n_99_12), .C2 (n_100_6) );
AOI211_X1 g_99_28 (.ZN (n_99_28), .A (n_99_24), .B (n_100_18), .C1 (n_100_14), .C2 (n_99_8) );
AOI211_X1 g_100_30 (.ZN (n_100_30), .A (n_100_26), .B (n_99_20), .C1 (n_99_16), .C2 (n_100_10) );
AOI211_X1 g_99_32 (.ZN (n_99_32), .A (n_99_28), .B (n_100_22), .C1 (n_100_18), .C2 (n_99_12) );
AOI211_X1 g_100_34 (.ZN (n_100_34), .A (n_100_30), .B (n_99_24), .C1 (n_99_20), .C2 (n_100_14) );
AOI211_X1 g_99_36 (.ZN (n_99_36), .A (n_99_32), .B (n_100_26), .C1 (n_100_22), .C2 (n_99_16) );
AOI211_X1 g_100_38 (.ZN (n_100_38), .A (n_100_34), .B (n_99_28), .C1 (n_99_24), .C2 (n_100_18) );
AOI211_X1 g_99_40 (.ZN (n_99_40), .A (n_99_36), .B (n_100_30), .C1 (n_100_26), .C2 (n_99_20) );
AOI211_X1 g_100_42 (.ZN (n_100_42), .A (n_100_38), .B (n_99_32), .C1 (n_99_28), .C2 (n_100_22) );
AOI211_X1 g_99_44 (.ZN (n_99_44), .A (n_99_40), .B (n_100_34), .C1 (n_100_30), .C2 (n_99_24) );
AOI211_X1 g_100_46 (.ZN (n_100_46), .A (n_100_42), .B (n_99_36), .C1 (n_99_32), .C2 (n_100_26) );
AOI211_X1 g_99_48 (.ZN (n_99_48), .A (n_99_44), .B (n_100_38), .C1 (n_100_34), .C2 (n_99_28) );
AOI211_X1 g_100_50 (.ZN (n_100_50), .A (n_100_46), .B (n_99_40), .C1 (n_99_36), .C2 (n_100_30) );
AOI211_X1 g_99_52 (.ZN (n_99_52), .A (n_99_48), .B (n_100_42), .C1 (n_100_38), .C2 (n_99_32) );
AOI211_X1 g_100_54 (.ZN (n_100_54), .A (n_100_50), .B (n_99_44), .C1 (n_99_40), .C2 (n_100_34) );
AOI211_X1 g_99_56 (.ZN (n_99_56), .A (n_99_52), .B (n_100_46), .C1 (n_100_42), .C2 (n_99_36) );
AOI211_X1 g_100_58 (.ZN (n_100_58), .A (n_100_54), .B (n_99_48), .C1 (n_99_44), .C2 (n_100_38) );
AOI211_X1 g_99_60 (.ZN (n_99_60), .A (n_99_56), .B (n_100_50), .C1 (n_100_46), .C2 (n_99_40) );
AOI211_X1 g_100_62 (.ZN (n_100_62), .A (n_100_58), .B (n_99_52), .C1 (n_99_48), .C2 (n_100_42) );
AOI211_X1 g_99_64 (.ZN (n_99_64), .A (n_99_60), .B (n_100_54), .C1 (n_100_50), .C2 (n_99_44) );
AOI211_X1 g_100_66 (.ZN (n_100_66), .A (n_100_62), .B (n_99_56), .C1 (n_99_52), .C2 (n_100_46) );
AOI211_X1 g_99_68 (.ZN (n_99_68), .A (n_99_64), .B (n_100_58), .C1 (n_100_54), .C2 (n_99_48) );
AOI211_X1 g_100_70 (.ZN (n_100_70), .A (n_100_66), .B (n_99_60), .C1 (n_99_56), .C2 (n_100_50) );
AOI211_X1 g_99_72 (.ZN (n_99_72), .A (n_99_68), .B (n_100_62), .C1 (n_100_58), .C2 (n_99_52) );
AOI211_X1 g_100_74 (.ZN (n_100_74), .A (n_100_70), .B (n_99_64), .C1 (n_99_60), .C2 (n_100_54) );
AOI211_X1 g_99_76 (.ZN (n_99_76), .A (n_99_72), .B (n_100_66), .C1 (n_100_62), .C2 (n_99_56) );
AOI211_X1 g_100_78 (.ZN (n_100_78), .A (n_100_74), .B (n_99_68), .C1 (n_99_64), .C2 (n_100_58) );
AOI211_X1 g_99_80 (.ZN (n_99_80), .A (n_99_76), .B (n_100_70), .C1 (n_100_66), .C2 (n_99_60) );
AOI211_X1 g_100_82 (.ZN (n_100_82), .A (n_100_78), .B (n_99_72), .C1 (n_99_68), .C2 (n_100_62) );
AOI211_X1 g_99_84 (.ZN (n_99_84), .A (n_99_80), .B (n_100_74), .C1 (n_100_70), .C2 (n_99_64) );
AOI211_X1 g_100_86 (.ZN (n_100_86), .A (n_100_82), .B (n_99_76), .C1 (n_99_72), .C2 (n_100_66) );
AOI211_X1 g_99_88 (.ZN (n_99_88), .A (n_99_84), .B (n_100_78), .C1 (n_100_74), .C2 (n_99_68) );
AOI211_X1 g_100_90 (.ZN (n_100_90), .A (n_100_86), .B (n_99_80), .C1 (n_99_76), .C2 (n_100_70) );
AOI211_X1 g_99_92 (.ZN (n_99_92), .A (n_99_88), .B (n_100_82), .C1 (n_100_78), .C2 (n_99_72) );
AOI211_X1 g_100_94 (.ZN (n_100_94), .A (n_100_90), .B (n_99_84), .C1 (n_99_80), .C2 (n_100_74) );
AOI211_X1 g_99_96 (.ZN (n_99_96), .A (n_99_92), .B (n_100_86), .C1 (n_100_82), .C2 (n_99_76) );
AOI211_X1 g_100_98 (.ZN (n_100_98), .A (n_100_94), .B (n_99_88), .C1 (n_99_84), .C2 (n_100_78) );
AOI211_X1 g_99_100 (.ZN (n_99_100), .A (n_99_96), .B (n_100_90), .C1 (n_100_86), .C2 (n_99_80) );
AOI211_X1 g_97_99 (.ZN (n_97_99), .A (n_100_98), .B (n_99_92), .C1 (n_99_88), .C2 (n_100_82) );
AOI211_X1 g_95_100 (.ZN (n_95_100), .A (n_99_100), .B (n_100_94), .C1 (n_100_90), .C2 (n_99_84) );
AOI211_X1 g_93_99 (.ZN (n_93_99), .A (n_97_99), .B (n_99_96), .C1 (n_99_92), .C2 (n_100_86) );
AOI211_X1 g_91_100 (.ZN (n_91_100), .A (n_95_100), .B (n_100_98), .C1 (n_100_94), .C2 (n_99_88) );
AOI211_X1 g_89_99 (.ZN (n_89_99), .A (n_93_99), .B (n_99_100), .C1 (n_99_96), .C2 (n_100_90) );
AOI211_X1 g_87_100 (.ZN (n_87_100), .A (n_91_100), .B (n_97_99), .C1 (n_100_98), .C2 (n_99_92) );
AOI211_X1 g_85_99 (.ZN (n_85_99), .A (n_89_99), .B (n_95_100), .C1 (n_99_100), .C2 (n_100_94) );
AOI211_X1 g_83_100 (.ZN (n_83_100), .A (n_87_100), .B (n_93_99), .C1 (n_97_99), .C2 (n_99_96) );
AOI211_X1 g_81_99 (.ZN (n_81_99), .A (n_85_99), .B (n_91_100), .C1 (n_95_100), .C2 (n_100_98) );
AOI211_X1 g_79_100 (.ZN (n_79_100), .A (n_83_100), .B (n_89_99), .C1 (n_93_99), .C2 (n_99_100) );
AOI211_X1 g_77_99 (.ZN (n_77_99), .A (n_81_99), .B (n_87_100), .C1 (n_91_100), .C2 (n_97_99) );
AOI211_X1 g_75_100 (.ZN (n_75_100), .A (n_79_100), .B (n_85_99), .C1 (n_89_99), .C2 (n_95_100) );
AOI211_X1 g_73_99 (.ZN (n_73_99), .A (n_77_99), .B (n_83_100), .C1 (n_87_100), .C2 (n_93_99) );
AOI211_X1 g_71_100 (.ZN (n_71_100), .A (n_75_100), .B (n_81_99), .C1 (n_85_99), .C2 (n_91_100) );
AOI211_X1 g_69_99 (.ZN (n_69_99), .A (n_73_99), .B (n_79_100), .C1 (n_83_100), .C2 (n_89_99) );
AOI211_X1 g_67_100 (.ZN (n_67_100), .A (n_71_100), .B (n_77_99), .C1 (n_81_99), .C2 (n_87_100) );
AOI211_X1 g_65_99 (.ZN (n_65_99), .A (n_69_99), .B (n_75_100), .C1 (n_79_100), .C2 (n_85_99) );
AOI211_X1 g_63_100 (.ZN (n_63_100), .A (n_67_100), .B (n_73_99), .C1 (n_77_99), .C2 (n_83_100) );
AOI211_X1 g_61_99 (.ZN (n_61_99), .A (n_65_99), .B (n_71_100), .C1 (n_75_100), .C2 (n_81_99) );
AOI211_X1 g_59_100 (.ZN (n_59_100), .A (n_63_100), .B (n_69_99), .C1 (n_73_99), .C2 (n_79_100) );
AOI211_X1 g_57_99 (.ZN (n_57_99), .A (n_61_99), .B (n_67_100), .C1 (n_71_100), .C2 (n_77_99) );
AOI211_X1 g_55_100 (.ZN (n_55_100), .A (n_59_100), .B (n_65_99), .C1 (n_69_99), .C2 (n_75_100) );
AOI211_X1 g_53_99 (.ZN (n_53_99), .A (n_57_99), .B (n_63_100), .C1 (n_67_100), .C2 (n_73_99) );
AOI211_X1 g_51_100 (.ZN (n_51_100), .A (n_55_100), .B (n_61_99), .C1 (n_65_99), .C2 (n_71_100) );
AOI211_X1 g_49_99 (.ZN (n_49_99), .A (n_53_99), .B (n_59_100), .C1 (n_63_100), .C2 (n_69_99) );
AOI211_X1 g_47_100 (.ZN (n_47_100), .A (n_51_100), .B (n_57_99), .C1 (n_61_99), .C2 (n_67_100) );
AOI211_X1 g_45_99 (.ZN (n_45_99), .A (n_49_99), .B (n_55_100), .C1 (n_59_100), .C2 (n_65_99) );
AOI211_X1 g_43_100 (.ZN (n_43_100), .A (n_47_100), .B (n_53_99), .C1 (n_57_99), .C2 (n_63_100) );
AOI211_X1 g_41_99 (.ZN (n_41_99), .A (n_45_99), .B (n_51_100), .C1 (n_55_100), .C2 (n_61_99) );
AOI211_X1 g_39_100 (.ZN (n_39_100), .A (n_43_100), .B (n_49_99), .C1 (n_53_99), .C2 (n_59_100) );
AOI211_X1 g_37_99 (.ZN (n_37_99), .A (n_41_99), .B (n_47_100), .C1 (n_51_100), .C2 (n_57_99) );
AOI211_X1 g_35_100 (.ZN (n_35_100), .A (n_39_100), .B (n_45_99), .C1 (n_49_99), .C2 (n_55_100) );
AOI211_X1 g_33_99 (.ZN (n_33_99), .A (n_37_99), .B (n_43_100), .C1 (n_47_100), .C2 (n_53_99) );
AOI211_X1 g_31_100 (.ZN (n_31_100), .A (n_35_100), .B (n_41_99), .C1 (n_45_99), .C2 (n_51_100) );
AOI211_X1 g_29_99 (.ZN (n_29_99), .A (n_33_99), .B (n_39_100), .C1 (n_43_100), .C2 (n_49_99) );
AOI211_X1 g_27_100 (.ZN (n_27_100), .A (n_31_100), .B (n_37_99), .C1 (n_41_99), .C2 (n_47_100) );
AOI211_X1 g_25_99 (.ZN (n_25_99), .A (n_29_99), .B (n_35_100), .C1 (n_39_100), .C2 (n_45_99) );
AOI211_X1 g_23_100 (.ZN (n_23_100), .A (n_27_100), .B (n_33_99), .C1 (n_37_99), .C2 (n_43_100) );
AOI211_X1 g_21_99 (.ZN (n_21_99), .A (n_25_99), .B (n_31_100), .C1 (n_35_100), .C2 (n_41_99) );
AOI211_X1 g_19_100 (.ZN (n_19_100), .A (n_23_100), .B (n_29_99), .C1 (n_33_99), .C2 (n_39_100) );
AOI211_X1 g_17_99 (.ZN (n_17_99), .A (n_21_99), .B (n_27_100), .C1 (n_31_100), .C2 (n_37_99) );
AOI211_X1 g_15_100 (.ZN (n_15_100), .A (n_19_100), .B (n_25_99), .C1 (n_29_99), .C2 (n_35_100) );
AOI211_X1 g_13_99 (.ZN (n_13_99), .A (n_17_99), .B (n_23_100), .C1 (n_27_100), .C2 (n_33_99) );
AOI211_X1 g_11_100 (.ZN (n_11_100), .A (n_15_100), .B (n_21_99), .C1 (n_25_99), .C2 (n_31_100) );
AOI211_X1 g_9_99 (.ZN (n_9_99), .A (n_13_99), .B (n_19_100), .C1 (n_23_100), .C2 (n_29_99) );
AOI211_X1 g_7_100 (.ZN (n_7_100), .A (n_11_100), .B (n_17_99), .C1 (n_21_99), .C2 (n_27_100) );
AOI211_X1 g_5_99 (.ZN (n_5_99), .A (n_9_99), .B (n_15_100), .C1 (n_19_100), .C2 (n_25_99) );
AOI211_X1 g_3_100 (.ZN (n_3_100), .A (n_7_100), .B (n_13_99), .C1 (n_17_99), .C2 (n_23_100) );
AOI211_X1 g_1_99 (.ZN (n_1_99), .A (n_5_99), .B (n_11_100), .C1 (n_15_100), .C2 (n_21_99) );
AOI211_X1 g_2_97 (.ZN (n_2_97), .A (n_3_100), .B (n_9_99), .C1 (n_13_99), .C2 (n_19_100) );
AOI211_X1 g_1_95 (.ZN (n_1_95), .A (n_1_99), .B (n_7_100), .C1 (n_11_100), .C2 (n_17_99) );
AOI211_X1 g_2_93 (.ZN (n_2_93), .A (n_2_97), .B (n_5_99), .C1 (n_9_99), .C2 (n_15_100) );
AOI211_X1 g_1_91 (.ZN (n_1_91), .A (n_1_95), .B (n_3_100), .C1 (n_7_100), .C2 (n_13_99) );
AOI211_X1 g_2_89 (.ZN (n_2_89), .A (n_2_93), .B (n_1_99), .C1 (n_5_99), .C2 (n_11_100) );
AOI211_X1 g_1_87 (.ZN (n_1_87), .A (n_1_91), .B (n_2_97), .C1 (n_3_100), .C2 (n_9_99) );
AOI211_X1 g_2_85 (.ZN (n_2_85), .A (n_2_89), .B (n_1_95), .C1 (n_1_99), .C2 (n_7_100) );
AOI211_X1 g_1_83 (.ZN (n_1_83), .A (n_1_87), .B (n_2_93), .C1 (n_2_97), .C2 (n_5_99) );
AOI211_X1 g_2_81 (.ZN (n_2_81), .A (n_2_85), .B (n_1_91), .C1 (n_1_95), .C2 (n_3_100) );
AOI211_X1 g_1_79 (.ZN (n_1_79), .A (n_1_83), .B (n_2_89), .C1 (n_2_93), .C2 (n_1_99) );
AOI211_X1 g_2_77 (.ZN (n_2_77), .A (n_2_81), .B (n_1_87), .C1 (n_1_91), .C2 (n_2_97) );
AOI211_X1 g_1_75 (.ZN (n_1_75), .A (n_1_79), .B (n_2_85), .C1 (n_2_89), .C2 (n_1_95) );
AOI211_X1 g_2_73 (.ZN (n_2_73), .A (n_2_77), .B (n_1_83), .C1 (n_1_87), .C2 (n_2_93) );
AOI211_X1 g_1_71 (.ZN (n_1_71), .A (n_1_75), .B (n_2_81), .C1 (n_2_85), .C2 (n_1_91) );
AOI211_X1 g_2_69 (.ZN (n_2_69), .A (n_2_73), .B (n_1_79), .C1 (n_1_83), .C2 (n_2_89) );
AOI211_X1 g_1_67 (.ZN (n_1_67), .A (n_1_71), .B (n_2_77), .C1 (n_2_81), .C2 (n_1_87) );
AOI211_X1 g_2_65 (.ZN (n_2_65), .A (n_2_69), .B (n_1_75), .C1 (n_1_79), .C2 (n_2_85) );
AOI211_X1 g_1_63 (.ZN (n_1_63), .A (n_1_67), .B (n_2_73), .C1 (n_2_77), .C2 (n_1_83) );
AOI211_X1 g_2_61 (.ZN (n_2_61), .A (n_2_65), .B (n_1_71), .C1 (n_1_75), .C2 (n_2_81) );
AOI211_X1 g_1_59 (.ZN (n_1_59), .A (n_1_63), .B (n_2_69), .C1 (n_2_73), .C2 (n_1_79) );
AOI211_X1 g_2_57 (.ZN (n_2_57), .A (n_2_61), .B (n_1_67), .C1 (n_1_71), .C2 (n_2_77) );
AOI211_X1 g_1_55 (.ZN (n_1_55), .A (n_1_59), .B (n_2_65), .C1 (n_2_69), .C2 (n_1_75) );
AOI211_X1 g_2_53 (.ZN (n_2_53), .A (n_2_57), .B (n_1_63), .C1 (n_1_67), .C2 (n_2_73) );
AOI211_X1 g_1_51 (.ZN (n_1_51), .A (n_1_55), .B (n_2_61), .C1 (n_2_65), .C2 (n_1_71) );
AOI211_X1 g_2_49 (.ZN (n_2_49), .A (n_2_53), .B (n_1_59), .C1 (n_1_63), .C2 (n_2_69) );
AOI211_X1 g_1_47 (.ZN (n_1_47), .A (n_1_51), .B (n_2_57), .C1 (n_2_61), .C2 (n_1_67) );
AOI211_X1 g_2_45 (.ZN (n_2_45), .A (n_2_49), .B (n_1_55), .C1 (n_1_59), .C2 (n_2_65) );
AOI211_X1 g_1_43 (.ZN (n_1_43), .A (n_1_47), .B (n_2_53), .C1 (n_2_57), .C2 (n_1_63) );
AOI211_X1 g_2_41 (.ZN (n_2_41), .A (n_2_45), .B (n_1_51), .C1 (n_1_55), .C2 (n_2_61) );
AOI211_X1 g_1_39 (.ZN (n_1_39), .A (n_1_43), .B (n_2_49), .C1 (n_2_53), .C2 (n_1_59) );
AOI211_X1 g_2_37 (.ZN (n_2_37), .A (n_2_41), .B (n_1_47), .C1 (n_1_51), .C2 (n_2_57) );
AOI211_X1 g_1_35 (.ZN (n_1_35), .A (n_1_39), .B (n_2_45), .C1 (n_2_49), .C2 (n_1_55) );
AOI211_X1 g_2_33 (.ZN (n_2_33), .A (n_2_37), .B (n_1_43), .C1 (n_1_47), .C2 (n_2_53) );
AOI211_X1 g_1_31 (.ZN (n_1_31), .A (n_1_35), .B (n_2_41), .C1 (n_2_45), .C2 (n_1_51) );
AOI211_X1 g_2_29 (.ZN (n_2_29), .A (n_2_33), .B (n_1_39), .C1 (n_1_43), .C2 (n_2_49) );
AOI211_X1 g_1_27 (.ZN (n_1_27), .A (n_1_31), .B (n_2_37), .C1 (n_2_41), .C2 (n_1_47) );
AOI211_X1 g_2_25 (.ZN (n_2_25), .A (n_2_29), .B (n_1_35), .C1 (n_1_39), .C2 (n_2_45) );
AOI211_X1 g_1_23 (.ZN (n_1_23), .A (n_1_27), .B (n_2_33), .C1 (n_2_37), .C2 (n_1_43) );
AOI211_X1 g_2_21 (.ZN (n_2_21), .A (n_2_25), .B (n_1_31), .C1 (n_1_35), .C2 (n_2_41) );
AOI211_X1 g_1_19 (.ZN (n_1_19), .A (n_1_23), .B (n_2_29), .C1 (n_2_33), .C2 (n_1_39) );
AOI211_X1 g_2_17 (.ZN (n_2_17), .A (n_2_21), .B (n_1_27), .C1 (n_1_31), .C2 (n_2_37) );
AOI211_X1 g_1_15 (.ZN (n_1_15), .A (n_1_19), .B (n_2_25), .C1 (n_2_29), .C2 (n_1_35) );
AOI211_X1 g_2_13 (.ZN (n_2_13), .A (n_2_17), .B (n_1_23), .C1 (n_1_27), .C2 (n_2_33) );
AOI211_X1 g_1_11 (.ZN (n_1_11), .A (n_1_15), .B (n_2_21), .C1 (n_2_25), .C2 (n_1_31) );
AOI211_X1 g_2_9 (.ZN (n_2_9), .A (n_2_13), .B (n_1_19), .C1 (n_1_23), .C2 (n_2_29) );
AOI211_X1 g_1_7 (.ZN (n_1_7), .A (n_1_11), .B (n_2_17), .C1 (n_2_21), .C2 (n_1_27) );
AOI211_X1 g_2_5 (.ZN (n_2_5), .A (n_2_9), .B (n_1_15), .C1 (n_1_19), .C2 (n_2_25) );
AOI211_X1 g_1_3 (.ZN (n_1_3), .A (n_1_7), .B (n_2_13), .C1 (n_2_17), .C2 (n_1_23) );
AOI211_X1 g_2_1 (.ZN (n_2_1), .A (n_2_5), .B (n_1_11), .C1 (n_1_15), .C2 (n_2_21) );
AOI211_X1 g_3_3 (.ZN (n_3_3), .A (n_1_3), .B (n_2_9), .C1 (n_2_13), .C2 (n_1_19) );
AOI211_X1 g_1_2 (.ZN (n_1_2), .A (n_2_1), .B (n_1_7), .C1 (n_1_11), .C2 (n_2_17) );
AOI211_X1 g_3_1 (.ZN (n_3_1), .A (n_3_3), .B (n_2_5), .C1 (n_2_9), .C2 (n_1_15) );
AOI211_X1 g_2_3 (.ZN (n_2_3), .A (n_1_2), .B (n_1_3), .C1 (n_1_7), .C2 (n_2_13) );
AOI211_X1 g_1_1 (.ZN (n_1_1), .A (n_3_1), .B (n_2_1), .C1 (n_2_5), .C2 (n_1_11) );
AOI211_X1 g_3_2 (.ZN (n_3_2), .A (n_2_3), .B (n_3_3), .C1 (n_1_3), .C2 (n_2_9) );
AOI211_X1 g_5_1 (.ZN (n_5_1), .A (n_1_1), .B (n_1_2), .C1 (n_2_1), .C2 (n_1_7) );
AOI211_X1 g_6_3 (.ZN (n_6_3), .A (n_3_2), .B (n_3_1), .C1 (n_3_3), .C2 (n_2_5) );
AOI211_X1 g_4_2 (.ZN (n_4_2), .A (n_5_1), .B (n_2_3), .C1 (n_1_2), .C2 (n_1_3) );
AOI211_X1 g_6_1 (.ZN (n_6_1), .A (n_6_3), .B (n_1_1), .C1 (n_3_1), .C2 (n_2_1) );
AOI211_X1 g_8_2 (.ZN (n_8_2), .A (n_4_2), .B (n_3_2), .C1 (n_2_3), .C2 (n_3_3) );
AOI211_X1 g_10_1 (.ZN (n_10_1), .A (n_6_1), .B (n_5_1), .C1 (n_1_1), .C2 (n_1_2) );
AOI211_X1 g_11_3 (.ZN (n_11_3), .A (n_8_2), .B (n_6_3), .C1 (n_3_2), .C2 (n_3_1) );
AOI211_X1 g_12_1 (.ZN (n_12_1), .A (n_10_1), .B (n_4_2), .C1 (n_5_1), .C2 (n_2_3) );
AOI211_X1 g_10_2 (.ZN (n_10_2), .A (n_11_3), .B (n_6_1), .C1 (n_6_3), .C2 (n_1_1) );
AOI211_X1 g_8_1 (.ZN (n_8_1), .A (n_12_1), .B (n_8_2), .C1 (n_4_2), .C2 (n_3_2) );
AOI211_X1 g_7_3 (.ZN (n_7_3), .A (n_10_2), .B (n_10_1), .C1 (n_6_1), .C2 (n_5_1) );
AOI211_X1 g_9_4 (.ZN (n_9_4), .A (n_8_1), .B (n_11_3), .C1 (n_8_2), .C2 (n_6_3) );
AOI211_X1 g_7_5 (.ZN (n_7_5), .A (n_7_3), .B (n_12_1), .C1 (n_10_1), .C2 (n_4_2) );
AOI211_X1 g_5_4 (.ZN (n_5_4), .A (n_9_4), .B (n_10_2), .C1 (n_11_3), .C2 (n_6_1) );
AOI211_X1 g_6_2 (.ZN (n_6_2), .A (n_7_5), .B (n_8_1), .C1 (n_12_1), .C2 (n_8_2) );
AOI211_X1 g_4_1 (.ZN (n_4_1), .A (n_5_4), .B (n_7_3), .C1 (n_10_2), .C2 (n_10_1) );
AOI211_X1 g_2_2 (.ZN (n_2_2), .A (n_6_2), .B (n_9_4), .C1 (n_8_1), .C2 (n_11_3) );
AOI211_X1 g_1_4 (.ZN (n_1_4), .A (n_4_1), .B (n_7_5), .C1 (n_7_3), .C2 (n_12_1) );
AOI211_X1 g_2_6 (.ZN (n_2_6), .A (n_2_2), .B (n_5_4), .C1 (n_9_4), .C2 (n_10_2) );
AOI211_X1 g_1_8 (.ZN (n_1_8), .A (n_1_4), .B (n_6_2), .C1 (n_7_5), .C2 (n_8_1) );
AOI211_X1 g_3_7 (.ZN (n_3_7), .A (n_2_6), .B (n_4_1), .C1 (n_5_4), .C2 (n_7_3) );
AOI211_X1 g_1_6 (.ZN (n_1_6), .A (n_1_8), .B (n_2_2), .C1 (n_6_2), .C2 (n_9_4) );
AOI211_X1 g_2_4 (.ZN (n_2_4), .A (n_3_7), .B (n_1_4), .C1 (n_4_1), .C2 (n_7_5) );
AOI211_X1 g_4_3 (.ZN (n_4_3), .A (n_1_6), .B (n_2_6), .C1 (n_2_2), .C2 (n_5_4) );
AOI211_X1 g_3_5 (.ZN (n_3_5), .A (n_2_4), .B (n_1_8), .C1 (n_1_4), .C2 (n_6_2) );
AOI211_X1 g_5_6 (.ZN (n_5_6), .A (n_4_3), .B (n_3_7), .C1 (n_2_6), .C2 (n_4_1) );
AOI211_X1 g_6_4 (.ZN (n_6_4), .A (n_3_5), .B (n_1_6), .C1 (n_1_8), .C2 (n_2_2) );
AOI211_X1 g_8_3 (.ZN (n_8_3), .A (n_5_6), .B (n_2_4), .C1 (n_3_7), .C2 (n_1_4) );
AOI211_X1 g_9_1 (.ZN (n_9_1), .A (n_6_4), .B (n_4_3), .C1 (n_1_6), .C2 (n_2_6) );
AOI211_X1 g_7_2 (.ZN (n_7_2), .A (n_8_3), .B (n_3_5), .C1 (n_2_4), .C2 (n_1_8) );
AOI211_X1 g_5_3 (.ZN (n_5_3), .A (n_9_1), .B (n_5_6), .C1 (n_4_3), .C2 (n_3_7) );
AOI211_X1 g_4_5 (.ZN (n_4_5), .A (n_7_2), .B (n_6_4), .C1 (n_3_5), .C2 (n_1_6) );
AOI211_X1 g_6_6 (.ZN (n_6_6), .A (n_5_3), .B (n_8_3), .C1 (n_5_6), .C2 (n_2_4) );
AOI211_X1 g_7_4 (.ZN (n_7_4), .A (n_4_5), .B (n_9_1), .C1 (n_6_4), .C2 (n_4_3) );
AOI211_X1 g_9_3 (.ZN (n_9_3), .A (n_6_6), .B (n_7_2), .C1 (n_8_3), .C2 (n_3_5) );
AOI211_X1 g_11_2 (.ZN (n_11_2), .A (n_7_4), .B (n_5_3), .C1 (n_9_1), .C2 (n_5_6) );
AOI211_X1 g_13_1 (.ZN (n_13_1), .A (n_9_3), .B (n_4_5), .C1 (n_7_2), .C2 (n_6_4) );
AOI211_X1 g_12_3 (.ZN (n_12_3), .A (n_11_2), .B (n_6_6), .C1 (n_5_3), .C2 (n_8_3) );
AOI211_X1 g_14_2 (.ZN (n_14_2), .A (n_13_1), .B (n_7_4), .C1 (n_4_5), .C2 (n_9_1) );
AOI211_X1 g_16_1 (.ZN (n_16_1), .A (n_12_3), .B (n_9_3), .C1 (n_6_6), .C2 (n_7_2) );
AOI211_X1 g_15_3 (.ZN (n_15_3), .A (n_14_2), .B (n_11_2), .C1 (n_7_4), .C2 (n_5_3) );
AOI211_X1 g_14_1 (.ZN (n_14_1), .A (n_16_1), .B (n_13_1), .C1 (n_9_3), .C2 (n_4_5) );
AOI211_X1 g_12_2 (.ZN (n_12_2), .A (n_15_3), .B (n_12_3), .C1 (n_11_2), .C2 (n_6_6) );
AOI211_X1 g_10_3 (.ZN (n_10_3), .A (n_14_1), .B (n_14_2), .C1 (n_13_1), .C2 (n_7_4) );
AOI211_X1 g_8_4 (.ZN (n_8_4), .A (n_12_2), .B (n_16_1), .C1 (n_12_3), .C2 (n_9_3) );
AOI211_X1 g_6_5 (.ZN (n_6_5), .A (n_10_3), .B (n_15_3), .C1 (n_14_2), .C2 (n_11_2) );
AOI211_X1 g_4_6 (.ZN (n_4_6), .A (n_8_4), .B (n_14_1), .C1 (n_16_1), .C2 (n_13_1) );
AOI211_X1 g_3_4 (.ZN (n_3_4), .A (n_6_5), .B (n_12_2), .C1 (n_15_3), .C2 (n_12_3) );
AOI211_X1 g_1_5 (.ZN (n_1_5), .A (n_4_6), .B (n_10_3), .C1 (n_14_1), .C2 (n_14_2) );
AOI211_X1 g_2_7 (.ZN (n_2_7), .A (n_3_4), .B (n_8_4), .C1 (n_12_2), .C2 (n_16_1) );
AOI211_X1 g_1_9 (.ZN (n_1_9), .A (n_1_5), .B (n_6_5), .C1 (n_10_3), .C2 (n_15_3) );
AOI211_X1 g_3_8 (.ZN (n_3_8), .A (n_2_7), .B (n_4_6), .C1 (n_8_4), .C2 (n_14_1) );
AOI211_X1 g_2_10 (.ZN (n_2_10), .A (n_1_9), .B (n_3_4), .C1 (n_6_5), .C2 (n_12_2) );
AOI211_X1 g_1_12 (.ZN (n_1_12), .A (n_3_8), .B (n_1_5), .C1 (n_4_6), .C2 (n_10_3) );
AOI211_X1 g_3_11 (.ZN (n_3_11), .A (n_2_10), .B (n_2_7), .C1 (n_3_4), .C2 (n_8_4) );
AOI211_X1 g_1_10 (.ZN (n_1_10), .A (n_1_12), .B (n_1_9), .C1 (n_1_5), .C2 (n_6_5) );
AOI211_X1 g_2_8 (.ZN (n_2_8), .A (n_3_11), .B (n_3_8), .C1 (n_2_7), .C2 (n_4_6) );
AOI211_X1 g_3_6 (.ZN (n_3_6), .A (n_1_10), .B (n_2_10), .C1 (n_1_9), .C2 (n_3_4) );
AOI211_X1 g_5_5 (.ZN (n_5_5), .A (n_2_8), .B (n_1_12), .C1 (n_3_8), .C2 (n_1_5) );
AOI211_X1 g_4_7 (.ZN (n_4_7), .A (n_3_6), .B (n_3_11), .C1 (n_2_10), .C2 (n_2_7) );
AOI211_X1 g_3_9 (.ZN (n_3_9), .A (n_5_5), .B (n_1_10), .C1 (n_1_12), .C2 (n_1_9) );
AOI211_X1 g_5_8 (.ZN (n_5_8), .A (n_4_7), .B (n_2_8), .C1 (n_3_11), .C2 (n_3_8) );
AOI211_X1 g_7_7 (.ZN (n_7_7), .A (n_3_9), .B (n_3_6), .C1 (n_1_10), .C2 (n_2_10) );
AOI211_X1 g_8_5 (.ZN (n_8_5), .A (n_5_8), .B (n_5_5), .C1 (n_2_8), .C2 (n_1_12) );
AOI211_X1 g_10_4 (.ZN (n_10_4), .A (n_7_7), .B (n_4_7), .C1 (n_3_6), .C2 (n_3_11) );
AOI211_X1 g_9_6 (.ZN (n_9_6), .A (n_8_5), .B (n_3_9), .C1 (n_5_5), .C2 (n_1_10) );
AOI211_X1 g_11_5 (.ZN (n_11_5), .A (n_10_4), .B (n_5_8), .C1 (n_4_7), .C2 (n_2_8) );
AOI211_X1 g_13_4 (.ZN (n_13_4), .A (n_9_6), .B (n_7_7), .C1 (n_3_9), .C2 (n_3_6) );
AOI211_X1 g_12_6 (.ZN (n_12_6), .A (n_11_5), .B (n_8_5), .C1 (n_5_8), .C2 (n_5_5) );
AOI211_X1 g_11_4 (.ZN (n_11_4), .A (n_13_4), .B (n_10_4), .C1 (n_7_7), .C2 (n_4_7) );
AOI211_X1 g_13_3 (.ZN (n_13_3), .A (n_12_6), .B (n_9_6), .C1 (n_8_5), .C2 (n_3_9) );
AOI211_X1 g_15_2 (.ZN (n_15_2), .A (n_11_4), .B (n_11_5), .C1 (n_10_4), .C2 (n_5_8) );
AOI211_X1 g_17_1 (.ZN (n_17_1), .A (n_13_3), .B (n_13_4), .C1 (n_9_6), .C2 (n_7_7) );
AOI211_X1 g_16_3 (.ZN (n_16_3), .A (n_15_2), .B (n_12_6), .C1 (n_11_5), .C2 (n_8_5) );
AOI211_X1 g_18_2 (.ZN (n_18_2), .A (n_17_1), .B (n_11_4), .C1 (n_13_4), .C2 (n_10_4) );
AOI211_X1 g_20_1 (.ZN (n_20_1), .A (n_16_3), .B (n_13_3), .C1 (n_12_6), .C2 (n_9_6) );
AOI211_X1 g_19_3 (.ZN (n_19_3), .A (n_18_2), .B (n_15_2), .C1 (n_11_4), .C2 (n_11_5) );
AOI211_X1 g_18_1 (.ZN (n_18_1), .A (n_20_1), .B (n_17_1), .C1 (n_13_3), .C2 (n_13_4) );
AOI211_X1 g_16_2 (.ZN (n_16_2), .A (n_19_3), .B (n_16_3), .C1 (n_15_2), .C2 (n_12_6) );
AOI211_X1 g_14_3 (.ZN (n_14_3), .A (n_18_1), .B (n_18_2), .C1 (n_17_1), .C2 (n_11_4) );
AOI211_X1 g_12_4 (.ZN (n_12_4), .A (n_16_2), .B (n_20_1), .C1 (n_16_3), .C2 (n_13_3) );
AOI211_X1 g_10_5 (.ZN (n_10_5), .A (n_14_3), .B (n_19_3), .C1 (n_18_2), .C2 (n_15_2) );
AOI211_X1 g_8_6 (.ZN (n_8_6), .A (n_12_4), .B (n_18_1), .C1 (n_20_1), .C2 (n_17_1) );
AOI211_X1 g_6_7 (.ZN (n_6_7), .A (n_10_5), .B (n_16_2), .C1 (n_19_3), .C2 (n_16_3) );
AOI211_X1 g_4_8 (.ZN (n_4_8), .A (n_8_6), .B (n_14_3), .C1 (n_18_1), .C2 (n_18_2) );
AOI211_X1 g_3_10 (.ZN (n_3_10), .A (n_6_7), .B (n_12_4), .C1 (n_16_2), .C2 (n_20_1) );
AOI211_X1 g_5_9 (.ZN (n_5_9), .A (n_4_8), .B (n_10_5), .C1 (n_14_3), .C2 (n_19_3) );
AOI211_X1 g_7_8 (.ZN (n_7_8), .A (n_3_10), .B (n_8_6), .C1 (n_12_4), .C2 (n_18_1) );
AOI211_X1 g_5_7 (.ZN (n_5_7), .A (n_5_9), .B (n_6_7), .C1 (n_10_5), .C2 (n_16_2) );
AOI211_X1 g_4_9 (.ZN (n_4_9), .A (n_7_8), .B (n_4_8), .C1 (n_8_6), .C2 (n_14_3) );
AOI211_X1 g_6_8 (.ZN (n_6_8), .A (n_5_7), .B (n_3_10), .C1 (n_6_7), .C2 (n_12_4) );
AOI211_X1 g_7_6 (.ZN (n_7_6), .A (n_4_9), .B (n_5_9), .C1 (n_4_8), .C2 (n_10_5) );
AOI211_X1 g_9_5 (.ZN (n_9_5), .A (n_6_8), .B (n_7_8), .C1 (n_3_10), .C2 (n_8_6) );
AOI211_X1 g_8_7 (.ZN (n_8_7), .A (n_7_6), .B (n_5_7), .C1 (n_5_9), .C2 (n_6_7) );
AOI211_X1 g_10_6 (.ZN (n_10_6), .A (n_9_5), .B (n_4_9), .C1 (n_7_8), .C2 (n_4_8) );
AOI211_X1 g_12_5 (.ZN (n_12_5), .A (n_8_7), .B (n_6_8), .C1 (n_5_7), .C2 (n_3_10) );
AOI211_X1 g_14_4 (.ZN (n_14_4), .A (n_10_6), .B (n_7_6), .C1 (n_4_9), .C2 (n_5_9) );
AOI211_X1 g_13_6 (.ZN (n_13_6), .A (n_12_5), .B (n_9_5), .C1 (n_6_8), .C2 (n_7_8) );
AOI211_X1 g_15_5 (.ZN (n_15_5), .A (n_14_4), .B (n_8_7), .C1 (n_7_6), .C2 (n_5_7) );
AOI211_X1 g_17_4 (.ZN (n_17_4), .A (n_13_6), .B (n_10_6), .C1 (n_9_5), .C2 (n_4_9) );
AOI211_X1 g_16_6 (.ZN (n_16_6), .A (n_15_5), .B (n_12_5), .C1 (n_8_7), .C2 (n_6_8) );
AOI211_X1 g_14_5 (.ZN (n_14_5), .A (n_17_4), .B (n_14_4), .C1 (n_10_6), .C2 (n_7_6) );
AOI211_X1 g_16_4 (.ZN (n_16_4), .A (n_16_6), .B (n_13_6), .C1 (n_12_5), .C2 (n_9_5) );
AOI211_X1 g_18_3 (.ZN (n_18_3), .A (n_14_5), .B (n_15_5), .C1 (n_14_4), .C2 (n_8_7) );
AOI211_X1 g_20_2 (.ZN (n_20_2), .A (n_16_4), .B (n_17_4), .C1 (n_13_6), .C2 (n_10_6) );
AOI211_X1 g_22_1 (.ZN (n_22_1), .A (n_18_3), .B (n_16_6), .C1 (n_15_5), .C2 (n_12_5) );
AOI211_X1 g_23_3 (.ZN (n_23_3), .A (n_20_2), .B (n_14_5), .C1 (n_17_4), .C2 (n_14_4) );
AOI211_X1 g_24_1 (.ZN (n_24_1), .A (n_22_1), .B (n_16_4), .C1 (n_16_6), .C2 (n_13_6) );
AOI211_X1 g_22_2 (.ZN (n_22_2), .A (n_23_3), .B (n_18_3), .C1 (n_14_5), .C2 (n_15_5) );
AOI211_X1 g_21_4 (.ZN (n_21_4), .A (n_24_1), .B (n_20_2), .C1 (n_16_4), .C2 (n_17_4) );
AOI211_X1 g_19_5 (.ZN (n_19_5), .A (n_22_2), .B (n_22_1), .C1 (n_18_3), .C2 (n_16_6) );
AOI211_X1 g_20_3 (.ZN (n_20_3), .A (n_21_4), .B (n_23_3), .C1 (n_20_2), .C2 (n_14_5) );
AOI211_X1 g_21_1 (.ZN (n_21_1), .A (n_19_5), .B (n_24_1), .C1 (n_22_1), .C2 (n_16_4) );
AOI211_X1 g_19_2 (.ZN (n_19_2), .A (n_20_3), .B (n_22_2), .C1 (n_23_3), .C2 (n_18_3) );
AOI211_X1 g_17_3 (.ZN (n_17_3), .A (n_21_1), .B (n_21_4), .C1 (n_24_1), .C2 (n_20_2) );
AOI211_X1 g_15_4 (.ZN (n_15_4), .A (n_19_2), .B (n_19_5), .C1 (n_22_2), .C2 (n_22_1) );
AOI211_X1 g_13_5 (.ZN (n_13_5), .A (n_17_3), .B (n_20_3), .C1 (n_21_4), .C2 (n_23_3) );
AOI211_X1 g_11_6 (.ZN (n_11_6), .A (n_15_4), .B (n_21_1), .C1 (n_19_5), .C2 (n_24_1) );
AOI211_X1 g_9_7 (.ZN (n_9_7), .A (n_13_5), .B (n_19_2), .C1 (n_20_3), .C2 (n_22_2) );
AOI211_X1 g_8_9 (.ZN (n_8_9), .A (n_11_6), .B (n_17_3), .C1 (n_21_1), .C2 (n_21_4) );
AOI211_X1 g_10_8 (.ZN (n_10_8), .A (n_9_7), .B (n_15_4), .C1 (n_19_2), .C2 (n_19_5) );
AOI211_X1 g_12_7 (.ZN (n_12_7), .A (n_8_9), .B (n_13_5), .C1 (n_17_3), .C2 (n_20_3) );
AOI211_X1 g_14_6 (.ZN (n_14_6), .A (n_10_8), .B (n_11_6), .C1 (n_15_4), .C2 (n_21_1) );
AOI211_X1 g_16_5 (.ZN (n_16_5), .A (n_12_7), .B (n_9_7), .C1 (n_13_5), .C2 (n_19_2) );
AOI211_X1 g_18_4 (.ZN (n_18_4), .A (n_14_6), .B (n_8_9), .C1 (n_11_6), .C2 (n_17_3) );
AOI211_X1 g_17_6 (.ZN (n_17_6), .A (n_16_5), .B (n_10_8), .C1 (n_9_7), .C2 (n_15_4) );
AOI211_X1 g_15_7 (.ZN (n_15_7), .A (n_18_4), .B (n_12_7), .C1 (n_8_9), .C2 (n_13_5) );
AOI211_X1 g_13_8 (.ZN (n_13_8), .A (n_17_6), .B (n_14_6), .C1 (n_10_8), .C2 (n_11_6) );
AOI211_X1 g_11_7 (.ZN (n_11_7), .A (n_15_7), .B (n_16_5), .C1 (n_12_7), .C2 (n_9_7) );
AOI211_X1 g_9_8 (.ZN (n_9_8), .A (n_13_8), .B (n_18_4), .C1 (n_14_6), .C2 (n_8_9) );
AOI211_X1 g_7_9 (.ZN (n_7_9), .A (n_11_7), .B (n_17_6), .C1 (n_16_5), .C2 (n_10_8) );
AOI211_X1 g_5_10 (.ZN (n_5_10), .A (n_9_8), .B (n_15_7), .C1 (n_18_4), .C2 (n_12_7) );
AOI211_X1 g_4_12 (.ZN (n_4_12), .A (n_7_9), .B (n_13_8), .C1 (n_17_6), .C2 (n_14_6) );
AOI211_X1 g_2_11 (.ZN (n_2_11), .A (n_5_10), .B (n_11_7), .C1 (n_15_7), .C2 (n_16_5) );
AOI211_X1 g_1_13 (.ZN (n_1_13), .A (n_4_12), .B (n_9_8), .C1 (n_13_8), .C2 (n_18_4) );
AOI211_X1 g_3_12 (.ZN (n_3_12), .A (n_2_11), .B (n_7_9), .C1 (n_11_7), .C2 (n_17_6) );
AOI211_X1 g_4_10 (.ZN (n_4_10), .A (n_1_13), .B (n_5_10), .C1 (n_9_8), .C2 (n_15_7) );
AOI211_X1 g_6_9 (.ZN (n_6_9), .A (n_3_12), .B (n_4_12), .C1 (n_7_9), .C2 (n_13_8) );
AOI211_X1 g_8_8 (.ZN (n_8_8), .A (n_4_10), .B (n_2_11), .C1 (n_5_10), .C2 (n_11_7) );
AOI211_X1 g_10_7 (.ZN (n_10_7), .A (n_6_9), .B (n_1_13), .C1 (n_4_12), .C2 (n_9_8) );
AOI211_X1 g_11_9 (.ZN (n_11_9), .A (n_8_8), .B (n_3_12), .C1 (n_2_11), .C2 (n_7_9) );
AOI211_X1 g_9_10 (.ZN (n_9_10), .A (n_10_7), .B (n_4_10), .C1 (n_1_13), .C2 (n_5_10) );
AOI211_X1 g_7_11 (.ZN (n_7_11), .A (n_11_9), .B (n_6_9), .C1 (n_3_12), .C2 (n_4_12) );
AOI211_X1 g_5_12 (.ZN (n_5_12), .A (n_9_10), .B (n_8_8), .C1 (n_4_10), .C2 (n_2_11) );
AOI211_X1 g_6_10 (.ZN (n_6_10), .A (n_7_11), .B (n_10_7), .C1 (n_6_9), .C2 (n_1_13) );
AOI211_X1 g_4_11 (.ZN (n_4_11), .A (n_5_12), .B (n_11_9), .C1 (n_8_8), .C2 (n_3_12) );
AOI211_X1 g_2_12 (.ZN (n_2_12), .A (n_6_10), .B (n_9_10), .C1 (n_10_7), .C2 (n_4_10) );
AOI211_X1 g_1_14 (.ZN (n_1_14), .A (n_4_11), .B (n_7_11), .C1 (n_11_9), .C2 (n_6_9) );
AOI211_X1 g_3_13 (.ZN (n_3_13), .A (n_2_12), .B (n_5_12), .C1 (n_9_10), .C2 (n_8_8) );
AOI211_X1 g_2_15 (.ZN (n_2_15), .A (n_1_14), .B (n_6_10), .C1 (n_7_11), .C2 (n_10_7) );
AOI211_X1 g_1_17 (.ZN (n_1_17), .A (n_3_13), .B (n_4_11), .C1 (n_5_12), .C2 (n_11_9) );
AOI211_X1 g_2_19 (.ZN (n_2_19), .A (n_2_15), .B (n_2_12), .C1 (n_6_10), .C2 (n_9_10) );
AOI211_X1 g_1_21 (.ZN (n_1_21), .A (n_1_17), .B (n_1_14), .C1 (n_4_11), .C2 (n_7_11) );
AOI211_X1 g_2_23 (.ZN (n_2_23), .A (n_2_19), .B (n_3_13), .C1 (n_2_12), .C2 (n_5_12) );
AOI211_X1 g_1_25 (.ZN (n_1_25), .A (n_1_21), .B (n_2_15), .C1 (n_1_14), .C2 (n_6_10) );
AOI211_X1 g_2_27 (.ZN (n_2_27), .A (n_2_23), .B (n_1_17), .C1 (n_3_13), .C2 (n_4_11) );
AOI211_X1 g_1_29 (.ZN (n_1_29), .A (n_1_25), .B (n_2_19), .C1 (n_2_15), .C2 (n_2_12) );
AOI211_X1 g_2_31 (.ZN (n_2_31), .A (n_2_27), .B (n_1_21), .C1 (n_1_17), .C2 (n_1_14) );
AOI211_X1 g_1_33 (.ZN (n_1_33), .A (n_1_29), .B (n_2_23), .C1 (n_2_19), .C2 (n_3_13) );
AOI211_X1 g_2_35 (.ZN (n_2_35), .A (n_2_31), .B (n_1_25), .C1 (n_1_21), .C2 (n_2_15) );
AOI211_X1 g_1_37 (.ZN (n_1_37), .A (n_1_33), .B (n_2_27), .C1 (n_2_23), .C2 (n_1_17) );
AOI211_X1 g_2_39 (.ZN (n_2_39), .A (n_2_35), .B (n_1_29), .C1 (n_1_25), .C2 (n_2_19) );
AOI211_X1 g_1_41 (.ZN (n_1_41), .A (n_1_37), .B (n_2_31), .C1 (n_2_27), .C2 (n_1_21) );
AOI211_X1 g_2_43 (.ZN (n_2_43), .A (n_2_39), .B (n_1_33), .C1 (n_1_29), .C2 (n_2_23) );
AOI211_X1 g_1_45 (.ZN (n_1_45), .A (n_1_41), .B (n_2_35), .C1 (n_2_31), .C2 (n_1_25) );
AOI211_X1 g_2_47 (.ZN (n_2_47), .A (n_2_43), .B (n_1_37), .C1 (n_1_33), .C2 (n_2_27) );
AOI211_X1 g_1_49 (.ZN (n_1_49), .A (n_1_45), .B (n_2_39), .C1 (n_2_35), .C2 (n_1_29) );
AOI211_X1 g_2_51 (.ZN (n_2_51), .A (n_2_47), .B (n_1_41), .C1 (n_1_37), .C2 (n_2_31) );
AOI211_X1 g_1_53 (.ZN (n_1_53), .A (n_1_49), .B (n_2_43), .C1 (n_2_39), .C2 (n_1_33) );
AOI211_X1 g_2_55 (.ZN (n_2_55), .A (n_2_51), .B (n_1_45), .C1 (n_1_41), .C2 (n_2_35) );
AOI211_X1 g_1_57 (.ZN (n_1_57), .A (n_1_53), .B (n_2_47), .C1 (n_2_43), .C2 (n_1_37) );
AOI211_X1 g_2_59 (.ZN (n_2_59), .A (n_2_55), .B (n_1_49), .C1 (n_1_45), .C2 (n_2_39) );
AOI211_X1 g_1_61 (.ZN (n_1_61), .A (n_1_57), .B (n_2_51), .C1 (n_2_47), .C2 (n_1_41) );
AOI211_X1 g_2_63 (.ZN (n_2_63), .A (n_2_59), .B (n_1_53), .C1 (n_1_49), .C2 (n_2_43) );
AOI211_X1 g_1_65 (.ZN (n_1_65), .A (n_1_61), .B (n_2_55), .C1 (n_2_51), .C2 (n_1_45) );
AOI211_X1 g_2_67 (.ZN (n_2_67), .A (n_2_63), .B (n_1_57), .C1 (n_1_53), .C2 (n_2_47) );
AOI211_X1 g_1_69 (.ZN (n_1_69), .A (n_1_65), .B (n_2_59), .C1 (n_2_55), .C2 (n_1_49) );
AOI211_X1 g_2_71 (.ZN (n_2_71), .A (n_2_67), .B (n_1_61), .C1 (n_1_57), .C2 (n_2_51) );
AOI211_X1 g_1_73 (.ZN (n_1_73), .A (n_1_69), .B (n_2_63), .C1 (n_2_59), .C2 (n_1_53) );
AOI211_X1 g_2_75 (.ZN (n_2_75), .A (n_2_71), .B (n_1_65), .C1 (n_1_61), .C2 (n_2_55) );
AOI211_X1 g_1_77 (.ZN (n_1_77), .A (n_1_73), .B (n_2_67), .C1 (n_2_63), .C2 (n_1_57) );
AOI211_X1 g_2_79 (.ZN (n_2_79), .A (n_2_75), .B (n_1_69), .C1 (n_1_65), .C2 (n_2_59) );
AOI211_X1 g_1_81 (.ZN (n_1_81), .A (n_1_77), .B (n_2_71), .C1 (n_2_67), .C2 (n_1_61) );
AOI211_X1 g_2_83 (.ZN (n_2_83), .A (n_2_79), .B (n_1_73), .C1 (n_1_69), .C2 (n_2_63) );
AOI211_X1 g_1_85 (.ZN (n_1_85), .A (n_1_81), .B (n_2_75), .C1 (n_2_71), .C2 (n_1_65) );
AOI211_X1 g_2_87 (.ZN (n_2_87), .A (n_2_83), .B (n_1_77), .C1 (n_1_73), .C2 (n_2_67) );
AOI211_X1 g_1_89 (.ZN (n_1_89), .A (n_1_85), .B (n_2_79), .C1 (n_2_75), .C2 (n_1_69) );
AOI211_X1 g_2_91 (.ZN (n_2_91), .A (n_2_87), .B (n_1_81), .C1 (n_1_77), .C2 (n_2_71) );
AOI211_X1 g_1_93 (.ZN (n_1_93), .A (n_1_89), .B (n_2_83), .C1 (n_2_79), .C2 (n_1_73) );
AOI211_X1 g_2_95 (.ZN (n_2_95), .A (n_2_91), .B (n_1_85), .C1 (n_1_81), .C2 (n_2_75) );
AOI211_X1 g_1_97 (.ZN (n_1_97), .A (n_1_93), .B (n_2_87), .C1 (n_2_83), .C2 (n_1_77) );
AOI211_X1 g_2_99 (.ZN (n_2_99), .A (n_2_95), .B (n_1_89), .C1 (n_1_85), .C2 (n_2_79) );
AOI211_X1 g_4_100 (.ZN (n_4_100), .A (n_1_97), .B (n_2_91), .C1 (n_2_87), .C2 (n_1_81) );
AOI211_X1 g_3_98 (.ZN (n_3_98), .A (n_2_99), .B (n_1_93), .C1 (n_1_89), .C2 (n_2_83) );
AOI211_X1 g_2_100 (.ZN (n_2_100), .A (n_4_100), .B (n_2_95), .C1 (n_2_91), .C2 (n_1_85) );
AOI211_X1 g_1_98 (.ZN (n_1_98), .A (n_3_98), .B (n_1_97), .C1 (n_1_93), .C2 (n_2_87) );
AOI211_X1 g_2_96 (.ZN (n_2_96), .A (n_2_100), .B (n_2_99), .C1 (n_2_95), .C2 (n_1_89) );
AOI211_X1 g_1_94 (.ZN (n_1_94), .A (n_1_98), .B (n_4_100), .C1 (n_1_97), .C2 (n_2_91) );
AOI211_X1 g_3_93 (.ZN (n_3_93), .A (n_2_96), .B (n_3_98), .C1 (n_2_99), .C2 (n_1_93) );
AOI211_X1 g_1_92 (.ZN (n_1_92), .A (n_1_94), .B (n_2_100), .C1 (n_4_100), .C2 (n_2_95) );
AOI211_X1 g_3_91 (.ZN (n_3_91), .A (n_3_93), .B (n_1_98), .C1 (n_3_98), .C2 (n_1_97) );
AOI211_X1 g_1_90 (.ZN (n_1_90), .A (n_1_92), .B (n_2_96), .C1 (n_2_100), .C2 (n_2_99) );
AOI211_X1 g_2_92 (.ZN (n_2_92), .A (n_3_91), .B (n_1_94), .C1 (n_1_98), .C2 (n_4_100) );
AOI211_X1 g_3_94 (.ZN (n_3_94), .A (n_1_90), .B (n_3_93), .C1 (n_2_96), .C2 (n_3_98) );
AOI211_X1 g_4_96 (.ZN (n_4_96), .A (n_2_92), .B (n_1_92), .C1 (n_1_94), .C2 (n_2_100) );
AOI211_X1 g_5_94 (.ZN (n_5_94), .A (n_3_94), .B (n_3_91), .C1 (n_3_93), .C2 (n_1_98) );
AOI211_X1 g_4_92 (.ZN (n_4_92), .A (n_4_96), .B (n_1_90), .C1 (n_1_92), .C2 (n_2_96) );
AOI211_X1 g_3_90 (.ZN (n_3_90), .A (n_5_94), .B (n_2_92), .C1 (n_3_91), .C2 (n_1_94) );
AOI211_X1 g_2_88 (.ZN (n_2_88), .A (n_4_92), .B (n_3_94), .C1 (n_1_90), .C2 (n_3_93) );
AOI211_X1 g_1_86 (.ZN (n_1_86), .A (n_3_90), .B (n_4_96), .C1 (n_2_92), .C2 (n_1_92) );
AOI211_X1 g_3_85 (.ZN (n_3_85), .A (n_2_88), .B (n_5_94), .C1 (n_3_94), .C2 (n_3_91) );
AOI211_X1 g_1_84 (.ZN (n_1_84), .A (n_1_86), .B (n_4_92), .C1 (n_4_96), .C2 (n_1_90) );
AOI211_X1 g_3_83 (.ZN (n_3_83), .A (n_3_85), .B (n_3_90), .C1 (n_5_94), .C2 (n_2_92) );
AOI211_X1 g_1_82 (.ZN (n_1_82), .A (n_1_84), .B (n_2_88), .C1 (n_4_92), .C2 (n_3_94) );
AOI211_X1 g_2_84 (.ZN (n_2_84), .A (n_3_83), .B (n_1_86), .C1 (n_3_90), .C2 (n_4_96) );
AOI211_X1 g_3_86 (.ZN (n_3_86), .A (n_1_82), .B (n_3_85), .C1 (n_2_88), .C2 (n_5_94) );
AOI211_X1 g_4_88 (.ZN (n_4_88), .A (n_2_84), .B (n_1_84), .C1 (n_1_86), .C2 (n_4_92) );
AOI211_X1 g_5_90 (.ZN (n_5_90), .A (n_3_86), .B (n_3_83), .C1 (n_3_85), .C2 (n_3_90) );
AOI211_X1 g_3_89 (.ZN (n_3_89), .A (n_4_88), .B (n_1_82), .C1 (n_1_84), .C2 (n_2_88) );
AOI211_X1 g_1_88 (.ZN (n_1_88), .A (n_5_90), .B (n_2_84), .C1 (n_3_83), .C2 (n_1_86) );
AOI211_X1 g_3_87 (.ZN (n_3_87), .A (n_3_89), .B (n_3_86), .C1 (n_1_82), .C2 (n_3_85) );
AOI211_X1 g_5_86 (.ZN (n_5_86), .A (n_1_88), .B (n_4_88), .C1 (n_2_84), .C2 (n_1_84) );
AOI211_X1 g_4_84 (.ZN (n_4_84), .A (n_3_87), .B (n_5_90), .C1 (n_3_86), .C2 (n_3_83) );
AOI211_X1 g_3_82 (.ZN (n_3_82), .A (n_5_86), .B (n_3_89), .C1 (n_4_88), .C2 (n_1_82) );
AOI211_X1 g_2_80 (.ZN (n_2_80), .A (n_4_84), .B (n_1_88), .C1 (n_5_90), .C2 (n_2_84) );
AOI211_X1 g_1_78 (.ZN (n_1_78), .A (n_3_82), .B (n_3_87), .C1 (n_3_89), .C2 (n_3_86) );
AOI211_X1 g_3_77 (.ZN (n_3_77), .A (n_2_80), .B (n_5_86), .C1 (n_1_88), .C2 (n_4_88) );
AOI211_X1 g_1_76 (.ZN (n_1_76), .A (n_1_78), .B (n_4_84), .C1 (n_3_87), .C2 (n_5_90) );
AOI211_X1 g_3_75 (.ZN (n_3_75), .A (n_3_77), .B (n_3_82), .C1 (n_5_86), .C2 (n_3_89) );
AOI211_X1 g_1_74 (.ZN (n_1_74), .A (n_1_76), .B (n_2_80), .C1 (n_4_84), .C2 (n_1_88) );
AOI211_X1 g_2_76 (.ZN (n_2_76), .A (n_3_75), .B (n_1_78), .C1 (n_3_82), .C2 (n_3_87) );
AOI211_X1 g_3_78 (.ZN (n_3_78), .A (n_1_74), .B (n_3_77), .C1 (n_2_80), .C2 (n_5_86) );
AOI211_X1 g_4_80 (.ZN (n_4_80), .A (n_2_76), .B (n_1_76), .C1 (n_1_78), .C2 (n_4_84) );
AOI211_X1 g_5_82 (.ZN (n_5_82), .A (n_3_78), .B (n_3_75), .C1 (n_3_77), .C2 (n_3_82) );
AOI211_X1 g_3_81 (.ZN (n_3_81), .A (n_4_80), .B (n_1_74), .C1 (n_1_76), .C2 (n_2_80) );
AOI211_X1 g_1_80 (.ZN (n_1_80), .A (n_5_82), .B (n_2_76), .C1 (n_3_75), .C2 (n_1_78) );
AOI211_X1 g_3_79 (.ZN (n_3_79), .A (n_3_81), .B (n_3_78), .C1 (n_1_74), .C2 (n_3_77) );
AOI211_X1 g_5_78 (.ZN (n_5_78), .A (n_1_80), .B (n_4_80), .C1 (n_2_76), .C2 (n_1_76) );
AOI211_X1 g_4_76 (.ZN (n_4_76), .A (n_3_79), .B (n_5_82), .C1 (n_3_78), .C2 (n_3_75) );
AOI211_X1 g_3_74 (.ZN (n_3_74), .A (n_5_78), .B (n_3_81), .C1 (n_4_80), .C2 (n_1_74) );
AOI211_X1 g_2_72 (.ZN (n_2_72), .A (n_4_76), .B (n_1_80), .C1 (n_5_82), .C2 (n_2_76) );
AOI211_X1 g_1_70 (.ZN (n_1_70), .A (n_3_74), .B (n_3_79), .C1 (n_3_81), .C2 (n_3_78) );
AOI211_X1 g_3_69 (.ZN (n_3_69), .A (n_2_72), .B (n_5_78), .C1 (n_1_80), .C2 (n_4_80) );
AOI211_X1 g_1_68 (.ZN (n_1_68), .A (n_1_70), .B (n_4_76), .C1 (n_3_79), .C2 (n_5_82) );
AOI211_X1 g_3_67 (.ZN (n_3_67), .A (n_3_69), .B (n_3_74), .C1 (n_5_78), .C2 (n_3_81) );
AOI211_X1 g_1_66 (.ZN (n_1_66), .A (n_1_68), .B (n_2_72), .C1 (n_4_76), .C2 (n_1_80) );
AOI211_X1 g_2_68 (.ZN (n_2_68), .A (n_3_67), .B (n_1_70), .C1 (n_3_74), .C2 (n_3_79) );
AOI211_X1 g_3_70 (.ZN (n_3_70), .A (n_1_66), .B (n_3_69), .C1 (n_2_72), .C2 (n_5_78) );
AOI211_X1 g_4_72 (.ZN (n_4_72), .A (n_2_68), .B (n_1_68), .C1 (n_1_70), .C2 (n_4_76) );
AOI211_X1 g_5_74 (.ZN (n_5_74), .A (n_3_70), .B (n_3_67), .C1 (n_3_69), .C2 (n_3_74) );
AOI211_X1 g_3_73 (.ZN (n_3_73), .A (n_4_72), .B (n_1_66), .C1 (n_1_68), .C2 (n_2_72) );
AOI211_X1 g_1_72 (.ZN (n_1_72), .A (n_5_74), .B (n_2_68), .C1 (n_3_67), .C2 (n_1_70) );
AOI211_X1 g_3_71 (.ZN (n_3_71), .A (n_3_73), .B (n_3_70), .C1 (n_1_66), .C2 (n_3_69) );
AOI211_X1 g_5_70 (.ZN (n_5_70), .A (n_1_72), .B (n_4_72), .C1 (n_2_68), .C2 (n_1_68) );
AOI211_X1 g_4_68 (.ZN (n_4_68), .A (n_3_71), .B (n_5_74), .C1 (n_3_70), .C2 (n_3_67) );
AOI211_X1 g_3_66 (.ZN (n_3_66), .A (n_5_70), .B (n_3_73), .C1 (n_4_72), .C2 (n_1_66) );
AOI211_X1 g_2_64 (.ZN (n_2_64), .A (n_4_68), .B (n_1_72), .C1 (n_5_74), .C2 (n_2_68) );
AOI211_X1 g_1_62 (.ZN (n_1_62), .A (n_3_66), .B (n_3_71), .C1 (n_3_73), .C2 (n_3_70) );
AOI211_X1 g_3_61 (.ZN (n_3_61), .A (n_2_64), .B (n_5_70), .C1 (n_1_72), .C2 (n_4_72) );
AOI211_X1 g_1_60 (.ZN (n_1_60), .A (n_1_62), .B (n_4_68), .C1 (n_3_71), .C2 (n_5_74) );
AOI211_X1 g_3_59 (.ZN (n_3_59), .A (n_3_61), .B (n_3_66), .C1 (n_5_70), .C2 (n_3_73) );
AOI211_X1 g_1_58 (.ZN (n_1_58), .A (n_1_60), .B (n_2_64), .C1 (n_4_68), .C2 (n_1_72) );
AOI211_X1 g_2_60 (.ZN (n_2_60), .A (n_3_59), .B (n_1_62), .C1 (n_3_66), .C2 (n_3_71) );
AOI211_X1 g_3_62 (.ZN (n_3_62), .A (n_1_58), .B (n_3_61), .C1 (n_2_64), .C2 (n_5_70) );
AOI211_X1 g_4_64 (.ZN (n_4_64), .A (n_2_60), .B (n_1_60), .C1 (n_1_62), .C2 (n_4_68) );
AOI211_X1 g_5_66 (.ZN (n_5_66), .A (n_3_62), .B (n_3_59), .C1 (n_3_61), .C2 (n_3_66) );
AOI211_X1 g_3_65 (.ZN (n_3_65), .A (n_4_64), .B (n_1_58), .C1 (n_1_60), .C2 (n_2_64) );
AOI211_X1 g_1_64 (.ZN (n_1_64), .A (n_5_66), .B (n_2_60), .C1 (n_3_59), .C2 (n_1_62) );
AOI211_X1 g_3_63 (.ZN (n_3_63), .A (n_3_65), .B (n_3_62), .C1 (n_1_58), .C2 (n_3_61) );
AOI211_X1 g_5_62 (.ZN (n_5_62), .A (n_1_64), .B (n_4_64), .C1 (n_2_60), .C2 (n_1_60) );
AOI211_X1 g_4_60 (.ZN (n_4_60), .A (n_3_63), .B (n_5_66), .C1 (n_3_62), .C2 (n_3_59) );
AOI211_X1 g_3_58 (.ZN (n_3_58), .A (n_5_62), .B (n_3_65), .C1 (n_4_64), .C2 (n_1_58) );
AOI211_X1 g_2_56 (.ZN (n_2_56), .A (n_4_60), .B (n_1_64), .C1 (n_5_66), .C2 (n_2_60) );
AOI211_X1 g_1_54 (.ZN (n_1_54), .A (n_3_58), .B (n_3_63), .C1 (n_3_65), .C2 (n_3_62) );
AOI211_X1 g_3_53 (.ZN (n_3_53), .A (n_2_56), .B (n_5_62), .C1 (n_1_64), .C2 (n_4_64) );
AOI211_X1 g_1_52 (.ZN (n_1_52), .A (n_1_54), .B (n_4_60), .C1 (n_3_63), .C2 (n_5_66) );
AOI211_X1 g_3_51 (.ZN (n_3_51), .A (n_3_53), .B (n_3_58), .C1 (n_5_62), .C2 (n_3_65) );
AOI211_X1 g_1_50 (.ZN (n_1_50), .A (n_1_52), .B (n_2_56), .C1 (n_4_60), .C2 (n_1_64) );
AOI211_X1 g_2_52 (.ZN (n_2_52), .A (n_3_51), .B (n_1_54), .C1 (n_3_58), .C2 (n_3_63) );
AOI211_X1 g_3_54 (.ZN (n_3_54), .A (n_1_50), .B (n_3_53), .C1 (n_2_56), .C2 (n_5_62) );
AOI211_X1 g_4_56 (.ZN (n_4_56), .A (n_2_52), .B (n_1_52), .C1 (n_1_54), .C2 (n_4_60) );
AOI211_X1 g_5_58 (.ZN (n_5_58), .A (n_3_54), .B (n_3_51), .C1 (n_3_53), .C2 (n_3_58) );
AOI211_X1 g_3_57 (.ZN (n_3_57), .A (n_4_56), .B (n_1_50), .C1 (n_1_52), .C2 (n_2_56) );
AOI211_X1 g_1_56 (.ZN (n_1_56), .A (n_5_58), .B (n_2_52), .C1 (n_3_51), .C2 (n_1_54) );
AOI211_X1 g_3_55 (.ZN (n_3_55), .A (n_3_57), .B (n_3_54), .C1 (n_1_50), .C2 (n_3_53) );
AOI211_X1 g_5_54 (.ZN (n_5_54), .A (n_1_56), .B (n_4_56), .C1 (n_2_52), .C2 (n_1_52) );
AOI211_X1 g_4_52 (.ZN (n_4_52), .A (n_3_55), .B (n_5_58), .C1 (n_3_54), .C2 (n_3_51) );
AOI211_X1 g_3_50 (.ZN (n_3_50), .A (n_5_54), .B (n_3_57), .C1 (n_4_56), .C2 (n_1_50) );
AOI211_X1 g_2_48 (.ZN (n_2_48), .A (n_4_52), .B (n_1_56), .C1 (n_5_58), .C2 (n_2_52) );
AOI211_X1 g_1_46 (.ZN (n_1_46), .A (n_3_50), .B (n_3_55), .C1 (n_3_57), .C2 (n_3_54) );
AOI211_X1 g_3_45 (.ZN (n_3_45), .A (n_2_48), .B (n_5_54), .C1 (n_1_56), .C2 (n_4_56) );
AOI211_X1 g_1_44 (.ZN (n_1_44), .A (n_1_46), .B (n_4_52), .C1 (n_3_55), .C2 (n_5_58) );
AOI211_X1 g_3_43 (.ZN (n_3_43), .A (n_3_45), .B (n_3_50), .C1 (n_5_54), .C2 (n_3_57) );
AOI211_X1 g_1_42 (.ZN (n_1_42), .A (n_1_44), .B (n_2_48), .C1 (n_4_52), .C2 (n_1_56) );
AOI211_X1 g_2_44 (.ZN (n_2_44), .A (n_3_43), .B (n_1_46), .C1 (n_3_50), .C2 (n_3_55) );
AOI211_X1 g_3_46 (.ZN (n_3_46), .A (n_1_42), .B (n_3_45), .C1 (n_2_48), .C2 (n_5_54) );
AOI211_X1 g_4_48 (.ZN (n_4_48), .A (n_2_44), .B (n_1_44), .C1 (n_1_46), .C2 (n_4_52) );
AOI211_X1 g_5_50 (.ZN (n_5_50), .A (n_3_46), .B (n_3_43), .C1 (n_3_45), .C2 (n_3_50) );
AOI211_X1 g_3_49 (.ZN (n_3_49), .A (n_4_48), .B (n_1_42), .C1 (n_1_44), .C2 (n_2_48) );
AOI211_X1 g_1_48 (.ZN (n_1_48), .A (n_5_50), .B (n_2_44), .C1 (n_3_43), .C2 (n_1_46) );
AOI211_X1 g_3_47 (.ZN (n_3_47), .A (n_3_49), .B (n_3_46), .C1 (n_1_42), .C2 (n_3_45) );
AOI211_X1 g_5_46 (.ZN (n_5_46), .A (n_1_48), .B (n_4_48), .C1 (n_2_44), .C2 (n_1_44) );
AOI211_X1 g_4_44 (.ZN (n_4_44), .A (n_3_47), .B (n_5_50), .C1 (n_3_46), .C2 (n_3_43) );
AOI211_X1 g_3_42 (.ZN (n_3_42), .A (n_5_46), .B (n_3_49), .C1 (n_4_48), .C2 (n_1_42) );
AOI211_X1 g_2_40 (.ZN (n_2_40), .A (n_4_44), .B (n_1_48), .C1 (n_5_50), .C2 (n_2_44) );
AOI211_X1 g_1_38 (.ZN (n_1_38), .A (n_3_42), .B (n_3_47), .C1 (n_3_49), .C2 (n_3_46) );
AOI211_X1 g_3_37 (.ZN (n_3_37), .A (n_2_40), .B (n_5_46), .C1 (n_1_48), .C2 (n_4_48) );
AOI211_X1 g_1_36 (.ZN (n_1_36), .A (n_1_38), .B (n_4_44), .C1 (n_3_47), .C2 (n_5_50) );
AOI211_X1 g_3_35 (.ZN (n_3_35), .A (n_3_37), .B (n_3_42), .C1 (n_5_46), .C2 (n_3_49) );
AOI211_X1 g_1_34 (.ZN (n_1_34), .A (n_1_36), .B (n_2_40), .C1 (n_4_44), .C2 (n_1_48) );
AOI211_X1 g_2_36 (.ZN (n_2_36), .A (n_3_35), .B (n_1_38), .C1 (n_3_42), .C2 (n_3_47) );
AOI211_X1 g_3_38 (.ZN (n_3_38), .A (n_1_34), .B (n_3_37), .C1 (n_2_40), .C2 (n_5_46) );
AOI211_X1 g_4_40 (.ZN (n_4_40), .A (n_2_36), .B (n_1_36), .C1 (n_1_38), .C2 (n_4_44) );
AOI211_X1 g_5_42 (.ZN (n_5_42), .A (n_3_38), .B (n_3_35), .C1 (n_3_37), .C2 (n_3_42) );
AOI211_X1 g_3_41 (.ZN (n_3_41), .A (n_4_40), .B (n_1_34), .C1 (n_1_36), .C2 (n_2_40) );
AOI211_X1 g_1_40 (.ZN (n_1_40), .A (n_5_42), .B (n_2_36), .C1 (n_3_35), .C2 (n_1_38) );
AOI211_X1 g_3_39 (.ZN (n_3_39), .A (n_3_41), .B (n_3_38), .C1 (n_1_34), .C2 (n_3_37) );
AOI211_X1 g_5_38 (.ZN (n_5_38), .A (n_1_40), .B (n_4_40), .C1 (n_2_36), .C2 (n_1_36) );
AOI211_X1 g_4_36 (.ZN (n_4_36), .A (n_3_39), .B (n_5_42), .C1 (n_3_38), .C2 (n_3_35) );
AOI211_X1 g_3_34 (.ZN (n_3_34), .A (n_5_38), .B (n_3_41), .C1 (n_4_40), .C2 (n_1_34) );
AOI211_X1 g_2_32 (.ZN (n_2_32), .A (n_4_36), .B (n_1_40), .C1 (n_5_42), .C2 (n_2_36) );
AOI211_X1 g_1_30 (.ZN (n_1_30), .A (n_3_34), .B (n_3_39), .C1 (n_3_41), .C2 (n_3_38) );
AOI211_X1 g_3_29 (.ZN (n_3_29), .A (n_2_32), .B (n_5_38), .C1 (n_1_40), .C2 (n_4_40) );
AOI211_X1 g_1_28 (.ZN (n_1_28), .A (n_1_30), .B (n_4_36), .C1 (n_3_39), .C2 (n_5_42) );
AOI211_X1 g_3_27 (.ZN (n_3_27), .A (n_3_29), .B (n_3_34), .C1 (n_5_38), .C2 (n_3_41) );
AOI211_X1 g_1_26 (.ZN (n_1_26), .A (n_1_28), .B (n_2_32), .C1 (n_4_36), .C2 (n_1_40) );
AOI211_X1 g_2_28 (.ZN (n_2_28), .A (n_3_27), .B (n_1_30), .C1 (n_3_34), .C2 (n_3_39) );
AOI211_X1 g_3_30 (.ZN (n_3_30), .A (n_1_26), .B (n_3_29), .C1 (n_2_32), .C2 (n_5_38) );
AOI211_X1 g_4_32 (.ZN (n_4_32), .A (n_2_28), .B (n_1_28), .C1 (n_1_30), .C2 (n_4_36) );
AOI211_X1 g_5_34 (.ZN (n_5_34), .A (n_3_30), .B (n_3_27), .C1 (n_3_29), .C2 (n_3_34) );
AOI211_X1 g_3_33 (.ZN (n_3_33), .A (n_4_32), .B (n_1_26), .C1 (n_1_28), .C2 (n_2_32) );
AOI211_X1 g_1_32 (.ZN (n_1_32), .A (n_5_34), .B (n_2_28), .C1 (n_3_27), .C2 (n_1_30) );
AOI211_X1 g_3_31 (.ZN (n_3_31), .A (n_3_33), .B (n_3_30), .C1 (n_1_26), .C2 (n_3_29) );
AOI211_X1 g_5_30 (.ZN (n_5_30), .A (n_1_32), .B (n_4_32), .C1 (n_2_28), .C2 (n_1_28) );
AOI211_X1 g_4_28 (.ZN (n_4_28), .A (n_3_31), .B (n_5_34), .C1 (n_3_30), .C2 (n_3_27) );
AOI211_X1 g_3_26 (.ZN (n_3_26), .A (n_5_30), .B (n_3_33), .C1 (n_4_32), .C2 (n_1_26) );
AOI211_X1 g_2_24 (.ZN (n_2_24), .A (n_4_28), .B (n_1_32), .C1 (n_5_34), .C2 (n_2_28) );
AOI211_X1 g_1_22 (.ZN (n_1_22), .A (n_3_26), .B (n_3_31), .C1 (n_3_33), .C2 (n_3_30) );
AOI211_X1 g_3_21 (.ZN (n_3_21), .A (n_2_24), .B (n_5_30), .C1 (n_1_32), .C2 (n_4_32) );
AOI211_X1 g_1_20 (.ZN (n_1_20), .A (n_1_22), .B (n_4_28), .C1 (n_3_31), .C2 (n_5_34) );
AOI211_X1 g_3_19 (.ZN (n_3_19), .A (n_3_21), .B (n_3_26), .C1 (n_5_30), .C2 (n_3_33) );
AOI211_X1 g_1_18 (.ZN (n_1_18), .A (n_1_20), .B (n_2_24), .C1 (n_4_28), .C2 (n_1_32) );
AOI211_X1 g_2_16 (.ZN (n_2_16), .A (n_3_19), .B (n_1_22), .C1 (n_3_26), .C2 (n_3_31) );
AOI211_X1 g_3_14 (.ZN (n_3_14), .A (n_1_18), .B (n_3_21), .C1 (n_2_24), .C2 (n_5_30) );
AOI211_X1 g_5_13 (.ZN (n_5_13), .A (n_2_16), .B (n_1_20), .C1 (n_1_22), .C2 (n_4_28) );
AOI211_X1 g_6_11 (.ZN (n_6_11), .A (n_3_14), .B (n_3_19), .C1 (n_3_21), .C2 (n_3_26) );
AOI211_X1 g_8_10 (.ZN (n_8_10), .A (n_5_13), .B (n_1_18), .C1 (n_1_20), .C2 (n_2_24) );
AOI211_X1 g_10_9 (.ZN (n_10_9), .A (n_6_11), .B (n_2_16), .C1 (n_3_19), .C2 (n_1_22) );
AOI211_X1 g_12_8 (.ZN (n_12_8), .A (n_8_10), .B (n_3_14), .C1 (n_1_18), .C2 (n_3_21) );
AOI211_X1 g_14_7 (.ZN (n_14_7), .A (n_10_9), .B (n_5_13), .C1 (n_2_16), .C2 (n_1_20) );
AOI211_X1 g_13_9 (.ZN (n_13_9), .A (n_12_8), .B (n_6_11), .C1 (n_3_14), .C2 (n_3_19) );
AOI211_X1 g_11_8 (.ZN (n_11_8), .A (n_14_7), .B (n_8_10), .C1 (n_5_13), .C2 (n_1_18) );
AOI211_X1 g_13_7 (.ZN (n_13_7), .A (n_13_9), .B (n_10_9), .C1 (n_6_11), .C2 (n_2_16) );
AOI211_X1 g_15_6 (.ZN (n_15_6), .A (n_11_8), .B (n_12_8), .C1 (n_8_10), .C2 (n_3_14) );
AOI211_X1 g_17_5 (.ZN (n_17_5), .A (n_13_7), .B (n_14_7), .C1 (n_10_9), .C2 (n_5_13) );
AOI211_X1 g_19_4 (.ZN (n_19_4), .A (n_15_6), .B (n_13_9), .C1 (n_12_8), .C2 (n_6_11) );
AOI211_X1 g_21_3 (.ZN (n_21_3), .A (n_17_5), .B (n_11_8), .C1 (n_14_7), .C2 (n_8_10) );
AOI211_X1 g_23_2 (.ZN (n_23_2), .A (n_19_4), .B (n_13_7), .C1 (n_13_9), .C2 (n_10_9) );
AOI211_X1 g_25_1 (.ZN (n_25_1), .A (n_21_3), .B (n_15_6), .C1 (n_11_8), .C2 (n_12_8) );
AOI211_X1 g_24_3 (.ZN (n_24_3), .A (n_23_2), .B (n_17_5), .C1 (n_13_7), .C2 (n_14_7) );
AOI211_X1 g_26_2 (.ZN (n_26_2), .A (n_25_1), .B (n_19_4), .C1 (n_15_6), .C2 (n_13_9) );
AOI211_X1 g_28_1 (.ZN (n_28_1), .A (n_24_3), .B (n_21_3), .C1 (n_17_5), .C2 (n_11_8) );
AOI211_X1 g_27_3 (.ZN (n_27_3), .A (n_26_2), .B (n_23_2), .C1 (n_19_4), .C2 (n_13_7) );
AOI211_X1 g_26_1 (.ZN (n_26_1), .A (n_28_1), .B (n_25_1), .C1 (n_21_3), .C2 (n_15_6) );
AOI211_X1 g_24_2 (.ZN (n_24_2), .A (n_27_3), .B (n_24_3), .C1 (n_23_2), .C2 (n_17_5) );
AOI211_X1 g_22_3 (.ZN (n_22_3), .A (n_26_1), .B (n_26_2), .C1 (n_25_1), .C2 (n_19_4) );
AOI211_X1 g_20_4 (.ZN (n_20_4), .A (n_24_2), .B (n_28_1), .C1 (n_24_3), .C2 (n_21_3) );
AOI211_X1 g_18_5 (.ZN (n_18_5), .A (n_22_3), .B (n_27_3), .C1 (n_26_2), .C2 (n_23_2) );
AOI211_X1 g_17_7 (.ZN (n_17_7), .A (n_20_4), .B (n_26_1), .C1 (n_28_1), .C2 (n_25_1) );
AOI211_X1 g_15_8 (.ZN (n_15_8), .A (n_18_5), .B (n_24_2), .C1 (n_27_3), .C2 (n_24_3) );
AOI211_X1 g_14_10 (.ZN (n_14_10), .A (n_17_7), .B (n_22_3), .C1 (n_26_1), .C2 (n_26_2) );
AOI211_X1 g_12_9 (.ZN (n_12_9), .A (n_15_8), .B (n_20_4), .C1 (n_24_2), .C2 (n_28_1) );
AOI211_X1 g_14_8 (.ZN (n_14_8), .A (n_14_10), .B (n_18_5), .C1 (n_22_3), .C2 (n_27_3) );
AOI211_X1 g_16_7 (.ZN (n_16_7), .A (n_12_9), .B (n_17_7), .C1 (n_20_4), .C2 (n_26_1) );
AOI211_X1 g_18_6 (.ZN (n_18_6), .A (n_14_8), .B (n_15_8), .C1 (n_18_5), .C2 (n_24_2) );
AOI211_X1 g_20_5 (.ZN (n_20_5), .A (n_16_7), .B (n_14_10), .C1 (n_17_7), .C2 (n_22_3) );
AOI211_X1 g_22_4 (.ZN (n_22_4), .A (n_18_6), .B (n_12_9), .C1 (n_15_8), .C2 (n_20_4) );
AOI211_X1 g_21_6 (.ZN (n_21_6), .A (n_20_5), .B (n_14_8), .C1 (n_14_10), .C2 (n_18_5) );
AOI211_X1 g_23_5 (.ZN (n_23_5), .A (n_22_4), .B (n_16_7), .C1 (n_12_9), .C2 (n_17_7) );
AOI211_X1 g_25_4 (.ZN (n_25_4), .A (n_21_6), .B (n_18_6), .C1 (n_14_8), .C2 (n_15_8) );
AOI211_X1 g_24_6 (.ZN (n_24_6), .A (n_23_5), .B (n_20_5), .C1 (n_16_7), .C2 (n_14_10) );
AOI211_X1 g_23_4 (.ZN (n_23_4), .A (n_25_4), .B (n_22_4), .C1 (n_18_6), .C2 (n_12_9) );
AOI211_X1 g_25_3 (.ZN (n_25_3), .A (n_24_6), .B (n_21_6), .C1 (n_20_5), .C2 (n_14_8) );
AOI211_X1 g_27_2 (.ZN (n_27_2), .A (n_23_4), .B (n_23_5), .C1 (n_22_4), .C2 (n_16_7) );
AOI211_X1 g_29_1 (.ZN (n_29_1), .A (n_25_3), .B (n_25_4), .C1 (n_21_6), .C2 (n_18_6) );
AOI211_X1 g_28_3 (.ZN (n_28_3), .A (n_27_2), .B (n_24_6), .C1 (n_23_5), .C2 (n_20_5) );
AOI211_X1 g_30_2 (.ZN (n_30_2), .A (n_29_1), .B (n_23_4), .C1 (n_25_4), .C2 (n_22_4) );
AOI211_X1 g_32_1 (.ZN (n_32_1), .A (n_28_3), .B (n_25_3), .C1 (n_24_6), .C2 (n_21_6) );
AOI211_X1 g_31_3 (.ZN (n_31_3), .A (n_30_2), .B (n_27_2), .C1 (n_23_4), .C2 (n_23_5) );
AOI211_X1 g_30_1 (.ZN (n_30_1), .A (n_32_1), .B (n_29_1), .C1 (n_25_3), .C2 (n_25_4) );
AOI211_X1 g_28_2 (.ZN (n_28_2), .A (n_31_3), .B (n_28_3), .C1 (n_27_2), .C2 (n_24_6) );
AOI211_X1 g_26_3 (.ZN (n_26_3), .A (n_30_1), .B (n_30_2), .C1 (n_29_1), .C2 (n_23_4) );
AOI211_X1 g_24_4 (.ZN (n_24_4), .A (n_28_2), .B (n_32_1), .C1 (n_28_3), .C2 (n_25_3) );
AOI211_X1 g_22_5 (.ZN (n_22_5), .A (n_26_3), .B (n_31_3), .C1 (n_30_2), .C2 (n_27_2) );
AOI211_X1 g_20_6 (.ZN (n_20_6), .A (n_24_4), .B (n_30_1), .C1 (n_32_1), .C2 (n_29_1) );
AOI211_X1 g_18_7 (.ZN (n_18_7), .A (n_22_5), .B (n_28_2), .C1 (n_31_3), .C2 (n_28_3) );
AOI211_X1 g_16_8 (.ZN (n_16_8), .A (n_20_6), .B (n_26_3), .C1 (n_30_1), .C2 (n_30_2) );
AOI211_X1 g_14_9 (.ZN (n_14_9), .A (n_18_7), .B (n_24_4), .C1 (n_28_2), .C2 (n_32_1) );
AOI211_X1 g_12_10 (.ZN (n_12_10), .A (n_16_8), .B (n_22_5), .C1 (n_26_3), .C2 (n_31_3) );
AOI211_X1 g_10_11 (.ZN (n_10_11), .A (n_14_9), .B (n_20_6), .C1 (n_24_4), .C2 (n_30_1) );
AOI211_X1 g_9_9 (.ZN (n_9_9), .A (n_12_10), .B (n_18_7), .C1 (n_22_5), .C2 (n_28_2) );
AOI211_X1 g_7_10 (.ZN (n_7_10), .A (n_10_11), .B (n_16_8), .C1 (n_20_6), .C2 (n_26_3) );
AOI211_X1 g_5_11 (.ZN (n_5_11), .A (n_9_9), .B (n_14_9), .C1 (n_18_7), .C2 (n_24_4) );
AOI211_X1 g_7_12 (.ZN (n_7_12), .A (n_7_10), .B (n_12_10), .C1 (n_16_8), .C2 (n_22_5) );
AOI211_X1 g_9_11 (.ZN (n_9_11), .A (n_5_11), .B (n_10_11), .C1 (n_14_9), .C2 (n_20_6) );
AOI211_X1 g_11_10 (.ZN (n_11_10), .A (n_7_12), .B (n_9_9), .C1 (n_12_10), .C2 (n_18_7) );
AOI211_X1 g_13_11 (.ZN (n_13_11), .A (n_9_11), .B (n_7_10), .C1 (n_10_11), .C2 (n_16_8) );
AOI211_X1 g_15_10 (.ZN (n_15_10), .A (n_11_10), .B (n_5_11), .C1 (n_9_9), .C2 (n_14_9) );
AOI211_X1 g_17_9 (.ZN (n_17_9), .A (n_13_11), .B (n_7_12), .C1 (n_7_10), .C2 (n_12_10) );
AOI211_X1 g_19_8 (.ZN (n_19_8), .A (n_15_10), .B (n_9_11), .C1 (n_5_11), .C2 (n_10_11) );
AOI211_X1 g_21_7 (.ZN (n_21_7), .A (n_17_9), .B (n_11_10), .C1 (n_7_12), .C2 (n_9_9) );
AOI211_X1 g_19_6 (.ZN (n_19_6), .A (n_19_8), .B (n_13_11), .C1 (n_9_11), .C2 (n_7_10) );
AOI211_X1 g_21_5 (.ZN (n_21_5), .A (n_21_7), .B (n_15_10), .C1 (n_11_10), .C2 (n_5_11) );
AOI211_X1 g_22_7 (.ZN (n_22_7), .A (n_19_6), .B (n_17_9), .C1 (n_13_11), .C2 (n_7_12) );
AOI211_X1 g_20_8 (.ZN (n_20_8), .A (n_21_5), .B (n_19_8), .C1 (n_15_10), .C2 (n_9_11) );
AOI211_X1 g_18_9 (.ZN (n_18_9), .A (n_22_7), .B (n_21_7), .C1 (n_17_9), .C2 (n_11_10) );
AOI211_X1 g_19_7 (.ZN (n_19_7), .A (n_20_8), .B (n_19_6), .C1 (n_19_8), .C2 (n_13_11) );
AOI211_X1 g_17_8 (.ZN (n_17_8), .A (n_18_9), .B (n_21_5), .C1 (n_21_7), .C2 (n_15_10) );
AOI211_X1 g_15_9 (.ZN (n_15_9), .A (n_19_7), .B (n_22_7), .C1 (n_19_6), .C2 (n_17_9) );
AOI211_X1 g_13_10 (.ZN (n_13_10), .A (n_17_8), .B (n_20_8), .C1 (n_21_5), .C2 (n_19_8) );
AOI211_X1 g_11_11 (.ZN (n_11_11), .A (n_15_9), .B (n_18_9), .C1 (n_22_7), .C2 (n_21_7) );
AOI211_X1 g_9_12 (.ZN (n_9_12), .A (n_13_10), .B (n_19_7), .C1 (n_20_8), .C2 (n_19_6) );
AOI211_X1 g_10_10 (.ZN (n_10_10), .A (n_11_11), .B (n_17_8), .C1 (n_18_9), .C2 (n_21_5) );
AOI211_X1 g_8_11 (.ZN (n_8_11), .A (n_9_12), .B (n_15_9), .C1 (n_19_7), .C2 (n_22_7) );
AOI211_X1 g_6_12 (.ZN (n_6_12), .A (n_10_10), .B (n_13_10), .C1 (n_17_8), .C2 (n_20_8) );
AOI211_X1 g_4_13 (.ZN (n_4_13), .A (n_8_11), .B (n_11_11), .C1 (n_15_9), .C2 (n_18_9) );
AOI211_X1 g_2_14 (.ZN (n_2_14), .A (n_6_12), .B (n_9_12), .C1 (n_13_10), .C2 (n_19_7) );
AOI211_X1 g_1_16 (.ZN (n_1_16), .A (n_4_13), .B (n_10_10), .C1 (n_11_11), .C2 (n_17_8) );
AOI211_X1 g_3_15 (.ZN (n_3_15), .A (n_2_14), .B (n_8_11), .C1 (n_9_12), .C2 (n_15_9) );
AOI211_X1 g_5_14 (.ZN (n_5_14), .A (n_1_16), .B (n_6_12), .C1 (n_10_10), .C2 (n_13_10) );
AOI211_X1 g_7_13 (.ZN (n_7_13), .A (n_3_15), .B (n_4_13), .C1 (n_8_11), .C2 (n_11_11) );
AOI211_X1 g_6_15 (.ZN (n_6_15), .A (n_5_14), .B (n_2_14), .C1 (n_6_12), .C2 (n_9_12) );
AOI211_X1 g_4_14 (.ZN (n_4_14), .A (n_7_13), .B (n_1_16), .C1 (n_4_13), .C2 (n_10_10) );
AOI211_X1 g_6_13 (.ZN (n_6_13), .A (n_6_15), .B (n_3_15), .C1 (n_2_14), .C2 (n_8_11) );
AOI211_X1 g_8_12 (.ZN (n_8_12), .A (n_4_14), .B (n_5_14), .C1 (n_1_16), .C2 (n_6_12) );
AOI211_X1 g_7_14 (.ZN (n_7_14), .A (n_6_13), .B (n_7_13), .C1 (n_3_15), .C2 (n_4_13) );
AOI211_X1 g_9_13 (.ZN (n_9_13), .A (n_8_12), .B (n_6_15), .C1 (n_5_14), .C2 (n_2_14) );
AOI211_X1 g_11_12 (.ZN (n_11_12), .A (n_7_14), .B (n_4_14), .C1 (n_7_13), .C2 (n_1_16) );
AOI211_X1 g_10_14 (.ZN (n_10_14), .A (n_9_13), .B (n_6_13), .C1 (n_6_15), .C2 (n_3_15) );
AOI211_X1 g_8_13 (.ZN (n_8_13), .A (n_11_12), .B (n_8_12), .C1 (n_4_14), .C2 (n_5_14) );
AOI211_X1 g_10_12 (.ZN (n_10_12), .A (n_10_14), .B (n_7_14), .C1 (n_6_13), .C2 (n_7_13) );
AOI211_X1 g_12_11 (.ZN (n_12_11), .A (n_8_13), .B (n_9_13), .C1 (n_8_12), .C2 (n_6_15) );
AOI211_X1 g_11_13 (.ZN (n_11_13), .A (n_10_12), .B (n_11_12), .C1 (n_7_14), .C2 (n_4_14) );
AOI211_X1 g_13_12 (.ZN (n_13_12), .A (n_12_11), .B (n_10_14), .C1 (n_9_13), .C2 (n_6_13) );
AOI211_X1 g_15_11 (.ZN (n_15_11), .A (n_11_13), .B (n_8_13), .C1 (n_11_12), .C2 (n_8_12) );
AOI211_X1 g_16_9 (.ZN (n_16_9), .A (n_13_12), .B (n_10_12), .C1 (n_10_14), .C2 (n_7_14) );
AOI211_X1 g_18_8 (.ZN (n_18_8), .A (n_15_11), .B (n_12_11), .C1 (n_8_13), .C2 (n_9_13) );
AOI211_X1 g_20_7 (.ZN (n_20_7), .A (n_16_9), .B (n_11_13), .C1 (n_10_12), .C2 (n_11_12) );
AOI211_X1 g_22_6 (.ZN (n_22_6), .A (n_18_8), .B (n_13_12), .C1 (n_12_11), .C2 (n_10_14) );
AOI211_X1 g_24_5 (.ZN (n_24_5), .A (n_20_7), .B (n_15_11), .C1 (n_11_13), .C2 (n_8_13) );
AOI211_X1 g_26_4 (.ZN (n_26_4), .A (n_22_6), .B (n_16_9), .C1 (n_13_12), .C2 (n_10_12) );
AOI211_X1 g_25_6 (.ZN (n_25_6), .A (n_24_5), .B (n_18_8), .C1 (n_15_11), .C2 (n_12_11) );
AOI211_X1 g_27_5 (.ZN (n_27_5), .A (n_26_4), .B (n_20_7), .C1 (n_16_9), .C2 (n_11_13) );
AOI211_X1 g_29_4 (.ZN (n_29_4), .A (n_25_6), .B (n_22_6), .C1 (n_18_8), .C2 (n_13_12) );
AOI211_X1 g_28_6 (.ZN (n_28_6), .A (n_27_5), .B (n_24_5), .C1 (n_20_7), .C2 (n_15_11) );
AOI211_X1 g_26_5 (.ZN (n_26_5), .A (n_29_4), .B (n_26_4), .C1 (n_22_6), .C2 (n_16_9) );
AOI211_X1 g_28_4 (.ZN (n_28_4), .A (n_28_6), .B (n_25_6), .C1 (n_24_5), .C2 (n_18_8) );
AOI211_X1 g_30_3 (.ZN (n_30_3), .A (n_26_5), .B (n_27_5), .C1 (n_26_4), .C2 (n_20_7) );
AOI211_X1 g_32_2 (.ZN (n_32_2), .A (n_28_4), .B (n_29_4), .C1 (n_25_6), .C2 (n_22_6) );
AOI211_X1 g_34_1 (.ZN (n_34_1), .A (n_30_3), .B (n_28_6), .C1 (n_27_5), .C2 (n_24_5) );
AOI211_X1 g_35_3 (.ZN (n_35_3), .A (n_32_2), .B (n_26_5), .C1 (n_29_4), .C2 (n_26_4) );
AOI211_X1 g_36_1 (.ZN (n_36_1), .A (n_34_1), .B (n_28_4), .C1 (n_28_6), .C2 (n_25_6) );
AOI211_X1 g_34_2 (.ZN (n_34_2), .A (n_35_3), .B (n_30_3), .C1 (n_26_5), .C2 (n_27_5) );
AOI211_X1 g_33_4 (.ZN (n_33_4), .A (n_36_1), .B (n_32_2), .C1 (n_28_4), .C2 (n_29_4) );
AOI211_X1 g_31_5 (.ZN (n_31_5), .A (n_34_2), .B (n_34_1), .C1 (n_30_3), .C2 (n_28_6) );
AOI211_X1 g_32_3 (.ZN (n_32_3), .A (n_33_4), .B (n_35_3), .C1 (n_32_2), .C2 (n_26_5) );
AOI211_X1 g_33_1 (.ZN (n_33_1), .A (n_31_5), .B (n_36_1), .C1 (n_34_1), .C2 (n_28_4) );
AOI211_X1 g_31_2 (.ZN (n_31_2), .A (n_32_3), .B (n_34_2), .C1 (n_35_3), .C2 (n_30_3) );
AOI211_X1 g_29_3 (.ZN (n_29_3), .A (n_33_1), .B (n_33_4), .C1 (n_36_1), .C2 (n_32_2) );
AOI211_X1 g_27_4 (.ZN (n_27_4), .A (n_31_2), .B (n_31_5), .C1 (n_34_2), .C2 (n_34_1) );
AOI211_X1 g_25_5 (.ZN (n_25_5), .A (n_29_3), .B (n_32_3), .C1 (n_33_4), .C2 (n_35_3) );
AOI211_X1 g_23_6 (.ZN (n_23_6), .A (n_27_4), .B (n_33_1), .C1 (n_31_5), .C2 (n_36_1) );
AOI211_X1 g_22_8 (.ZN (n_22_8), .A (n_25_5), .B (n_31_2), .C1 (n_32_3), .C2 (n_34_2) );
AOI211_X1 g_24_7 (.ZN (n_24_7), .A (n_23_6), .B (n_29_3), .C1 (n_33_1), .C2 (n_33_4) );
AOI211_X1 g_26_6 (.ZN (n_26_6), .A (n_22_8), .B (n_27_4), .C1 (n_31_2), .C2 (n_31_5) );
AOI211_X1 g_28_5 (.ZN (n_28_5), .A (n_24_7), .B (n_25_5), .C1 (n_29_3), .C2 (n_32_3) );
AOI211_X1 g_30_4 (.ZN (n_30_4), .A (n_26_6), .B (n_23_6), .C1 (n_27_4), .C2 (n_33_1) );
AOI211_X1 g_29_6 (.ZN (n_29_6), .A (n_28_5), .B (n_22_8), .C1 (n_25_5), .C2 (n_31_2) );
AOI211_X1 g_27_7 (.ZN (n_27_7), .A (n_30_4), .B (n_24_7), .C1 (n_23_6), .C2 (n_29_3) );
AOI211_X1 g_25_8 (.ZN (n_25_8), .A (n_29_6), .B (n_26_6), .C1 (n_22_8), .C2 (n_27_4) );
AOI211_X1 g_23_7 (.ZN (n_23_7), .A (n_27_7), .B (n_28_5), .C1 (n_24_7), .C2 (n_25_5) );
AOI211_X1 g_21_8 (.ZN (n_21_8), .A (n_25_8), .B (n_30_4), .C1 (n_26_6), .C2 (n_23_6) );
AOI211_X1 g_19_9 (.ZN (n_19_9), .A (n_23_7), .B (n_29_6), .C1 (n_28_5), .C2 (n_22_8) );
AOI211_X1 g_17_10 (.ZN (n_17_10), .A (n_21_8), .B (n_27_7), .C1 (n_30_4), .C2 (n_24_7) );
AOI211_X1 g_16_12 (.ZN (n_16_12), .A (n_19_9), .B (n_25_8), .C1 (n_29_6), .C2 (n_26_6) );
AOI211_X1 g_14_11 (.ZN (n_14_11), .A (n_17_10), .B (n_23_7), .C1 (n_27_7), .C2 (n_28_5) );
AOI211_X1 g_16_10 (.ZN (n_16_10), .A (n_16_12), .B (n_21_8), .C1 (n_25_8), .C2 (n_30_4) );
AOI211_X1 g_18_11 (.ZN (n_18_11), .A (n_14_11), .B (n_19_9), .C1 (n_23_7), .C2 (n_29_6) );
AOI211_X1 g_20_10 (.ZN (n_20_10), .A (n_16_10), .B (n_17_10), .C1 (n_21_8), .C2 (n_27_7) );
AOI211_X1 g_22_9 (.ZN (n_22_9), .A (n_18_11), .B (n_16_12), .C1 (n_19_9), .C2 (n_25_8) );
AOI211_X1 g_24_8 (.ZN (n_24_8), .A (n_20_10), .B (n_14_11), .C1 (n_17_10), .C2 (n_23_7) );
AOI211_X1 g_26_7 (.ZN (n_26_7), .A (n_22_9), .B (n_16_10), .C1 (n_16_12), .C2 (n_21_8) );
AOI211_X1 g_25_9 (.ZN (n_25_9), .A (n_24_8), .B (n_18_11), .C1 (n_14_11), .C2 (n_19_9) );
AOI211_X1 g_23_8 (.ZN (n_23_8), .A (n_26_7), .B (n_20_10), .C1 (n_16_10), .C2 (n_17_10) );
AOI211_X1 g_25_7 (.ZN (n_25_7), .A (n_25_9), .B (n_22_9), .C1 (n_18_11), .C2 (n_16_12) );
AOI211_X1 g_27_6 (.ZN (n_27_6), .A (n_23_8), .B (n_24_8), .C1 (n_20_10), .C2 (n_14_11) );
AOI211_X1 g_29_5 (.ZN (n_29_5), .A (n_25_7), .B (n_26_7), .C1 (n_22_9), .C2 (n_16_10) );
AOI211_X1 g_31_4 (.ZN (n_31_4), .A (n_27_6), .B (n_25_9), .C1 (n_24_8), .C2 (n_18_11) );
AOI211_X1 g_33_3 (.ZN (n_33_3), .A (n_29_5), .B (n_23_8), .C1 (n_26_7), .C2 (n_20_10) );
AOI211_X1 g_35_2 (.ZN (n_35_2), .A (n_31_4), .B (n_25_7), .C1 (n_25_9), .C2 (n_22_9) );
AOI211_X1 g_37_1 (.ZN (n_37_1), .A (n_33_3), .B (n_27_6), .C1 (n_23_8), .C2 (n_24_8) );
AOI211_X1 g_36_3 (.ZN (n_36_3), .A (n_35_2), .B (n_29_5), .C1 (n_25_7), .C2 (n_26_7) );
AOI211_X1 g_38_2 (.ZN (n_38_2), .A (n_37_1), .B (n_31_4), .C1 (n_27_6), .C2 (n_25_9) );
AOI211_X1 g_40_1 (.ZN (n_40_1), .A (n_36_3), .B (n_33_3), .C1 (n_29_5), .C2 (n_23_8) );
AOI211_X1 g_39_3 (.ZN (n_39_3), .A (n_38_2), .B (n_35_2), .C1 (n_31_4), .C2 (n_25_7) );
AOI211_X1 g_38_1 (.ZN (n_38_1), .A (n_40_1), .B (n_37_1), .C1 (n_33_3), .C2 (n_27_6) );
AOI211_X1 g_36_2 (.ZN (n_36_2), .A (n_39_3), .B (n_36_3), .C1 (n_35_2), .C2 (n_29_5) );
AOI211_X1 g_34_3 (.ZN (n_34_3), .A (n_38_1), .B (n_38_2), .C1 (n_37_1), .C2 (n_31_4) );
AOI211_X1 g_32_4 (.ZN (n_32_4), .A (n_36_2), .B (n_40_1), .C1 (n_36_3), .C2 (n_33_3) );
AOI211_X1 g_30_5 (.ZN (n_30_5), .A (n_34_3), .B (n_39_3), .C1 (n_38_2), .C2 (n_35_2) );
AOI211_X1 g_29_7 (.ZN (n_29_7), .A (n_32_4), .B (n_38_1), .C1 (n_40_1), .C2 (n_37_1) );
AOI211_X1 g_27_8 (.ZN (n_27_8), .A (n_30_5), .B (n_36_2), .C1 (n_39_3), .C2 (n_36_3) );
AOI211_X1 g_26_10 (.ZN (n_26_10), .A (n_29_7), .B (n_34_3), .C1 (n_38_1), .C2 (n_38_2) );
AOI211_X1 g_24_9 (.ZN (n_24_9), .A (n_27_8), .B (n_32_4), .C1 (n_36_2), .C2 (n_40_1) );
AOI211_X1 g_26_8 (.ZN (n_26_8), .A (n_26_10), .B (n_30_5), .C1 (n_34_3), .C2 (n_39_3) );
AOI211_X1 g_28_7 (.ZN (n_28_7), .A (n_24_9), .B (n_29_7), .C1 (n_32_4), .C2 (n_38_1) );
AOI211_X1 g_30_6 (.ZN (n_30_6), .A (n_26_8), .B (n_27_8), .C1 (n_30_5), .C2 (n_36_2) );
AOI211_X1 g_32_5 (.ZN (n_32_5), .A (n_28_7), .B (n_26_10), .C1 (n_29_7), .C2 (n_34_3) );
AOI211_X1 g_34_4 (.ZN (n_34_4), .A (n_30_6), .B (n_24_9), .C1 (n_27_8), .C2 (n_32_4) );
AOI211_X1 g_33_6 (.ZN (n_33_6), .A (n_32_5), .B (n_26_8), .C1 (n_26_10), .C2 (n_30_5) );
AOI211_X1 g_35_5 (.ZN (n_35_5), .A (n_34_4), .B (n_28_7), .C1 (n_24_9), .C2 (n_29_7) );
AOI211_X1 g_37_4 (.ZN (n_37_4), .A (n_33_6), .B (n_30_6), .C1 (n_26_8), .C2 (n_27_8) );
AOI211_X1 g_36_6 (.ZN (n_36_6), .A (n_35_5), .B (n_32_5), .C1 (n_28_7), .C2 (n_26_10) );
AOI211_X1 g_35_4 (.ZN (n_35_4), .A (n_37_4), .B (n_34_4), .C1 (n_30_6), .C2 (n_24_9) );
AOI211_X1 g_37_3 (.ZN (n_37_3), .A (n_36_6), .B (n_33_6), .C1 (n_32_5), .C2 (n_26_8) );
AOI211_X1 g_39_2 (.ZN (n_39_2), .A (n_35_4), .B (n_35_5), .C1 (n_34_4), .C2 (n_28_7) );
AOI211_X1 g_41_1 (.ZN (n_41_1), .A (n_37_3), .B (n_37_4), .C1 (n_33_6), .C2 (n_30_6) );
AOI211_X1 g_40_3 (.ZN (n_40_3), .A (n_39_2), .B (n_36_6), .C1 (n_35_5), .C2 (n_32_5) );
AOI211_X1 g_42_2 (.ZN (n_42_2), .A (n_41_1), .B (n_35_4), .C1 (n_37_4), .C2 (n_34_4) );
AOI211_X1 g_44_1 (.ZN (n_44_1), .A (n_40_3), .B (n_37_3), .C1 (n_36_6), .C2 (n_33_6) );
AOI211_X1 g_43_3 (.ZN (n_43_3), .A (n_42_2), .B (n_39_2), .C1 (n_35_4), .C2 (n_35_5) );
AOI211_X1 g_42_1 (.ZN (n_42_1), .A (n_44_1), .B (n_41_1), .C1 (n_37_3), .C2 (n_37_4) );
AOI211_X1 g_40_2 (.ZN (n_40_2), .A (n_43_3), .B (n_40_3), .C1 (n_39_2), .C2 (n_36_6) );
AOI211_X1 g_38_3 (.ZN (n_38_3), .A (n_42_1), .B (n_42_2), .C1 (n_41_1), .C2 (n_35_4) );
AOI211_X1 g_36_4 (.ZN (n_36_4), .A (n_40_2), .B (n_44_1), .C1 (n_40_3), .C2 (n_37_3) );
AOI211_X1 g_34_5 (.ZN (n_34_5), .A (n_38_3), .B (n_43_3), .C1 (n_42_2), .C2 (n_39_2) );
AOI211_X1 g_32_6 (.ZN (n_32_6), .A (n_36_4), .B (n_42_1), .C1 (n_44_1), .C2 (n_41_1) );
AOI211_X1 g_30_7 (.ZN (n_30_7), .A (n_34_5), .B (n_40_2), .C1 (n_43_3), .C2 (n_40_3) );
AOI211_X1 g_28_8 (.ZN (n_28_8), .A (n_32_6), .B (n_38_3), .C1 (n_42_1), .C2 (n_42_2) );
AOI211_X1 g_26_9 (.ZN (n_26_9), .A (n_30_7), .B (n_36_4), .C1 (n_40_2), .C2 (n_44_1) );
AOI211_X1 g_24_10 (.ZN (n_24_10), .A (n_28_8), .B (n_34_5), .C1 (n_38_3), .C2 (n_43_3) );
AOI211_X1 g_22_11 (.ZN (n_22_11), .A (n_26_9), .B (n_32_6), .C1 (n_36_4), .C2 (n_42_1) );
AOI211_X1 g_23_9 (.ZN (n_23_9), .A (n_24_10), .B (n_30_7), .C1 (n_34_5), .C2 (n_40_2) );
AOI211_X1 g_21_10 (.ZN (n_21_10), .A (n_22_11), .B (n_28_8), .C1 (n_32_6), .C2 (n_38_3) );
AOI211_X1 g_19_11 (.ZN (n_19_11), .A (n_23_9), .B (n_26_9), .C1 (n_30_7), .C2 (n_36_4) );
AOI211_X1 g_20_9 (.ZN (n_20_9), .A (n_21_10), .B (n_24_10), .C1 (n_28_8), .C2 (n_34_5) );
AOI211_X1 g_18_10 (.ZN (n_18_10), .A (n_19_11), .B (n_22_11), .C1 (n_26_9), .C2 (n_32_6) );
AOI211_X1 g_16_11 (.ZN (n_16_11), .A (n_20_9), .B (n_23_9), .C1 (n_24_10), .C2 (n_30_7) );
AOI211_X1 g_14_12 (.ZN (n_14_12), .A (n_18_10), .B (n_21_10), .C1 (n_22_11), .C2 (n_28_8) );
AOI211_X1 g_12_13 (.ZN (n_12_13), .A (n_16_11), .B (n_19_11), .C1 (n_23_9), .C2 (n_26_9) );
AOI211_X1 g_14_14 (.ZN (n_14_14), .A (n_14_12), .B (n_20_9), .C1 (n_21_10), .C2 (n_24_10) );
AOI211_X1 g_15_12 (.ZN (n_15_12), .A (n_12_13), .B (n_18_10), .C1 (n_19_11), .C2 (n_22_11) );
AOI211_X1 g_17_11 (.ZN (n_17_11), .A (n_14_14), .B (n_16_11), .C1 (n_20_9), .C2 (n_23_9) );
AOI211_X1 g_19_10 (.ZN (n_19_10), .A (n_15_12), .B (n_14_12), .C1 (n_18_10), .C2 (n_21_10) );
AOI211_X1 g_21_9 (.ZN (n_21_9), .A (n_17_11), .B (n_12_13), .C1 (n_16_11), .C2 (n_19_11) );
AOI211_X1 g_23_10 (.ZN (n_23_10), .A (n_19_10), .B (n_14_14), .C1 (n_14_12), .C2 (n_20_9) );
AOI211_X1 g_21_11 (.ZN (n_21_11), .A (n_21_9), .B (n_15_12), .C1 (n_12_13), .C2 (n_18_10) );
AOI211_X1 g_19_12 (.ZN (n_19_12), .A (n_23_10), .B (n_17_11), .C1 (n_14_14), .C2 (n_16_11) );
AOI211_X1 g_17_13 (.ZN (n_17_13), .A (n_21_11), .B (n_19_10), .C1 (n_15_12), .C2 (n_14_12) );
AOI211_X1 g_15_14 (.ZN (n_15_14), .A (n_19_12), .B (n_21_9), .C1 (n_17_11), .C2 (n_12_13) );
AOI211_X1 g_13_13 (.ZN (n_13_13), .A (n_17_13), .B (n_23_10), .C1 (n_19_10), .C2 (n_14_14) );
AOI211_X1 g_12_15 (.ZN (n_12_15), .A (n_15_14), .B (n_21_11), .C1 (n_21_9), .C2 (n_15_12) );
AOI211_X1 g_14_16 (.ZN (n_14_16), .A (n_13_13), .B (n_19_12), .C1 (n_23_10), .C2 (n_17_11) );
AOI211_X1 g_16_15 (.ZN (n_16_15), .A (n_12_15), .B (n_17_13), .C1 (n_21_11), .C2 (n_19_10) );
AOI211_X1 g_15_13 (.ZN (n_15_13), .A (n_14_16), .B (n_15_14), .C1 (n_19_12), .C2 (n_21_9) );
AOI211_X1 g_17_12 (.ZN (n_17_12), .A (n_16_15), .B (n_13_13), .C1 (n_17_13), .C2 (n_23_10) );
AOI211_X1 g_18_14 (.ZN (n_18_14), .A (n_15_13), .B (n_12_15), .C1 (n_15_14), .C2 (n_21_11) );
AOI211_X1 g_16_13 (.ZN (n_16_13), .A (n_17_12), .B (n_14_16), .C1 (n_13_13), .C2 (n_19_12) );
AOI211_X1 g_18_12 (.ZN (n_18_12), .A (n_18_14), .B (n_16_15), .C1 (n_12_15), .C2 (n_17_13) );
AOI211_X1 g_20_11 (.ZN (n_20_11), .A (n_16_13), .B (n_15_13), .C1 (n_14_16), .C2 (n_15_14) );
AOI211_X1 g_22_10 (.ZN (n_22_10), .A (n_18_12), .B (n_17_12), .C1 (n_16_15), .C2 (n_13_13) );
AOI211_X1 g_24_11 (.ZN (n_24_11), .A (n_20_11), .B (n_18_14), .C1 (n_15_13), .C2 (n_12_15) );
AOI211_X1 g_22_12 (.ZN (n_22_12), .A (n_22_10), .B (n_16_13), .C1 (n_17_12), .C2 (n_14_16) );
AOI211_X1 g_20_13 (.ZN (n_20_13), .A (n_24_11), .B (n_18_12), .C1 (n_18_14), .C2 (n_16_15) );
AOI211_X1 g_19_15 (.ZN (n_19_15), .A (n_22_12), .B (n_20_11), .C1 (n_16_13), .C2 (n_15_13) );
AOI211_X1 g_18_13 (.ZN (n_18_13), .A (n_20_13), .B (n_22_10), .C1 (n_18_12), .C2 (n_17_12) );
AOI211_X1 g_20_12 (.ZN (n_20_12), .A (n_19_15), .B (n_24_11), .C1 (n_20_11), .C2 (n_18_14) );
AOI211_X1 g_19_14 (.ZN (n_19_14), .A (n_18_13), .B (n_22_12), .C1 (n_22_10), .C2 (n_16_13) );
AOI211_X1 g_21_13 (.ZN (n_21_13), .A (n_20_12), .B (n_20_13), .C1 (n_24_11), .C2 (n_18_12) );
AOI211_X1 g_23_12 (.ZN (n_23_12), .A (n_19_14), .B (n_19_15), .C1 (n_22_12), .C2 (n_20_11) );
AOI211_X1 g_25_11 (.ZN (n_25_11), .A (n_21_13), .B (n_18_13), .C1 (n_20_13), .C2 (n_22_10) );
AOI211_X1 g_27_10 (.ZN (n_27_10), .A (n_23_12), .B (n_20_12), .C1 (n_19_15), .C2 (n_24_11) );
AOI211_X1 g_29_9 (.ZN (n_29_9), .A (n_25_11), .B (n_19_14), .C1 (n_18_13), .C2 (n_22_12) );
AOI211_X1 g_31_8 (.ZN (n_31_8), .A (n_27_10), .B (n_21_13), .C1 (n_20_12), .C2 (n_20_13) );
AOI211_X1 g_33_7 (.ZN (n_33_7), .A (n_29_9), .B (n_23_12), .C1 (n_19_14), .C2 (n_19_15) );
AOI211_X1 g_31_6 (.ZN (n_31_6), .A (n_31_8), .B (n_25_11), .C1 (n_21_13), .C2 (n_18_13) );
AOI211_X1 g_33_5 (.ZN (n_33_5), .A (n_33_7), .B (n_27_10), .C1 (n_23_12), .C2 (n_20_12) );
AOI211_X1 g_34_7 (.ZN (n_34_7), .A (n_31_6), .B (n_29_9), .C1 (n_25_11), .C2 (n_19_14) );
AOI211_X1 g_32_8 (.ZN (n_32_8), .A (n_33_5), .B (n_31_8), .C1 (n_27_10), .C2 (n_21_13) );
AOI211_X1 g_30_9 (.ZN (n_30_9), .A (n_34_7), .B (n_33_7), .C1 (n_29_9), .C2 (n_23_12) );
AOI211_X1 g_31_7 (.ZN (n_31_7), .A (n_32_8), .B (n_31_6), .C1 (n_31_8), .C2 (n_25_11) );
AOI211_X1 g_29_8 (.ZN (n_29_8), .A (n_30_9), .B (n_33_5), .C1 (n_33_7), .C2 (n_27_10) );
AOI211_X1 g_27_9 (.ZN (n_27_9), .A (n_31_7), .B (n_34_7), .C1 (n_31_6), .C2 (n_29_9) );
AOI211_X1 g_25_10 (.ZN (n_25_10), .A (n_29_8), .B (n_32_8), .C1 (n_33_5), .C2 (n_31_8) );
AOI211_X1 g_23_11 (.ZN (n_23_11), .A (n_27_9), .B (n_30_9), .C1 (n_34_7), .C2 (n_33_7) );
AOI211_X1 g_21_12 (.ZN (n_21_12), .A (n_25_10), .B (n_31_7), .C1 (n_32_8), .C2 (n_31_6) );
AOI211_X1 g_19_13 (.ZN (n_19_13), .A (n_23_11), .B (n_29_8), .C1 (n_30_9), .C2 (n_33_5) );
AOI211_X1 g_17_14 (.ZN (n_17_14), .A (n_21_12), .B (n_27_9), .C1 (n_31_7), .C2 (n_34_7) );
AOI211_X1 g_18_16 (.ZN (n_18_16), .A (n_19_13), .B (n_25_10), .C1 (n_29_8), .C2 (n_32_8) );
AOI211_X1 g_20_15 (.ZN (n_20_15), .A (n_17_14), .B (n_23_11), .C1 (n_27_9), .C2 (n_30_9) );
AOI211_X1 g_22_14 (.ZN (n_22_14), .A (n_18_16), .B (n_21_12), .C1 (n_25_10), .C2 (n_31_7) );
AOI211_X1 g_24_13 (.ZN (n_24_13), .A (n_20_15), .B (n_19_13), .C1 (n_23_11), .C2 (n_29_8) );
AOI211_X1 g_26_12 (.ZN (n_26_12), .A (n_22_14), .B (n_17_14), .C1 (n_21_12), .C2 (n_27_9) );
AOI211_X1 g_28_11 (.ZN (n_28_11), .A (n_24_13), .B (n_18_16), .C1 (n_19_13), .C2 (n_25_10) );
AOI211_X1 g_30_10 (.ZN (n_30_10), .A (n_26_12), .B (n_20_15), .C1 (n_17_14), .C2 (n_23_11) );
AOI211_X1 g_28_9 (.ZN (n_28_9), .A (n_28_11), .B (n_22_14), .C1 (n_18_16), .C2 (n_21_12) );
AOI211_X1 g_30_8 (.ZN (n_30_8), .A (n_30_10), .B (n_24_13), .C1 (n_20_15), .C2 (n_19_13) );
AOI211_X1 g_32_7 (.ZN (n_32_7), .A (n_28_9), .B (n_26_12), .C1 (n_22_14), .C2 (n_17_14) );
AOI211_X1 g_34_6 (.ZN (n_34_6), .A (n_30_8), .B (n_28_11), .C1 (n_24_13), .C2 (n_18_16) );
AOI211_X1 g_36_5 (.ZN (n_36_5), .A (n_32_7), .B (n_30_10), .C1 (n_26_12), .C2 (n_20_15) );
AOI211_X1 g_38_4 (.ZN (n_38_4), .A (n_34_6), .B (n_28_9), .C1 (n_28_11), .C2 (n_22_14) );
AOI211_X1 g_37_6 (.ZN (n_37_6), .A (n_36_5), .B (n_30_8), .C1 (n_30_10), .C2 (n_24_13) );
AOI211_X1 g_39_5 (.ZN (n_39_5), .A (n_38_4), .B (n_32_7), .C1 (n_28_9), .C2 (n_26_12) );
AOI211_X1 g_41_4 (.ZN (n_41_4), .A (n_37_6), .B (n_34_6), .C1 (n_30_8), .C2 (n_28_11) );
AOI211_X1 g_40_6 (.ZN (n_40_6), .A (n_39_5), .B (n_36_5), .C1 (n_32_7), .C2 (n_30_10) );
AOI211_X1 g_38_5 (.ZN (n_38_5), .A (n_41_4), .B (n_38_4), .C1 (n_34_6), .C2 (n_28_9) );
AOI211_X1 g_40_4 (.ZN (n_40_4), .A (n_40_6), .B (n_37_6), .C1 (n_36_5), .C2 (n_30_8) );
AOI211_X1 g_42_3 (.ZN (n_42_3), .A (n_38_5), .B (n_39_5), .C1 (n_38_4), .C2 (n_32_7) );
AOI211_X1 g_44_2 (.ZN (n_44_2), .A (n_40_4), .B (n_41_4), .C1 (n_37_6), .C2 (n_34_6) );
AOI211_X1 g_46_1 (.ZN (n_46_1), .A (n_42_3), .B (n_40_6), .C1 (n_39_5), .C2 (n_36_5) );
AOI211_X1 g_47_3 (.ZN (n_47_3), .A (n_44_2), .B (n_38_5), .C1 (n_41_4), .C2 (n_38_4) );
AOI211_X1 g_48_1 (.ZN (n_48_1), .A (n_46_1), .B (n_40_4), .C1 (n_40_6), .C2 (n_37_6) );
AOI211_X1 g_46_2 (.ZN (n_46_2), .A (n_47_3), .B (n_42_3), .C1 (n_38_5), .C2 (n_39_5) );
AOI211_X1 g_45_4 (.ZN (n_45_4), .A (n_48_1), .B (n_44_2), .C1 (n_40_4), .C2 (n_41_4) );
AOI211_X1 g_43_5 (.ZN (n_43_5), .A (n_46_2), .B (n_46_1), .C1 (n_42_3), .C2 (n_40_6) );
AOI211_X1 g_44_3 (.ZN (n_44_3), .A (n_45_4), .B (n_47_3), .C1 (n_44_2), .C2 (n_38_5) );
AOI211_X1 g_45_1 (.ZN (n_45_1), .A (n_43_5), .B (n_48_1), .C1 (n_46_1), .C2 (n_40_4) );
AOI211_X1 g_43_2 (.ZN (n_43_2), .A (n_44_3), .B (n_46_2), .C1 (n_47_3), .C2 (n_42_3) );
AOI211_X1 g_41_3 (.ZN (n_41_3), .A (n_45_1), .B (n_45_4), .C1 (n_48_1), .C2 (n_44_2) );
AOI211_X1 g_39_4 (.ZN (n_39_4), .A (n_43_2), .B (n_43_5), .C1 (n_46_2), .C2 (n_46_1) );
AOI211_X1 g_37_5 (.ZN (n_37_5), .A (n_41_3), .B (n_44_3), .C1 (n_45_4), .C2 (n_47_3) );
AOI211_X1 g_35_6 (.ZN (n_35_6), .A (n_39_4), .B (n_45_1), .C1 (n_43_5), .C2 (n_48_1) );
AOI211_X1 g_34_8 (.ZN (n_34_8), .A (n_37_5), .B (n_43_2), .C1 (n_44_3), .C2 (n_46_2) );
AOI211_X1 g_32_9 (.ZN (n_32_9), .A (n_35_6), .B (n_41_3), .C1 (n_45_1), .C2 (n_45_4) );
AOI211_X1 g_31_11 (.ZN (n_31_11), .A (n_34_8), .B (n_39_4), .C1 (n_43_2), .C2 (n_43_5) );
AOI211_X1 g_29_10 (.ZN (n_29_10), .A (n_32_9), .B (n_37_5), .C1 (n_41_3), .C2 (n_44_3) );
AOI211_X1 g_31_9 (.ZN (n_31_9), .A (n_31_11), .B (n_35_6), .C1 (n_39_4), .C2 (n_45_1) );
AOI211_X1 g_33_8 (.ZN (n_33_8), .A (n_29_10), .B (n_34_8), .C1 (n_37_5), .C2 (n_43_2) );
AOI211_X1 g_35_7 (.ZN (n_35_7), .A (n_31_9), .B (n_32_9), .C1 (n_35_6), .C2 (n_41_3) );
AOI211_X1 g_34_9 (.ZN (n_34_9), .A (n_33_8), .B (n_31_11), .C1 (n_34_8), .C2 (n_39_4) );
AOI211_X1 g_36_8 (.ZN (n_36_8), .A (n_35_7), .B (n_29_10), .C1 (n_32_9), .C2 (n_37_5) );
AOI211_X1 g_38_7 (.ZN (n_38_7), .A (n_34_9), .B (n_31_9), .C1 (n_31_11), .C2 (n_35_6) );
AOI211_X1 g_37_9 (.ZN (n_37_9), .A (n_36_8), .B (n_33_8), .C1 (n_29_10), .C2 (n_34_8) );
AOI211_X1 g_36_7 (.ZN (n_36_7), .A (n_38_7), .B (n_35_7), .C1 (n_31_9), .C2 (n_32_9) );
AOI211_X1 g_38_6 (.ZN (n_38_6), .A (n_37_9), .B (n_34_9), .C1 (n_33_8), .C2 (n_31_11) );
AOI211_X1 g_40_5 (.ZN (n_40_5), .A (n_36_7), .B (n_36_8), .C1 (n_35_7), .C2 (n_29_10) );
AOI211_X1 g_42_4 (.ZN (n_42_4), .A (n_38_6), .B (n_38_7), .C1 (n_34_9), .C2 (n_31_9) );
AOI211_X1 g_41_6 (.ZN (n_41_6), .A (n_40_5), .B (n_37_9), .C1 (n_36_8), .C2 (n_33_8) );
AOI211_X1 g_39_7 (.ZN (n_39_7), .A (n_42_4), .B (n_36_7), .C1 (n_38_7), .C2 (n_35_7) );
AOI211_X1 g_37_8 (.ZN (n_37_8), .A (n_41_6), .B (n_38_6), .C1 (n_37_9), .C2 (n_34_9) );
AOI211_X1 g_35_9 (.ZN (n_35_9), .A (n_39_7), .B (n_40_5), .C1 (n_36_7), .C2 (n_36_8) );
AOI211_X1 g_33_10 (.ZN (n_33_10), .A (n_37_8), .B (n_42_4), .C1 (n_38_6), .C2 (n_38_7) );
AOI211_X1 g_35_11 (.ZN (n_35_11), .A (n_35_9), .B (n_41_6), .C1 (n_40_5), .C2 (n_37_9) );
AOI211_X1 g_37_10 (.ZN (n_37_10), .A (n_33_10), .B (n_39_7), .C1 (n_42_4), .C2 (n_36_7) );
AOI211_X1 g_39_9 (.ZN (n_39_9), .A (n_35_11), .B (n_37_8), .C1 (n_41_6), .C2 (n_38_6) );
AOI211_X1 g_41_8 (.ZN (n_41_8), .A (n_37_10), .B (n_35_9), .C1 (n_39_7), .C2 (n_40_5) );
AOI211_X1 g_42_6 (.ZN (n_42_6), .A (n_39_9), .B (n_33_10), .C1 (n_37_8), .C2 (n_42_4) );
AOI211_X1 g_43_4 (.ZN (n_43_4), .A (n_41_8), .B (n_35_11), .C1 (n_35_9), .C2 (n_41_6) );
AOI211_X1 g_45_3 (.ZN (n_45_3), .A (n_42_6), .B (n_37_10), .C1 (n_33_10), .C2 (n_39_7) );
AOI211_X1 g_47_2 (.ZN (n_47_2), .A (n_43_4), .B (n_39_9), .C1 (n_35_11), .C2 (n_37_8) );
AOI211_X1 g_49_1 (.ZN (n_49_1), .A (n_45_3), .B (n_41_8), .C1 (n_37_10), .C2 (n_35_9) );
AOI211_X1 g_48_3 (.ZN (n_48_3), .A (n_47_2), .B (n_42_6), .C1 (n_39_9), .C2 (n_33_10) );
AOI211_X1 g_50_2 (.ZN (n_50_2), .A (n_49_1), .B (n_43_4), .C1 (n_41_8), .C2 (n_35_11) );
AOI211_X1 g_52_1 (.ZN (n_52_1), .A (n_48_3), .B (n_45_3), .C1 (n_42_6), .C2 (n_37_10) );
AOI211_X1 g_51_3 (.ZN (n_51_3), .A (n_50_2), .B (n_47_2), .C1 (n_43_4), .C2 (n_39_9) );
AOI211_X1 g_50_1 (.ZN (n_50_1), .A (n_52_1), .B (n_49_1), .C1 (n_45_3), .C2 (n_41_8) );
AOI211_X1 g_48_2 (.ZN (n_48_2), .A (n_51_3), .B (n_48_3), .C1 (n_47_2), .C2 (n_42_6) );
AOI211_X1 g_46_3 (.ZN (n_46_3), .A (n_50_1), .B (n_50_2), .C1 (n_49_1), .C2 (n_43_4) );
AOI211_X1 g_44_4 (.ZN (n_44_4), .A (n_48_2), .B (n_52_1), .C1 (n_48_3), .C2 (n_45_3) );
AOI211_X1 g_42_5 (.ZN (n_42_5), .A (n_46_3), .B (n_51_3), .C1 (n_50_2), .C2 (n_47_2) );
AOI211_X1 g_43_7 (.ZN (n_43_7), .A (n_44_4), .B (n_50_1), .C1 (n_52_1), .C2 (n_49_1) );
AOI211_X1 g_44_5 (.ZN (n_44_5), .A (n_42_5), .B (n_48_2), .C1 (n_51_3), .C2 (n_48_3) );
AOI211_X1 g_46_4 (.ZN (n_46_4), .A (n_43_7), .B (n_46_3), .C1 (n_50_1), .C2 (n_50_2) );
AOI211_X1 g_45_6 (.ZN (n_45_6), .A (n_44_5), .B (n_44_4), .C1 (n_48_2), .C2 (n_52_1) );
AOI211_X1 g_47_5 (.ZN (n_47_5), .A (n_46_4), .B (n_42_5), .C1 (n_46_3), .C2 (n_51_3) );
AOI211_X1 g_49_4 (.ZN (n_49_4), .A (n_45_6), .B (n_43_7), .C1 (n_44_4), .C2 (n_50_1) );
AOI211_X1 g_48_6 (.ZN (n_48_6), .A (n_47_5), .B (n_44_5), .C1 (n_42_5), .C2 (n_48_2) );
AOI211_X1 g_47_4 (.ZN (n_47_4), .A (n_49_4), .B (n_46_4), .C1 (n_43_7), .C2 (n_46_3) );
AOI211_X1 g_49_3 (.ZN (n_49_3), .A (n_48_6), .B (n_45_6), .C1 (n_44_5), .C2 (n_44_4) );
AOI211_X1 g_51_2 (.ZN (n_51_2), .A (n_47_4), .B (n_47_5), .C1 (n_46_4), .C2 (n_42_5) );
AOI211_X1 g_53_1 (.ZN (n_53_1), .A (n_49_3), .B (n_49_4), .C1 (n_45_6), .C2 (n_43_7) );
AOI211_X1 g_52_3 (.ZN (n_52_3), .A (n_51_2), .B (n_48_6), .C1 (n_47_5), .C2 (n_44_5) );
AOI211_X1 g_54_2 (.ZN (n_54_2), .A (n_53_1), .B (n_47_4), .C1 (n_49_4), .C2 (n_46_4) );
AOI211_X1 g_56_1 (.ZN (n_56_1), .A (n_52_3), .B (n_49_3), .C1 (n_48_6), .C2 (n_45_6) );
AOI211_X1 g_55_3 (.ZN (n_55_3), .A (n_54_2), .B (n_51_2), .C1 (n_47_4), .C2 (n_47_5) );
AOI211_X1 g_54_1 (.ZN (n_54_1), .A (n_56_1), .B (n_53_1), .C1 (n_49_3), .C2 (n_49_4) );
AOI211_X1 g_52_2 (.ZN (n_52_2), .A (n_55_3), .B (n_52_3), .C1 (n_51_2), .C2 (n_48_6) );
AOI211_X1 g_50_3 (.ZN (n_50_3), .A (n_54_1), .B (n_54_2), .C1 (n_53_1), .C2 (n_47_4) );
AOI211_X1 g_48_4 (.ZN (n_48_4), .A (n_52_2), .B (n_56_1), .C1 (n_52_3), .C2 (n_49_3) );
AOI211_X1 g_46_5 (.ZN (n_46_5), .A (n_50_3), .B (n_55_3), .C1 (n_54_2), .C2 (n_51_2) );
AOI211_X1 g_44_6 (.ZN (n_44_6), .A (n_48_4), .B (n_54_1), .C1 (n_56_1), .C2 (n_53_1) );
AOI211_X1 g_42_7 (.ZN (n_42_7), .A (n_46_5), .B (n_52_2), .C1 (n_55_3), .C2 (n_52_3) );
AOI211_X1 g_41_5 (.ZN (n_41_5), .A (n_44_6), .B (n_50_3), .C1 (n_54_1), .C2 (n_54_2) );
AOI211_X1 g_40_7 (.ZN (n_40_7), .A (n_42_7), .B (n_48_4), .C1 (n_52_2), .C2 (n_56_1) );
AOI211_X1 g_38_8 (.ZN (n_38_8), .A (n_41_5), .B (n_46_5), .C1 (n_50_3), .C2 (n_55_3) );
AOI211_X1 g_39_6 (.ZN (n_39_6), .A (n_40_7), .B (n_44_6), .C1 (n_48_4), .C2 (n_54_1) );
AOI211_X1 g_37_7 (.ZN (n_37_7), .A (n_38_8), .B (n_42_7), .C1 (n_46_5), .C2 (n_52_2) );
AOI211_X1 g_35_8 (.ZN (n_35_8), .A (n_39_6), .B (n_41_5), .C1 (n_44_6), .C2 (n_50_3) );
AOI211_X1 g_33_9 (.ZN (n_33_9), .A (n_37_7), .B (n_40_7), .C1 (n_42_7), .C2 (n_48_4) );
AOI211_X1 g_31_10 (.ZN (n_31_10), .A (n_35_8), .B (n_38_8), .C1 (n_41_5), .C2 (n_46_5) );
AOI211_X1 g_29_11 (.ZN (n_29_11), .A (n_33_9), .B (n_39_6), .C1 (n_40_7), .C2 (n_44_6) );
AOI211_X1 g_27_12 (.ZN (n_27_12), .A (n_31_10), .B (n_37_7), .C1 (n_38_8), .C2 (n_42_7) );
AOI211_X1 g_28_10 (.ZN (n_28_10), .A (n_29_11), .B (n_35_8), .C1 (n_39_6), .C2 (n_41_5) );
AOI211_X1 g_26_11 (.ZN (n_26_11), .A (n_27_12), .B (n_33_9), .C1 (n_37_7), .C2 (n_40_7) );
AOI211_X1 g_24_12 (.ZN (n_24_12), .A (n_28_10), .B (n_31_10), .C1 (n_35_8), .C2 (n_38_8) );
AOI211_X1 g_22_13 (.ZN (n_22_13), .A (n_26_11), .B (n_29_11), .C1 (n_33_9), .C2 (n_39_6) );
AOI211_X1 g_20_14 (.ZN (n_20_14), .A (n_24_12), .B (n_27_12), .C1 (n_31_10), .C2 (n_37_7) );
AOI211_X1 g_18_15 (.ZN (n_18_15), .A (n_22_13), .B (n_28_10), .C1 (n_29_11), .C2 (n_35_8) );
AOI211_X1 g_16_14 (.ZN (n_16_14), .A (n_20_14), .B (n_26_11), .C1 (n_27_12), .C2 (n_33_9) );
AOI211_X1 g_14_13 (.ZN (n_14_13), .A (n_18_15), .B (n_24_12), .C1 (n_28_10), .C2 (n_31_10) );
AOI211_X1 g_12_12 (.ZN (n_12_12), .A (n_16_14), .B (n_22_13), .C1 (n_26_11), .C2 (n_29_11) );
AOI211_X1 g_13_14 (.ZN (n_13_14), .A (n_14_13), .B (n_20_14), .C1 (n_24_12), .C2 (n_27_12) );
AOI211_X1 g_15_15 (.ZN (n_15_15), .A (n_12_12), .B (n_18_15), .C1 (n_22_13), .C2 (n_28_10) );
AOI211_X1 g_17_16 (.ZN (n_17_16), .A (n_13_14), .B (n_16_14), .C1 (n_20_14), .C2 (n_26_11) );
AOI211_X1 g_19_17 (.ZN (n_19_17), .A (n_15_15), .B (n_14_13), .C1 (n_18_15), .C2 (n_24_12) );
AOI211_X1 g_21_16 (.ZN (n_21_16), .A (n_17_16), .B (n_12_12), .C1 (n_16_14), .C2 (n_22_13) );
AOI211_X1 g_23_15 (.ZN (n_23_15), .A (n_19_17), .B (n_13_14), .C1 (n_14_13), .C2 (n_20_14) );
AOI211_X1 g_21_14 (.ZN (n_21_14), .A (n_21_16), .B (n_15_15), .C1 (n_12_12), .C2 (n_18_15) );
AOI211_X1 g_23_13 (.ZN (n_23_13), .A (n_23_15), .B (n_17_16), .C1 (n_13_14), .C2 (n_16_14) );
AOI211_X1 g_25_12 (.ZN (n_25_12), .A (n_21_14), .B (n_19_17), .C1 (n_15_15), .C2 (n_14_13) );
AOI211_X1 g_27_11 (.ZN (n_27_11), .A (n_23_13), .B (n_21_16), .C1 (n_17_16), .C2 (n_12_12) );
AOI211_X1 g_29_12 (.ZN (n_29_12), .A (n_25_12), .B (n_23_15), .C1 (n_19_17), .C2 (n_13_14) );
AOI211_X1 g_27_13 (.ZN (n_27_13), .A (n_27_11), .B (n_21_14), .C1 (n_21_16), .C2 (n_15_15) );
AOI211_X1 g_25_14 (.ZN (n_25_14), .A (n_29_12), .B (n_23_13), .C1 (n_23_15), .C2 (n_17_16) );
AOI211_X1 g_24_16 (.ZN (n_24_16), .A (n_27_13), .B (n_25_12), .C1 (n_21_14), .C2 (n_19_17) );
AOI211_X1 g_23_14 (.ZN (n_23_14), .A (n_25_14), .B (n_27_11), .C1 (n_23_13), .C2 (n_21_16) );
AOI211_X1 g_25_13 (.ZN (n_25_13), .A (n_24_16), .B (n_29_12), .C1 (n_25_12), .C2 (n_23_15) );
AOI211_X1 g_24_15 (.ZN (n_24_15), .A (n_23_14), .B (n_27_13), .C1 (n_27_11), .C2 (n_21_14) );
AOI211_X1 g_26_14 (.ZN (n_26_14), .A (n_25_13), .B (n_25_14), .C1 (n_29_12), .C2 (n_23_13) );
AOI211_X1 g_28_13 (.ZN (n_28_13), .A (n_24_15), .B (n_24_16), .C1 (n_27_13), .C2 (n_25_12) );
AOI211_X1 g_30_12 (.ZN (n_30_12), .A (n_26_14), .B (n_23_14), .C1 (n_25_14), .C2 (n_27_11) );
AOI211_X1 g_32_11 (.ZN (n_32_11), .A (n_28_13), .B (n_25_13), .C1 (n_24_16), .C2 (n_29_12) );
AOI211_X1 g_34_10 (.ZN (n_34_10), .A (n_30_12), .B (n_24_15), .C1 (n_23_14), .C2 (n_27_13) );
AOI211_X1 g_36_9 (.ZN (n_36_9), .A (n_32_11), .B (n_26_14), .C1 (n_25_13), .C2 (n_25_14) );
AOI211_X1 g_38_10 (.ZN (n_38_10), .A (n_34_10), .B (n_28_13), .C1 (n_24_15), .C2 (n_24_16) );
AOI211_X1 g_39_8 (.ZN (n_39_8), .A (n_36_9), .B (n_30_12), .C1 (n_26_14), .C2 (n_23_14) );
AOI211_X1 g_41_7 (.ZN (n_41_7), .A (n_38_10), .B (n_32_11), .C1 (n_28_13), .C2 (n_25_13) );
AOI211_X1 g_43_6 (.ZN (n_43_6), .A (n_39_8), .B (n_34_10), .C1 (n_30_12), .C2 (n_24_15) );
AOI211_X1 g_45_5 (.ZN (n_45_5), .A (n_41_7), .B (n_36_9), .C1 (n_32_11), .C2 (n_26_14) );
AOI211_X1 g_46_7 (.ZN (n_46_7), .A (n_43_6), .B (n_38_10), .C1 (n_34_10), .C2 (n_28_13) );
AOI211_X1 g_44_8 (.ZN (n_44_8), .A (n_45_5), .B (n_39_8), .C1 (n_36_9), .C2 (n_30_12) );
AOI211_X1 g_42_9 (.ZN (n_42_9), .A (n_46_7), .B (n_41_7), .C1 (n_38_10), .C2 (n_32_11) );
AOI211_X1 g_40_8 (.ZN (n_40_8), .A (n_44_8), .B (n_43_6), .C1 (n_39_8), .C2 (n_34_10) );
AOI211_X1 g_38_9 (.ZN (n_38_9), .A (n_42_9), .B (n_45_5), .C1 (n_41_7), .C2 (n_36_9) );
AOI211_X1 g_36_10 (.ZN (n_36_10), .A (n_40_8), .B (n_46_7), .C1 (n_43_6), .C2 (n_38_10) );
AOI211_X1 g_34_11 (.ZN (n_34_11), .A (n_38_9), .B (n_44_8), .C1 (n_45_5), .C2 (n_39_8) );
AOI211_X1 g_32_10 (.ZN (n_32_10), .A (n_36_10), .B (n_42_9), .C1 (n_46_7), .C2 (n_41_7) );
AOI211_X1 g_30_11 (.ZN (n_30_11), .A (n_34_11), .B (n_40_8), .C1 (n_44_8), .C2 (n_43_6) );
AOI211_X1 g_28_12 (.ZN (n_28_12), .A (n_32_10), .B (n_38_9), .C1 (n_42_9), .C2 (n_45_5) );
AOI211_X1 g_26_13 (.ZN (n_26_13), .A (n_30_11), .B (n_36_10), .C1 (n_40_8), .C2 (n_46_7) );
AOI211_X1 g_24_14 (.ZN (n_24_14), .A (n_28_12), .B (n_34_11), .C1 (n_38_9), .C2 (n_44_8) );
AOI211_X1 g_22_15 (.ZN (n_22_15), .A (n_26_13), .B (n_32_10), .C1 (n_36_10), .C2 (n_42_9) );
AOI211_X1 g_20_16 (.ZN (n_20_16), .A (n_24_14), .B (n_30_11), .C1 (n_34_11), .C2 (n_40_8) );
AOI211_X1 g_22_17 (.ZN (n_22_17), .A (n_22_15), .B (n_28_12), .C1 (n_32_10), .C2 (n_38_9) );
AOI211_X1 g_21_15 (.ZN (n_21_15), .A (n_20_16), .B (n_26_13), .C1 (n_30_11), .C2 (n_36_10) );
AOI211_X1 g_19_16 (.ZN (n_19_16), .A (n_22_17), .B (n_24_14), .C1 (n_28_12), .C2 (n_34_11) );
AOI211_X1 g_17_15 (.ZN (n_17_15), .A (n_21_15), .B (n_22_15), .C1 (n_26_13), .C2 (n_32_10) );
AOI211_X1 g_16_17 (.ZN (n_16_17), .A (n_19_16), .B (n_20_16), .C1 (n_24_14), .C2 (n_30_11) );
AOI211_X1 g_18_18 (.ZN (n_18_18), .A (n_17_15), .B (n_22_17), .C1 (n_22_15), .C2 (n_28_12) );
AOI211_X1 g_20_17 (.ZN (n_20_17), .A (n_16_17), .B (n_21_15), .C1 (n_20_16), .C2 (n_26_13) );
AOI211_X1 g_22_16 (.ZN (n_22_16), .A (n_18_18), .B (n_19_16), .C1 (n_22_17), .C2 (n_24_14) );
AOI211_X1 g_21_18 (.ZN (n_21_18), .A (n_20_17), .B (n_17_15), .C1 (n_21_15), .C2 (n_22_15) );
AOI211_X1 g_23_17 (.ZN (n_23_17), .A (n_22_16), .B (n_16_17), .C1 (n_19_16), .C2 (n_20_16) );
AOI211_X1 g_25_16 (.ZN (n_25_16), .A (n_21_18), .B (n_18_18), .C1 (n_17_15), .C2 (n_22_17) );
AOI211_X1 g_27_15 (.ZN (n_27_15), .A (n_23_17), .B (n_20_17), .C1 (n_16_17), .C2 (n_21_15) );
AOI211_X1 g_29_14 (.ZN (n_29_14), .A (n_25_16), .B (n_22_16), .C1 (n_18_18), .C2 (n_19_16) );
AOI211_X1 g_31_13 (.ZN (n_31_13), .A (n_27_15), .B (n_21_18), .C1 (n_20_17), .C2 (n_17_15) );
AOI211_X1 g_33_12 (.ZN (n_33_12), .A (n_29_14), .B (n_23_17), .C1 (n_22_16), .C2 (n_16_17) );
AOI211_X1 g_35_13 (.ZN (n_35_13), .A (n_31_13), .B (n_25_16), .C1 (n_21_18), .C2 (n_18_18) );
AOI211_X1 g_36_11 (.ZN (n_36_11), .A (n_33_12), .B (n_27_15), .C1 (n_23_17), .C2 (n_20_17) );
AOI211_X1 g_34_12 (.ZN (n_34_12), .A (n_35_13), .B (n_29_14), .C1 (n_25_16), .C2 (n_22_16) );
AOI211_X1 g_35_10 (.ZN (n_35_10), .A (n_36_11), .B (n_31_13), .C1 (n_27_15), .C2 (n_21_18) );
AOI211_X1 g_33_11 (.ZN (n_33_11), .A (n_34_12), .B (n_33_12), .C1 (n_29_14), .C2 (n_23_17) );
AOI211_X1 g_31_12 (.ZN (n_31_12), .A (n_35_10), .B (n_35_13), .C1 (n_31_13), .C2 (n_25_16) );
AOI211_X1 g_29_13 (.ZN (n_29_13), .A (n_33_11), .B (n_36_11), .C1 (n_33_12), .C2 (n_27_15) );
AOI211_X1 g_27_14 (.ZN (n_27_14), .A (n_31_12), .B (n_34_12), .C1 (n_35_13), .C2 (n_29_14) );
AOI211_X1 g_25_15 (.ZN (n_25_15), .A (n_29_13), .B (n_35_10), .C1 (n_36_11), .C2 (n_31_13) );
AOI211_X1 g_23_16 (.ZN (n_23_16), .A (n_27_14), .B (n_33_11), .C1 (n_34_12), .C2 (n_33_12) );
AOI211_X1 g_21_17 (.ZN (n_21_17), .A (n_25_15), .B (n_31_12), .C1 (n_35_10), .C2 (n_35_13) );
AOI211_X1 g_19_18 (.ZN (n_19_18), .A (n_23_16), .B (n_29_13), .C1 (n_33_11), .C2 (n_36_11) );
AOI211_X1 g_17_17 (.ZN (n_17_17), .A (n_21_17), .B (n_27_14), .C1 (n_31_12), .C2 (n_34_12) );
AOI211_X1 g_15_16 (.ZN (n_15_16), .A (n_19_18), .B (n_25_15), .C1 (n_29_13), .C2 (n_35_10) );
AOI211_X1 g_13_15 (.ZN (n_13_15), .A (n_17_17), .B (n_23_16), .C1 (n_27_14), .C2 (n_33_11) );
AOI211_X1 g_11_14 (.ZN (n_11_14), .A (n_15_16), .B (n_21_17), .C1 (n_25_15), .C2 (n_31_12) );
AOI211_X1 g_9_15 (.ZN (n_9_15), .A (n_13_15), .B (n_19_18), .C1 (n_23_16), .C2 (n_29_13) );
AOI211_X1 g_10_13 (.ZN (n_10_13), .A (n_11_14), .B (n_17_17), .C1 (n_21_17), .C2 (n_27_14) );
AOI211_X1 g_8_14 (.ZN (n_8_14), .A (n_9_15), .B (n_15_16), .C1 (n_19_18), .C2 (n_25_15) );
AOI211_X1 g_10_15 (.ZN (n_10_15), .A (n_10_13), .B (n_13_15), .C1 (n_17_17), .C2 (n_23_16) );
AOI211_X1 g_12_14 (.ZN (n_12_14), .A (n_8_14), .B (n_11_14), .C1 (n_15_16), .C2 (n_21_17) );
AOI211_X1 g_11_16 (.ZN (n_11_16), .A (n_10_15), .B (n_9_15), .C1 (n_13_15), .C2 (n_19_18) );
AOI211_X1 g_13_17 (.ZN (n_13_17), .A (n_12_14), .B (n_10_13), .C1 (n_11_14), .C2 (n_17_17) );
AOI211_X1 g_14_15 (.ZN (n_14_15), .A (n_11_16), .B (n_8_14), .C1 (n_9_15), .C2 (n_15_16) );
AOI211_X1 g_12_16 (.ZN (n_12_16), .A (n_13_17), .B (n_10_15), .C1 (n_10_13), .C2 (n_13_15) );
AOI211_X1 g_14_17 (.ZN (n_14_17), .A (n_14_15), .B (n_12_14), .C1 (n_8_14), .C2 (n_11_14) );
AOI211_X1 g_16_16 (.ZN (n_16_16), .A (n_12_16), .B (n_11_16), .C1 (n_10_15), .C2 (n_9_15) );
AOI211_X1 g_15_18 (.ZN (n_15_18), .A (n_14_17), .B (n_13_17), .C1 (n_12_14), .C2 (n_10_13) );
AOI211_X1 g_17_19 (.ZN (n_17_19), .A (n_16_16), .B (n_14_15), .C1 (n_11_16), .C2 (n_8_14) );
AOI211_X1 g_18_17 (.ZN (n_18_17), .A (n_15_18), .B (n_12_16), .C1 (n_13_17), .C2 (n_10_15) );
AOI211_X1 g_16_18 (.ZN (n_16_18), .A (n_17_19), .B (n_14_17), .C1 (n_14_15), .C2 (n_12_14) );
AOI211_X1 g_18_19 (.ZN (n_18_19), .A (n_18_17), .B (n_16_16), .C1 (n_12_16), .C2 (n_11_16) );
AOI211_X1 g_20_18 (.ZN (n_20_18), .A (n_16_18), .B (n_15_18), .C1 (n_14_17), .C2 (n_13_17) );
AOI211_X1 g_19_20 (.ZN (n_19_20), .A (n_18_19), .B (n_17_19), .C1 (n_16_16), .C2 (n_14_15) );
AOI211_X1 g_21_19 (.ZN (n_21_19), .A (n_20_18), .B (n_18_17), .C1 (n_15_18), .C2 (n_12_16) );
AOI211_X1 g_23_18 (.ZN (n_23_18), .A (n_19_20), .B (n_16_18), .C1 (n_17_19), .C2 (n_14_17) );
AOI211_X1 g_25_17 (.ZN (n_25_17), .A (n_21_19), .B (n_18_19), .C1 (n_18_17), .C2 (n_16_16) );
AOI211_X1 g_26_15 (.ZN (n_26_15), .A (n_23_18), .B (n_20_18), .C1 (n_16_18), .C2 (n_15_18) );
AOI211_X1 g_28_14 (.ZN (n_28_14), .A (n_25_17), .B (n_19_20), .C1 (n_18_19), .C2 (n_17_19) );
AOI211_X1 g_30_13 (.ZN (n_30_13), .A (n_26_15), .B (n_21_19), .C1 (n_20_18), .C2 (n_18_17) );
AOI211_X1 g_32_12 (.ZN (n_32_12), .A (n_28_14), .B (n_23_18), .C1 (n_19_20), .C2 (n_16_18) );
AOI211_X1 g_33_14 (.ZN (n_33_14), .A (n_30_13), .B (n_25_17), .C1 (n_21_19), .C2 (n_18_19) );
AOI211_X1 g_31_15 (.ZN (n_31_15), .A (n_32_12), .B (n_26_15), .C1 (n_23_18), .C2 (n_20_18) );
AOI211_X1 g_32_13 (.ZN (n_32_13), .A (n_33_14), .B (n_28_14), .C1 (n_25_17), .C2 (n_19_20) );
AOI211_X1 g_30_14 (.ZN (n_30_14), .A (n_31_15), .B (n_30_13), .C1 (n_26_15), .C2 (n_21_19) );
AOI211_X1 g_28_15 (.ZN (n_28_15), .A (n_32_13), .B (n_32_12), .C1 (n_28_14), .C2 (n_23_18) );
AOI211_X1 g_26_16 (.ZN (n_26_16), .A (n_30_14), .B (n_33_14), .C1 (n_30_13), .C2 (n_25_17) );
AOI211_X1 g_24_17 (.ZN (n_24_17), .A (n_28_15), .B (n_31_15), .C1 (n_32_12), .C2 (n_26_15) );
AOI211_X1 g_22_18 (.ZN (n_22_18), .A (n_26_16), .B (n_32_13), .C1 (n_33_14), .C2 (n_28_14) );
AOI211_X1 g_20_19 (.ZN (n_20_19), .A (n_24_17), .B (n_30_14), .C1 (n_31_15), .C2 (n_30_13) );
AOI211_X1 g_22_20 (.ZN (n_22_20), .A (n_22_18), .B (n_28_15), .C1 (n_32_13), .C2 (n_32_12) );
AOI211_X1 g_24_19 (.ZN (n_24_19), .A (n_20_19), .B (n_26_16), .C1 (n_30_14), .C2 (n_33_14) );
AOI211_X1 g_26_18 (.ZN (n_26_18), .A (n_22_20), .B (n_24_17), .C1 (n_28_15), .C2 (n_31_15) );
AOI211_X1 g_27_16 (.ZN (n_27_16), .A (n_24_19), .B (n_22_18), .C1 (n_26_16), .C2 (n_32_13) );
AOI211_X1 g_29_15 (.ZN (n_29_15), .A (n_26_18), .B (n_20_19), .C1 (n_24_17), .C2 (n_30_14) );
AOI211_X1 g_31_14 (.ZN (n_31_14), .A (n_27_16), .B (n_22_20), .C1 (n_22_18), .C2 (n_28_15) );
AOI211_X1 g_33_13 (.ZN (n_33_13), .A (n_29_15), .B (n_24_19), .C1 (n_20_19), .C2 (n_26_16) );
AOI211_X1 g_35_12 (.ZN (n_35_12), .A (n_31_14), .B (n_26_18), .C1 (n_22_20), .C2 (n_24_17) );
AOI211_X1 g_37_11 (.ZN (n_37_11), .A (n_33_13), .B (n_27_16), .C1 (n_24_19), .C2 (n_22_18) );
AOI211_X1 g_39_10 (.ZN (n_39_10), .A (n_35_12), .B (n_29_15), .C1 (n_26_18), .C2 (n_20_19) );
AOI211_X1 g_41_9 (.ZN (n_41_9), .A (n_37_11), .B (n_31_14), .C1 (n_27_16), .C2 (n_22_20) );
AOI211_X1 g_43_8 (.ZN (n_43_8), .A (n_39_10), .B (n_33_13), .C1 (n_29_15), .C2 (n_24_19) );
AOI211_X1 g_45_7 (.ZN (n_45_7), .A (n_41_9), .B (n_35_12), .C1 (n_31_14), .C2 (n_26_18) );
AOI211_X1 g_47_6 (.ZN (n_47_6), .A (n_43_8), .B (n_37_11), .C1 (n_33_13), .C2 (n_27_16) );
AOI211_X1 g_49_5 (.ZN (n_49_5), .A (n_45_7), .B (n_39_10), .C1 (n_35_12), .C2 (n_29_15) );
AOI211_X1 g_51_4 (.ZN (n_51_4), .A (n_47_6), .B (n_41_9), .C1 (n_37_11), .C2 (n_31_14) );
AOI211_X1 g_53_3 (.ZN (n_53_3), .A (n_49_5), .B (n_43_8), .C1 (n_39_10), .C2 (n_33_13) );
AOI211_X1 g_55_2 (.ZN (n_55_2), .A (n_51_4), .B (n_45_7), .C1 (n_41_9), .C2 (n_35_12) );
AOI211_X1 g_57_1 (.ZN (n_57_1), .A (n_53_3), .B (n_47_6), .C1 (n_43_8), .C2 (n_37_11) );
AOI211_X1 g_56_3 (.ZN (n_56_3), .A (n_55_2), .B (n_49_5), .C1 (n_45_7), .C2 (n_39_10) );
AOI211_X1 g_58_2 (.ZN (n_58_2), .A (n_57_1), .B (n_51_4), .C1 (n_47_6), .C2 (n_41_9) );
AOI211_X1 g_60_1 (.ZN (n_60_1), .A (n_56_3), .B (n_53_3), .C1 (n_49_5), .C2 (n_43_8) );
AOI211_X1 g_59_3 (.ZN (n_59_3), .A (n_58_2), .B (n_55_2), .C1 (n_51_4), .C2 (n_45_7) );
AOI211_X1 g_58_1 (.ZN (n_58_1), .A (n_60_1), .B (n_57_1), .C1 (n_53_3), .C2 (n_47_6) );
AOI211_X1 g_56_2 (.ZN (n_56_2), .A (n_59_3), .B (n_56_3), .C1 (n_55_2), .C2 (n_49_5) );
AOI211_X1 g_54_3 (.ZN (n_54_3), .A (n_58_1), .B (n_58_2), .C1 (n_57_1), .C2 (n_51_4) );
AOI211_X1 g_52_4 (.ZN (n_52_4), .A (n_56_2), .B (n_60_1), .C1 (n_56_3), .C2 (n_53_3) );
AOI211_X1 g_50_5 (.ZN (n_50_5), .A (n_54_3), .B (n_59_3), .C1 (n_58_2), .C2 (n_55_2) );
AOI211_X1 g_49_7 (.ZN (n_49_7), .A (n_52_4), .B (n_58_1), .C1 (n_60_1), .C2 (n_57_1) );
AOI211_X1 g_48_5 (.ZN (n_48_5), .A (n_50_5), .B (n_56_2), .C1 (n_59_3), .C2 (n_56_3) );
AOI211_X1 g_50_4 (.ZN (n_50_4), .A (n_49_7), .B (n_54_3), .C1 (n_58_1), .C2 (n_58_2) );
AOI211_X1 g_51_6 (.ZN (n_51_6), .A (n_48_5), .B (n_52_4), .C1 (n_56_2), .C2 (n_60_1) );
AOI211_X1 g_53_5 (.ZN (n_53_5), .A (n_50_4), .B (n_50_5), .C1 (n_54_3), .C2 (n_59_3) );
AOI211_X1 g_55_4 (.ZN (n_55_4), .A (n_51_6), .B (n_49_7), .C1 (n_52_4), .C2 (n_58_1) );
AOI211_X1 g_57_3 (.ZN (n_57_3), .A (n_53_5), .B (n_48_5), .C1 (n_50_5), .C2 (n_56_2) );
AOI211_X1 g_59_2 (.ZN (n_59_2), .A (n_55_4), .B (n_50_4), .C1 (n_49_7), .C2 (n_54_3) );
AOI211_X1 g_61_1 (.ZN (n_61_1), .A (n_57_3), .B (n_51_6), .C1 (n_48_5), .C2 (n_52_4) );
AOI211_X1 g_60_3 (.ZN (n_60_3), .A (n_59_2), .B (n_53_5), .C1 (n_50_4), .C2 (n_50_5) );
AOI211_X1 g_62_2 (.ZN (n_62_2), .A (n_61_1), .B (n_55_4), .C1 (n_51_6), .C2 (n_49_7) );
AOI211_X1 g_64_1 (.ZN (n_64_1), .A (n_60_3), .B (n_57_3), .C1 (n_53_5), .C2 (n_48_5) );
AOI211_X1 g_63_3 (.ZN (n_63_3), .A (n_62_2), .B (n_59_2), .C1 (n_55_4), .C2 (n_50_4) );
AOI211_X1 g_62_1 (.ZN (n_62_1), .A (n_64_1), .B (n_61_1), .C1 (n_57_3), .C2 (n_51_6) );
AOI211_X1 g_60_2 (.ZN (n_60_2), .A (n_63_3), .B (n_60_3), .C1 (n_59_2), .C2 (n_53_5) );
AOI211_X1 g_58_3 (.ZN (n_58_3), .A (n_62_1), .B (n_62_2), .C1 (n_61_1), .C2 (n_55_4) );
AOI211_X1 g_56_4 (.ZN (n_56_4), .A (n_60_2), .B (n_64_1), .C1 (n_60_3), .C2 (n_57_3) );
AOI211_X1 g_54_5 (.ZN (n_54_5), .A (n_58_3), .B (n_63_3), .C1 (n_62_2), .C2 (n_59_2) );
AOI211_X1 g_52_6 (.ZN (n_52_6), .A (n_56_4), .B (n_62_1), .C1 (n_64_1), .C2 (n_61_1) );
AOI211_X1 g_53_4 (.ZN (n_53_4), .A (n_54_5), .B (n_60_2), .C1 (n_63_3), .C2 (n_60_3) );
AOI211_X1 g_51_5 (.ZN (n_51_5), .A (n_52_6), .B (n_58_3), .C1 (n_62_1), .C2 (n_62_2) );
AOI211_X1 g_49_6 (.ZN (n_49_6), .A (n_53_4), .B (n_56_4), .C1 (n_60_2), .C2 (n_64_1) );
AOI211_X1 g_47_7 (.ZN (n_47_7), .A (n_51_5), .B (n_54_5), .C1 (n_58_3), .C2 (n_63_3) );
AOI211_X1 g_45_8 (.ZN (n_45_8), .A (n_49_6), .B (n_52_6), .C1 (n_56_4), .C2 (n_62_1) );
AOI211_X1 g_46_6 (.ZN (n_46_6), .A (n_47_7), .B (n_53_4), .C1 (n_54_5), .C2 (n_60_2) );
AOI211_X1 g_44_7 (.ZN (n_44_7), .A (n_45_8), .B (n_51_5), .C1 (n_52_6), .C2 (n_58_3) );
AOI211_X1 g_42_8 (.ZN (n_42_8), .A (n_46_6), .B (n_49_6), .C1 (n_53_4), .C2 (n_56_4) );
AOI211_X1 g_40_9 (.ZN (n_40_9), .A (n_44_7), .B (n_47_7), .C1 (n_51_5), .C2 (n_54_5) );
AOI211_X1 g_39_11 (.ZN (n_39_11), .A (n_42_8), .B (n_45_8), .C1 (n_49_6), .C2 (n_52_6) );
AOI211_X1 g_37_12 (.ZN (n_37_12), .A (n_40_9), .B (n_46_6), .C1 (n_47_7), .C2 (n_53_4) );
AOI211_X1 g_36_14 (.ZN (n_36_14), .A (n_39_11), .B (n_44_7), .C1 (n_45_8), .C2 (n_51_5) );
AOI211_X1 g_34_13 (.ZN (n_34_13), .A (n_37_12), .B (n_42_8), .C1 (n_46_6), .C2 (n_49_6) );
AOI211_X1 g_36_12 (.ZN (n_36_12), .A (n_36_14), .B (n_40_9), .C1 (n_44_7), .C2 (n_47_7) );
AOI211_X1 g_38_11 (.ZN (n_38_11), .A (n_34_13), .B (n_39_11), .C1 (n_42_8), .C2 (n_45_8) );
AOI211_X1 g_40_10 (.ZN (n_40_10), .A (n_36_12), .B (n_37_12), .C1 (n_40_9), .C2 (n_46_6) );
AOI211_X1 g_39_12 (.ZN (n_39_12), .A (n_38_11), .B (n_36_14), .C1 (n_39_11), .C2 (n_44_7) );
AOI211_X1 g_41_11 (.ZN (n_41_11), .A (n_40_10), .B (n_34_13), .C1 (n_37_12), .C2 (n_42_8) );
AOI211_X1 g_43_10 (.ZN (n_43_10), .A (n_39_12), .B (n_36_12), .C1 (n_36_14), .C2 (n_40_9) );
AOI211_X1 g_45_9 (.ZN (n_45_9), .A (n_41_11), .B (n_38_11), .C1 (n_34_13), .C2 (n_39_11) );
AOI211_X1 g_47_8 (.ZN (n_47_8), .A (n_43_10), .B (n_40_10), .C1 (n_36_12), .C2 (n_37_12) );
AOI211_X1 g_46_10 (.ZN (n_46_10), .A (n_45_9), .B (n_39_12), .C1 (n_38_11), .C2 (n_36_14) );
AOI211_X1 g_44_9 (.ZN (n_44_9), .A (n_47_8), .B (n_41_11), .C1 (n_40_10), .C2 (n_34_13) );
AOI211_X1 g_46_8 (.ZN (n_46_8), .A (n_46_10), .B (n_43_10), .C1 (n_39_12), .C2 (n_36_12) );
AOI211_X1 g_48_7 (.ZN (n_48_7), .A (n_44_9), .B (n_45_9), .C1 (n_41_11), .C2 (n_38_11) );
AOI211_X1 g_50_6 (.ZN (n_50_6), .A (n_46_8), .B (n_47_8), .C1 (n_43_10), .C2 (n_40_10) );
AOI211_X1 g_52_5 (.ZN (n_52_5), .A (n_48_7), .B (n_46_10), .C1 (n_45_9), .C2 (n_39_12) );
AOI211_X1 g_54_4 (.ZN (n_54_4), .A (n_50_6), .B (n_44_9), .C1 (n_47_8), .C2 (n_41_11) );
AOI211_X1 g_53_6 (.ZN (n_53_6), .A (n_52_5), .B (n_46_8), .C1 (n_46_10), .C2 (n_43_10) );
AOI211_X1 g_55_5 (.ZN (n_55_5), .A (n_54_4), .B (n_48_7), .C1 (n_44_9), .C2 (n_45_9) );
AOI211_X1 g_57_4 (.ZN (n_57_4), .A (n_53_6), .B (n_50_6), .C1 (n_46_8), .C2 (n_47_8) );
AOI211_X1 g_56_6 (.ZN (n_56_6), .A (n_55_5), .B (n_52_5), .C1 (n_48_7), .C2 (n_46_10) );
AOI211_X1 g_58_5 (.ZN (n_58_5), .A (n_57_4), .B (n_54_4), .C1 (n_50_6), .C2 (n_44_9) );
AOI211_X1 g_60_4 (.ZN (n_60_4), .A (n_56_6), .B (n_53_6), .C1 (n_52_5), .C2 (n_46_8) );
AOI211_X1 g_62_3 (.ZN (n_62_3), .A (n_58_5), .B (n_55_5), .C1 (n_54_4), .C2 (n_48_7) );
AOI211_X1 g_64_2 (.ZN (n_64_2), .A (n_60_4), .B (n_57_4), .C1 (n_53_6), .C2 (n_50_6) );
AOI211_X1 g_66_1 (.ZN (n_66_1), .A (n_62_3), .B (n_56_6), .C1 (n_55_5), .C2 (n_52_5) );
AOI211_X1 g_67_3 (.ZN (n_67_3), .A (n_64_2), .B (n_58_5), .C1 (n_57_4), .C2 (n_54_4) );
AOI211_X1 g_68_1 (.ZN (n_68_1), .A (n_66_1), .B (n_60_4), .C1 (n_56_6), .C2 (n_53_6) );
AOI211_X1 g_66_2 (.ZN (n_66_2), .A (n_67_3), .B (n_62_3), .C1 (n_58_5), .C2 (n_55_5) );
AOI211_X1 g_65_4 (.ZN (n_65_4), .A (n_68_1), .B (n_64_2), .C1 (n_60_4), .C2 (n_57_4) );
AOI211_X1 g_63_5 (.ZN (n_63_5), .A (n_66_2), .B (n_66_1), .C1 (n_62_3), .C2 (n_56_6) );
AOI211_X1 g_61_4 (.ZN (n_61_4), .A (n_65_4), .B (n_67_3), .C1 (n_64_2), .C2 (n_58_5) );
AOI211_X1 g_59_5 (.ZN (n_59_5), .A (n_63_5), .B (n_68_1), .C1 (n_66_1), .C2 (n_60_4) );
AOI211_X1 g_57_6 (.ZN (n_57_6), .A (n_61_4), .B (n_66_2), .C1 (n_67_3), .C2 (n_62_3) );
AOI211_X1 g_58_4 (.ZN (n_58_4), .A (n_59_5), .B (n_65_4), .C1 (n_68_1), .C2 (n_64_2) );
AOI211_X1 g_56_5 (.ZN (n_56_5), .A (n_57_6), .B (n_63_5), .C1 (n_66_2), .C2 (n_66_1) );
AOI211_X1 g_54_6 (.ZN (n_54_6), .A (n_58_4), .B (n_61_4), .C1 (n_65_4), .C2 (n_67_3) );
AOI211_X1 g_52_7 (.ZN (n_52_7), .A (n_56_5), .B (n_59_5), .C1 (n_63_5), .C2 (n_68_1) );
AOI211_X1 g_50_8 (.ZN (n_50_8), .A (n_54_6), .B (n_57_6), .C1 (n_61_4), .C2 (n_66_2) );
AOI211_X1 g_48_9 (.ZN (n_48_9), .A (n_52_7), .B (n_58_4), .C1 (n_59_5), .C2 (n_65_4) );
AOI211_X1 g_47_11 (.ZN (n_47_11), .A (n_50_8), .B (n_56_5), .C1 (n_57_6), .C2 (n_63_5) );
AOI211_X1 g_46_9 (.ZN (n_46_9), .A (n_48_9), .B (n_54_6), .C1 (n_58_4), .C2 (n_61_4) );
AOI211_X1 g_48_8 (.ZN (n_48_8), .A (n_47_11), .B (n_52_7), .C1 (n_56_5), .C2 (n_59_5) );
AOI211_X1 g_50_7 (.ZN (n_50_7), .A (n_46_9), .B (n_50_8), .C1 (n_54_6), .C2 (n_57_6) );
AOI211_X1 g_49_9 (.ZN (n_49_9), .A (n_48_8), .B (n_48_9), .C1 (n_52_7), .C2 (n_58_4) );
AOI211_X1 g_51_8 (.ZN (n_51_8), .A (n_50_7), .B (n_47_11), .C1 (n_50_8), .C2 (n_56_5) );
AOI211_X1 g_53_7 (.ZN (n_53_7), .A (n_49_9), .B (n_46_9), .C1 (n_48_9), .C2 (n_54_6) );
AOI211_X1 g_55_6 (.ZN (n_55_6), .A (n_51_8), .B (n_48_8), .C1 (n_47_11), .C2 (n_52_7) );
AOI211_X1 g_57_5 (.ZN (n_57_5), .A (n_53_7), .B (n_50_7), .C1 (n_46_9), .C2 (n_50_8) );
AOI211_X1 g_59_4 (.ZN (n_59_4), .A (n_55_6), .B (n_49_9), .C1 (n_48_8), .C2 (n_48_9) );
AOI211_X1 g_61_3 (.ZN (n_61_3), .A (n_57_5), .B (n_51_8), .C1 (n_50_7), .C2 (n_47_11) );
AOI211_X1 g_63_2 (.ZN (n_63_2), .A (n_59_4), .B (n_53_7), .C1 (n_49_9), .C2 (n_46_9) );
AOI211_X1 g_65_1 (.ZN (n_65_1), .A (n_61_3), .B (n_55_6), .C1 (n_51_8), .C2 (n_48_8) );
AOI211_X1 g_64_3 (.ZN (n_64_3), .A (n_63_2), .B (n_57_5), .C1 (n_53_7), .C2 (n_50_7) );
AOI211_X1 g_62_4 (.ZN (n_62_4), .A (n_65_1), .B (n_59_4), .C1 (n_55_6), .C2 (n_49_9) );
AOI211_X1 g_60_5 (.ZN (n_60_5), .A (n_64_3), .B (n_61_3), .C1 (n_57_5), .C2 (n_51_8) );
AOI211_X1 g_58_6 (.ZN (n_58_6), .A (n_62_4), .B (n_63_2), .C1 (n_59_4), .C2 (n_53_7) );
AOI211_X1 g_56_7 (.ZN (n_56_7), .A (n_60_5), .B (n_65_1), .C1 (n_61_3), .C2 (n_55_6) );
AOI211_X1 g_54_8 (.ZN (n_54_8), .A (n_58_6), .B (n_64_3), .C1 (n_63_2), .C2 (n_57_5) );
AOI211_X1 g_52_9 (.ZN (n_52_9), .A (n_56_7), .B (n_62_4), .C1 (n_65_1), .C2 (n_59_4) );
AOI211_X1 g_51_7 (.ZN (n_51_7), .A (n_54_8), .B (n_60_5), .C1 (n_64_3), .C2 (n_61_3) );
AOI211_X1 g_49_8 (.ZN (n_49_8), .A (n_52_9), .B (n_58_6), .C1 (n_62_4), .C2 (n_63_2) );
AOI211_X1 g_47_9 (.ZN (n_47_9), .A (n_51_7), .B (n_56_7), .C1 (n_60_5), .C2 (n_65_1) );
AOI211_X1 g_45_10 (.ZN (n_45_10), .A (n_49_8), .B (n_54_8), .C1 (n_58_6), .C2 (n_64_3) );
AOI211_X1 g_43_9 (.ZN (n_43_9), .A (n_47_9), .B (n_52_9), .C1 (n_56_7), .C2 (n_62_4) );
AOI211_X1 g_41_10 (.ZN (n_41_10), .A (n_45_10), .B (n_51_7), .C1 (n_54_8), .C2 (n_60_5) );
AOI211_X1 g_43_11 (.ZN (n_43_11), .A (n_43_9), .B (n_49_8), .C1 (n_52_9), .C2 (n_58_6) );
AOI211_X1 g_41_12 (.ZN (n_41_12), .A (n_41_10), .B (n_47_9), .C1 (n_51_7), .C2 (n_56_7) );
AOI211_X1 g_42_10 (.ZN (n_42_10), .A (n_43_11), .B (n_45_10), .C1 (n_49_8), .C2 (n_54_8) );
AOI211_X1 g_40_11 (.ZN (n_40_11), .A (n_41_12), .B (n_43_9), .C1 (n_47_9), .C2 (n_52_9) );
AOI211_X1 g_38_12 (.ZN (n_38_12), .A (n_42_10), .B (n_41_10), .C1 (n_45_10), .C2 (n_51_7) );
AOI211_X1 g_36_13 (.ZN (n_36_13), .A (n_40_11), .B (n_43_11), .C1 (n_43_9), .C2 (n_49_8) );
AOI211_X1 g_34_14 (.ZN (n_34_14), .A (n_38_12), .B (n_41_12), .C1 (n_41_10), .C2 (n_47_9) );
AOI211_X1 g_32_15 (.ZN (n_32_15), .A (n_36_13), .B (n_42_10), .C1 (n_43_11), .C2 (n_45_10) );
AOI211_X1 g_30_16 (.ZN (n_30_16), .A (n_34_14), .B (n_40_11), .C1 (n_41_12), .C2 (n_43_9) );
AOI211_X1 g_28_17 (.ZN (n_28_17), .A (n_32_15), .B (n_38_12), .C1 (n_42_10), .C2 (n_41_10) );
AOI211_X1 g_27_19 (.ZN (n_27_19), .A (n_30_16), .B (n_36_13), .C1 (n_40_11), .C2 (n_43_11) );
AOI211_X1 g_26_17 (.ZN (n_26_17), .A (n_28_17), .B (n_34_14), .C1 (n_38_12), .C2 (n_41_12) );
AOI211_X1 g_28_16 (.ZN (n_28_16), .A (n_27_19), .B (n_32_15), .C1 (n_36_13), .C2 (n_42_10) );
AOI211_X1 g_30_15 (.ZN (n_30_15), .A (n_26_17), .B (n_30_16), .C1 (n_34_14), .C2 (n_40_11) );
AOI211_X1 g_32_14 (.ZN (n_32_14), .A (n_28_16), .B (n_28_17), .C1 (n_32_15), .C2 (n_38_12) );
AOI211_X1 g_34_15 (.ZN (n_34_15), .A (n_30_15), .B (n_27_19), .C1 (n_30_16), .C2 (n_36_13) );
AOI211_X1 g_32_16 (.ZN (n_32_16), .A (n_32_14), .B (n_26_17), .C1 (n_28_17), .C2 (n_34_14) );
AOI211_X1 g_30_17 (.ZN (n_30_17), .A (n_34_15), .B (n_28_16), .C1 (n_27_19), .C2 (n_32_15) );
AOI211_X1 g_28_18 (.ZN (n_28_18), .A (n_32_16), .B (n_30_15), .C1 (n_26_17), .C2 (n_30_16) );
AOI211_X1 g_29_16 (.ZN (n_29_16), .A (n_30_17), .B (n_32_14), .C1 (n_28_16), .C2 (n_28_17) );
AOI211_X1 g_27_17 (.ZN (n_27_17), .A (n_28_18), .B (n_34_15), .C1 (n_30_15), .C2 (n_27_19) );
AOI211_X1 g_25_18 (.ZN (n_25_18), .A (n_29_16), .B (n_32_16), .C1 (n_32_14), .C2 (n_26_17) );
AOI211_X1 g_23_19 (.ZN (n_23_19), .A (n_27_17), .B (n_30_17), .C1 (n_34_15), .C2 (n_28_16) );
AOI211_X1 g_21_20 (.ZN (n_21_20), .A (n_25_18), .B (n_28_18), .C1 (n_32_16), .C2 (n_30_15) );
AOI211_X1 g_19_19 (.ZN (n_19_19), .A (n_23_19), .B (n_29_16), .C1 (n_30_17), .C2 (n_32_14) );
AOI211_X1 g_17_18 (.ZN (n_17_18), .A (n_21_20), .B (n_27_17), .C1 (n_28_18), .C2 (n_34_15) );
AOI211_X1 g_15_17 (.ZN (n_15_17), .A (n_19_19), .B (n_25_18), .C1 (n_29_16), .C2 (n_32_16) );
AOI211_X1 g_13_16 (.ZN (n_13_16), .A (n_17_18), .B (n_23_19), .C1 (n_27_17), .C2 (n_30_17) );
AOI211_X1 g_11_15 (.ZN (n_11_15), .A (n_15_17), .B (n_21_20), .C1 (n_25_18), .C2 (n_28_18) );
AOI211_X1 g_9_14 (.ZN (n_9_14), .A (n_13_16), .B (n_19_19), .C1 (n_23_19), .C2 (n_29_16) );
AOI211_X1 g_7_15 (.ZN (n_7_15), .A (n_11_15), .B (n_17_18), .C1 (n_21_20), .C2 (n_27_17) );
AOI211_X1 g_9_16 (.ZN (n_9_16), .A (n_9_14), .B (n_15_17), .C1 (n_19_19), .C2 (n_25_18) );
AOI211_X1 g_11_17 (.ZN (n_11_17), .A (n_7_15), .B (n_13_16), .C1 (n_17_18), .C2 (n_23_19) );
AOI211_X1 g_13_18 (.ZN (n_13_18), .A (n_9_16), .B (n_11_15), .C1 (n_15_17), .C2 (n_21_20) );
AOI211_X1 g_15_19 (.ZN (n_15_19), .A (n_11_17), .B (n_9_14), .C1 (n_13_16), .C2 (n_19_19) );
AOI211_X1 g_17_20 (.ZN (n_17_20), .A (n_13_18), .B (n_7_15), .C1 (n_11_15), .C2 (n_17_18) );
AOI211_X1 g_19_21 (.ZN (n_19_21), .A (n_15_19), .B (n_9_16), .C1 (n_9_14), .C2 (n_15_17) );
AOI211_X1 g_21_22 (.ZN (n_21_22), .A (n_17_20), .B (n_11_17), .C1 (n_7_15), .C2 (n_13_16) );
AOI211_X1 g_20_20 (.ZN (n_20_20), .A (n_19_21), .B (n_13_18), .C1 (n_9_16), .C2 (n_11_15) );
AOI211_X1 g_22_19 (.ZN (n_22_19), .A (n_21_22), .B (n_15_19), .C1 (n_11_17), .C2 (n_9_14) );
AOI211_X1 g_24_18 (.ZN (n_24_18), .A (n_20_20), .B (n_17_20), .C1 (n_13_18), .C2 (n_7_15) );
AOI211_X1 g_25_20 (.ZN (n_25_20), .A (n_22_19), .B (n_19_21), .C1 (n_15_19), .C2 (n_9_16) );
AOI211_X1 g_23_21 (.ZN (n_23_21), .A (n_24_18), .B (n_21_22), .C1 (n_17_20), .C2 (n_11_17) );
AOI211_X1 g_22_23 (.ZN (n_22_23), .A (n_25_20), .B (n_20_20), .C1 (n_19_21), .C2 (n_13_18) );
AOI211_X1 g_21_21 (.ZN (n_21_21), .A (n_23_21), .B (n_22_19), .C1 (n_21_22), .C2 (n_15_19) );
AOI211_X1 g_23_20 (.ZN (n_23_20), .A (n_22_23), .B (n_24_18), .C1 (n_20_20), .C2 (n_17_20) );
AOI211_X1 g_25_19 (.ZN (n_25_19), .A (n_21_21), .B (n_25_20), .C1 (n_22_19), .C2 (n_19_21) );
AOI211_X1 g_27_18 (.ZN (n_27_18), .A (n_23_20), .B (n_23_21), .C1 (n_24_18), .C2 (n_21_22) );
AOI211_X1 g_29_17 (.ZN (n_29_17), .A (n_25_19), .B (n_22_23), .C1 (n_25_20), .C2 (n_20_20) );
AOI211_X1 g_31_16 (.ZN (n_31_16), .A (n_27_18), .B (n_21_21), .C1 (n_23_21), .C2 (n_22_19) );
AOI211_X1 g_33_15 (.ZN (n_33_15), .A (n_29_17), .B (n_23_20), .C1 (n_22_23), .C2 (n_24_18) );
AOI211_X1 g_35_14 (.ZN (n_35_14), .A (n_31_16), .B (n_25_19), .C1 (n_21_21), .C2 (n_25_20) );
AOI211_X1 g_37_13 (.ZN (n_37_13), .A (n_33_15), .B (n_27_18), .C1 (n_23_20), .C2 (n_23_21) );
AOI211_X1 g_36_15 (.ZN (n_36_15), .A (n_35_14), .B (n_29_17), .C1 (n_25_19), .C2 (n_22_23) );
AOI211_X1 g_38_14 (.ZN (n_38_14), .A (n_37_13), .B (n_31_16), .C1 (n_27_18), .C2 (n_21_21) );
AOI211_X1 g_40_13 (.ZN (n_40_13), .A (n_36_15), .B (n_33_15), .C1 (n_29_17), .C2 (n_23_20) );
AOI211_X1 g_42_12 (.ZN (n_42_12), .A (n_38_14), .B (n_35_14), .C1 (n_31_16), .C2 (n_25_19) );
AOI211_X1 g_44_11 (.ZN (n_44_11), .A (n_40_13), .B (n_37_13), .C1 (n_33_15), .C2 (n_27_18) );
AOI211_X1 g_43_13 (.ZN (n_43_13), .A (n_42_12), .B (n_36_15), .C1 (n_35_14), .C2 (n_29_17) );
AOI211_X1 g_45_12 (.ZN (n_45_12), .A (n_44_11), .B (n_38_14), .C1 (n_37_13), .C2 (n_31_16) );
AOI211_X1 g_44_10 (.ZN (n_44_10), .A (n_43_13), .B (n_40_13), .C1 (n_36_15), .C2 (n_33_15) );
AOI211_X1 g_42_11 (.ZN (n_42_11), .A (n_45_12), .B (n_42_12), .C1 (n_38_14), .C2 (n_35_14) );
AOI211_X1 g_40_12 (.ZN (n_40_12), .A (n_44_10), .B (n_44_11), .C1 (n_40_13), .C2 (n_37_13) );
AOI211_X1 g_38_13 (.ZN (n_38_13), .A (n_42_11), .B (n_43_13), .C1 (n_42_12), .C2 (n_36_15) );
AOI211_X1 g_37_15 (.ZN (n_37_15), .A (n_40_12), .B (n_45_12), .C1 (n_44_11), .C2 (n_38_14) );
AOI211_X1 g_39_14 (.ZN (n_39_14), .A (n_38_13), .B (n_44_10), .C1 (n_43_13), .C2 (n_40_13) );
AOI211_X1 g_41_13 (.ZN (n_41_13), .A (n_37_15), .B (n_42_11), .C1 (n_45_12), .C2 (n_42_12) );
AOI211_X1 g_43_12 (.ZN (n_43_12), .A (n_39_14), .B (n_40_12), .C1 (n_44_10), .C2 (n_44_11) );
AOI211_X1 g_45_11 (.ZN (n_45_11), .A (n_41_13), .B (n_38_13), .C1 (n_42_11), .C2 (n_43_13) );
AOI211_X1 g_47_10 (.ZN (n_47_10), .A (n_43_12), .B (n_37_15), .C1 (n_40_12), .C2 (n_45_12) );
AOI211_X1 g_46_12 (.ZN (n_46_12), .A (n_45_11), .B (n_39_14), .C1 (n_38_13), .C2 (n_44_10) );
AOI211_X1 g_48_11 (.ZN (n_48_11), .A (n_47_10), .B (n_41_13), .C1 (n_37_15), .C2 (n_42_11) );
AOI211_X1 g_50_10 (.ZN (n_50_10), .A (n_46_12), .B (n_43_12), .C1 (n_39_14), .C2 (n_40_12) );
AOI211_X1 g_49_12 (.ZN (n_49_12), .A (n_48_11), .B (n_45_11), .C1 (n_41_13), .C2 (n_38_13) );
AOI211_X1 g_48_10 (.ZN (n_48_10), .A (n_50_10), .B (n_47_10), .C1 (n_43_12), .C2 (n_37_15) );
AOI211_X1 g_50_9 (.ZN (n_50_9), .A (n_49_12), .B (n_46_12), .C1 (n_45_11), .C2 (n_39_14) );
AOI211_X1 g_52_8 (.ZN (n_52_8), .A (n_48_10), .B (n_48_11), .C1 (n_47_10), .C2 (n_41_13) );
AOI211_X1 g_54_7 (.ZN (n_54_7), .A (n_50_9), .B (n_50_10), .C1 (n_46_12), .C2 (n_43_12) );
AOI211_X1 g_53_9 (.ZN (n_53_9), .A (n_52_8), .B (n_49_12), .C1 (n_48_11), .C2 (n_45_11) );
AOI211_X1 g_55_8 (.ZN (n_55_8), .A (n_54_7), .B (n_48_10), .C1 (n_50_10), .C2 (n_47_10) );
AOI211_X1 g_57_7 (.ZN (n_57_7), .A (n_53_9), .B (n_50_9), .C1 (n_49_12), .C2 (n_46_12) );
AOI211_X1 g_59_6 (.ZN (n_59_6), .A (n_55_8), .B (n_52_8), .C1 (n_48_10), .C2 (n_48_11) );
AOI211_X1 g_61_5 (.ZN (n_61_5), .A (n_57_7), .B (n_54_7), .C1 (n_50_9), .C2 (n_50_10) );
AOI211_X1 g_63_4 (.ZN (n_63_4), .A (n_59_6), .B (n_53_9), .C1 (n_52_8), .C2 (n_49_12) );
AOI211_X1 g_65_3 (.ZN (n_65_3), .A (n_61_5), .B (n_55_8), .C1 (n_54_7), .C2 (n_48_10) );
AOI211_X1 g_67_2 (.ZN (n_67_2), .A (n_63_4), .B (n_57_7), .C1 (n_53_9), .C2 (n_50_9) );
AOI211_X1 g_69_1 (.ZN (n_69_1), .A (n_65_3), .B (n_59_6), .C1 (n_55_8), .C2 (n_52_8) );
AOI211_X1 g_68_3 (.ZN (n_68_3), .A (n_67_2), .B (n_61_5), .C1 (n_57_7), .C2 (n_54_7) );
AOI211_X1 g_70_2 (.ZN (n_70_2), .A (n_69_1), .B (n_63_4), .C1 (n_59_6), .C2 (n_53_9) );
AOI211_X1 g_72_1 (.ZN (n_72_1), .A (n_68_3), .B (n_65_3), .C1 (n_61_5), .C2 (n_55_8) );
AOI211_X1 g_71_3 (.ZN (n_71_3), .A (n_70_2), .B (n_67_2), .C1 (n_63_4), .C2 (n_57_7) );
AOI211_X1 g_70_1 (.ZN (n_70_1), .A (n_72_1), .B (n_69_1), .C1 (n_65_3), .C2 (n_59_6) );
AOI211_X1 g_68_2 (.ZN (n_68_2), .A (n_71_3), .B (n_68_3), .C1 (n_67_2), .C2 (n_61_5) );
AOI211_X1 g_66_3 (.ZN (n_66_3), .A (n_70_1), .B (n_70_2), .C1 (n_69_1), .C2 (n_63_4) );
AOI211_X1 g_64_4 (.ZN (n_64_4), .A (n_68_2), .B (n_72_1), .C1 (n_68_3), .C2 (n_65_3) );
AOI211_X1 g_62_5 (.ZN (n_62_5), .A (n_66_3), .B (n_71_3), .C1 (n_70_2), .C2 (n_67_2) );
AOI211_X1 g_60_6 (.ZN (n_60_6), .A (n_64_4), .B (n_70_1), .C1 (n_72_1), .C2 (n_69_1) );
AOI211_X1 g_58_7 (.ZN (n_58_7), .A (n_62_5), .B (n_68_2), .C1 (n_71_3), .C2 (n_68_3) );
AOI211_X1 g_56_8 (.ZN (n_56_8), .A (n_60_6), .B (n_66_3), .C1 (n_70_1), .C2 (n_70_2) );
AOI211_X1 g_54_9 (.ZN (n_54_9), .A (n_58_7), .B (n_64_4), .C1 (n_68_2), .C2 (n_72_1) );
AOI211_X1 g_55_7 (.ZN (n_55_7), .A (n_56_8), .B (n_62_5), .C1 (n_66_3), .C2 (n_71_3) );
AOI211_X1 g_53_8 (.ZN (n_53_8), .A (n_54_9), .B (n_60_6), .C1 (n_64_4), .C2 (n_70_1) );
AOI211_X1 g_51_9 (.ZN (n_51_9), .A (n_55_7), .B (n_58_7), .C1 (n_62_5), .C2 (n_68_2) );
AOI211_X1 g_49_10 (.ZN (n_49_10), .A (n_53_8), .B (n_56_8), .C1 (n_60_6), .C2 (n_66_3) );
AOI211_X1 g_51_11 (.ZN (n_51_11), .A (n_51_9), .B (n_54_9), .C1 (n_58_7), .C2 (n_64_4) );
AOI211_X1 g_53_10 (.ZN (n_53_10), .A (n_49_10), .B (n_55_7), .C1 (n_56_8), .C2 (n_62_5) );
AOI211_X1 g_55_9 (.ZN (n_55_9), .A (n_51_11), .B (n_53_8), .C1 (n_54_9), .C2 (n_60_6) );
AOI211_X1 g_57_8 (.ZN (n_57_8), .A (n_53_10), .B (n_51_9), .C1 (n_55_7), .C2 (n_58_7) );
AOI211_X1 g_59_7 (.ZN (n_59_7), .A (n_55_9), .B (n_49_10), .C1 (n_53_8), .C2 (n_56_8) );
AOI211_X1 g_61_6 (.ZN (n_61_6), .A (n_57_8), .B (n_51_11), .C1 (n_51_9), .C2 (n_54_9) );
AOI211_X1 g_60_8 (.ZN (n_60_8), .A (n_59_7), .B (n_53_10), .C1 (n_49_10), .C2 (n_55_7) );
AOI211_X1 g_62_7 (.ZN (n_62_7), .A (n_61_6), .B (n_55_9), .C1 (n_51_11), .C2 (n_53_8) );
AOI211_X1 g_64_6 (.ZN (n_64_6), .A (n_60_8), .B (n_57_8), .C1 (n_53_10), .C2 (n_51_9) );
AOI211_X1 g_66_5 (.ZN (n_66_5), .A (n_62_7), .B (n_59_7), .C1 (n_55_9), .C2 (n_49_10) );
AOI211_X1 g_68_4 (.ZN (n_68_4), .A (n_64_6), .B (n_61_6), .C1 (n_57_8), .C2 (n_51_11) );
AOI211_X1 g_70_3 (.ZN (n_70_3), .A (n_66_5), .B (n_60_8), .C1 (n_59_7), .C2 (n_53_10) );
AOI211_X1 g_72_2 (.ZN (n_72_2), .A (n_68_4), .B (n_62_7), .C1 (n_61_6), .C2 (n_55_9) );
AOI211_X1 g_74_1 (.ZN (n_74_1), .A (n_70_3), .B (n_64_6), .C1 (n_60_8), .C2 (n_57_8) );
AOI211_X1 g_75_3 (.ZN (n_75_3), .A (n_72_2), .B (n_66_5), .C1 (n_62_7), .C2 (n_59_7) );
AOI211_X1 g_76_1 (.ZN (n_76_1), .A (n_74_1), .B (n_68_4), .C1 (n_64_6), .C2 (n_61_6) );
AOI211_X1 g_74_2 (.ZN (n_74_2), .A (n_75_3), .B (n_70_3), .C1 (n_66_5), .C2 (n_60_8) );
AOI211_X1 g_73_4 (.ZN (n_73_4), .A (n_76_1), .B (n_72_2), .C1 (n_68_4), .C2 (n_62_7) );
AOI211_X1 g_71_5 (.ZN (n_71_5), .A (n_74_2), .B (n_74_1), .C1 (n_70_3), .C2 (n_64_6) );
AOI211_X1 g_69_4 (.ZN (n_69_4), .A (n_73_4), .B (n_75_3), .C1 (n_72_2), .C2 (n_66_5) );
AOI211_X1 g_67_5 (.ZN (n_67_5), .A (n_71_5), .B (n_76_1), .C1 (n_74_1), .C2 (n_68_4) );
AOI211_X1 g_65_6 (.ZN (n_65_6), .A (n_69_4), .B (n_74_2), .C1 (n_75_3), .C2 (n_70_3) );
AOI211_X1 g_66_4 (.ZN (n_66_4), .A (n_67_5), .B (n_73_4), .C1 (n_76_1), .C2 (n_72_2) );
AOI211_X1 g_64_5 (.ZN (n_64_5), .A (n_65_6), .B (n_71_5), .C1 (n_74_2), .C2 (n_74_1) );
AOI211_X1 g_62_6 (.ZN (n_62_6), .A (n_66_4), .B (n_69_4), .C1 (n_73_4), .C2 (n_75_3) );
AOI211_X1 g_60_7 (.ZN (n_60_7), .A (n_64_5), .B (n_67_5), .C1 (n_71_5), .C2 (n_76_1) );
AOI211_X1 g_58_8 (.ZN (n_58_8), .A (n_62_6), .B (n_65_6), .C1 (n_69_4), .C2 (n_74_2) );
AOI211_X1 g_56_9 (.ZN (n_56_9), .A (n_60_7), .B (n_66_4), .C1 (n_67_5), .C2 (n_73_4) );
AOI211_X1 g_54_10 (.ZN (n_54_10), .A (n_58_8), .B (n_64_5), .C1 (n_65_6), .C2 (n_71_5) );
AOI211_X1 g_52_11 (.ZN (n_52_11), .A (n_56_9), .B (n_62_6), .C1 (n_66_4), .C2 (n_69_4) );
AOI211_X1 g_50_12 (.ZN (n_50_12), .A (n_54_10), .B (n_60_7), .C1 (n_64_5), .C2 (n_67_5) );
AOI211_X1 g_51_10 (.ZN (n_51_10), .A (n_52_11), .B (n_58_8), .C1 (n_62_6), .C2 (n_65_6) );
AOI211_X1 g_49_11 (.ZN (n_49_11), .A (n_50_12), .B (n_56_9), .C1 (n_60_7), .C2 (n_66_4) );
AOI211_X1 g_47_12 (.ZN (n_47_12), .A (n_51_10), .B (n_54_10), .C1 (n_58_8), .C2 (n_64_5) );
AOI211_X1 g_45_13 (.ZN (n_45_13), .A (n_49_11), .B (n_52_11), .C1 (n_56_9), .C2 (n_62_6) );
AOI211_X1 g_46_11 (.ZN (n_46_11), .A (n_47_12), .B (n_50_12), .C1 (n_54_10), .C2 (n_60_7) );
AOI211_X1 g_44_12 (.ZN (n_44_12), .A (n_45_13), .B (n_51_10), .C1 (n_52_11), .C2 (n_58_8) );
AOI211_X1 g_42_13 (.ZN (n_42_13), .A (n_46_11), .B (n_49_11), .C1 (n_50_12), .C2 (n_56_9) );
AOI211_X1 g_40_14 (.ZN (n_40_14), .A (n_44_12), .B (n_47_12), .C1 (n_51_10), .C2 (n_54_10) );
AOI211_X1 g_38_15 (.ZN (n_38_15), .A (n_42_13), .B (n_45_13), .C1 (n_49_11), .C2 (n_52_11) );
AOI211_X1 g_39_13 (.ZN (n_39_13), .A (n_40_14), .B (n_46_11), .C1 (n_47_12), .C2 (n_50_12) );
AOI211_X1 g_37_14 (.ZN (n_37_14), .A (n_38_15), .B (n_44_12), .C1 (n_45_13), .C2 (n_51_10) );
AOI211_X1 g_35_15 (.ZN (n_35_15), .A (n_39_13), .B (n_42_13), .C1 (n_46_11), .C2 (n_49_11) );
AOI211_X1 g_33_16 (.ZN (n_33_16), .A (n_37_14), .B (n_40_14), .C1 (n_44_12), .C2 (n_47_12) );
AOI211_X1 g_31_17 (.ZN (n_31_17), .A (n_35_15), .B (n_38_15), .C1 (n_42_13), .C2 (n_45_13) );
AOI211_X1 g_29_18 (.ZN (n_29_18), .A (n_33_16), .B (n_39_13), .C1 (n_40_14), .C2 (n_46_11) );
AOI211_X1 g_28_20 (.ZN (n_28_20), .A (n_31_17), .B (n_37_14), .C1 (n_38_15), .C2 (n_44_12) );
AOI211_X1 g_26_19 (.ZN (n_26_19), .A (n_29_18), .B (n_35_15), .C1 (n_39_13), .C2 (n_42_13) );
AOI211_X1 g_24_20 (.ZN (n_24_20), .A (n_28_20), .B (n_33_16), .C1 (n_37_14), .C2 (n_40_14) );
AOI211_X1 g_22_21 (.ZN (n_22_21), .A (n_26_19), .B (n_31_17), .C1 (n_35_15), .C2 (n_38_15) );
AOI211_X1 g_20_22 (.ZN (n_20_22), .A (n_24_20), .B (n_29_18), .C1 (n_33_16), .C2 (n_39_13) );
AOI211_X1 g_18_21 (.ZN (n_18_21), .A (n_22_21), .B (n_28_20), .C1 (n_31_17), .C2 (n_37_14) );
AOI211_X1 g_16_20 (.ZN (n_16_20), .A (n_20_22), .B (n_26_19), .C1 (n_29_18), .C2 (n_35_15) );
AOI211_X1 g_14_19 (.ZN (n_14_19), .A (n_18_21), .B (n_24_20), .C1 (n_28_20), .C2 (n_33_16) );
AOI211_X1 g_12_18 (.ZN (n_12_18), .A (n_16_20), .B (n_22_21), .C1 (n_26_19), .C2 (n_31_17) );
AOI211_X1 g_10_17 (.ZN (n_10_17), .A (n_14_19), .B (n_20_22), .C1 (n_24_20), .C2 (n_29_18) );
AOI211_X1 g_8_16 (.ZN (n_8_16), .A (n_12_18), .B (n_18_21), .C1 (n_22_21), .C2 (n_28_20) );
AOI211_X1 g_6_17 (.ZN (n_6_17), .A (n_10_17), .B (n_16_20), .C1 (n_20_22), .C2 (n_26_19) );
AOI211_X1 g_4_16 (.ZN (n_4_16), .A (n_8_16), .B (n_14_19), .C1 (n_18_21), .C2 (n_24_20) );
AOI211_X1 g_3_18 (.ZN (n_3_18), .A (n_6_17), .B (n_12_18), .C1 (n_16_20), .C2 (n_22_21) );
AOI211_X1 g_2_20 (.ZN (n_2_20), .A (n_4_16), .B (n_10_17), .C1 (n_14_19), .C2 (n_20_22) );
AOI211_X1 g_3_22 (.ZN (n_3_22), .A (n_3_18), .B (n_8_16), .C1 (n_12_18), .C2 (n_18_21) );
AOI211_X1 g_4_20 (.ZN (n_4_20), .A (n_2_20), .B (n_6_17), .C1 (n_10_17), .C2 (n_16_20) );
AOI211_X1 g_5_18 (.ZN (n_5_18), .A (n_3_22), .B (n_4_16), .C1 (n_8_16), .C2 (n_14_19) );
AOI211_X1 g_3_17 (.ZN (n_3_17), .A (n_4_20), .B (n_3_18), .C1 (n_6_17), .C2 (n_12_18) );
AOI211_X1 g_4_15 (.ZN (n_4_15), .A (n_5_18), .B (n_2_20), .C1 (n_4_16), .C2 (n_10_17) );
AOI211_X1 g_6_14 (.ZN (n_6_14), .A (n_3_17), .B (n_3_22), .C1 (n_3_18), .C2 (n_8_16) );
AOI211_X1 g_5_16 (.ZN (n_5_16), .A (n_4_15), .B (n_4_20), .C1 (n_2_20), .C2 (n_6_17) );
AOI211_X1 g_4_18 (.ZN (n_4_18), .A (n_6_14), .B (n_5_18), .C1 (n_3_22), .C2 (n_4_16) );
AOI211_X1 g_3_16 (.ZN (n_3_16), .A (n_5_16), .B (n_3_17), .C1 (n_4_20), .C2 (n_3_18) );
AOI211_X1 g_5_15 (.ZN (n_5_15), .A (n_4_18), .B (n_4_15), .C1 (n_5_18), .C2 (n_2_20) );
AOI211_X1 g_4_17 (.ZN (n_4_17), .A (n_3_16), .B (n_6_14), .C1 (n_3_17), .C2 (n_3_22) );
AOI211_X1 g_2_18 (.ZN (n_2_18), .A (n_5_15), .B (n_5_16), .C1 (n_4_15), .C2 (n_4_20) );
AOI211_X1 g_3_20 (.ZN (n_3_20), .A (n_4_17), .B (n_4_18), .C1 (n_6_14), .C2 (n_5_18) );
AOI211_X1 g_5_19 (.ZN (n_5_19), .A (n_2_18), .B (n_3_16), .C1 (n_5_16), .C2 (n_3_17) );
AOI211_X1 g_4_21 (.ZN (n_4_21), .A (n_3_20), .B (n_5_15), .C1 (n_4_18), .C2 (n_4_15) );
AOI211_X1 g_2_22 (.ZN (n_2_22), .A (n_5_19), .B (n_4_17), .C1 (n_3_16), .C2 (n_6_14) );
AOI211_X1 g_1_24 (.ZN (n_1_24), .A (n_4_21), .B (n_2_18), .C1 (n_5_15), .C2 (n_5_16) );
AOI211_X1 g_3_23 (.ZN (n_3_23), .A (n_2_22), .B (n_3_20), .C1 (n_4_17), .C2 (n_4_18) );
AOI211_X1 g_5_22 (.ZN (n_5_22), .A (n_1_24), .B (n_5_19), .C1 (n_2_18), .C2 (n_3_16) );
AOI211_X1 g_4_24 (.ZN (n_4_24), .A (n_3_23), .B (n_4_21), .C1 (n_3_20), .C2 (n_5_15) );
AOI211_X1 g_5_26 (.ZN (n_5_26), .A (n_5_22), .B (n_2_22), .C1 (n_5_19), .C2 (n_4_17) );
AOI211_X1 g_3_25 (.ZN (n_3_25), .A (n_4_24), .B (n_1_24), .C1 (n_4_21), .C2 (n_2_18) );
AOI211_X1 g_4_23 (.ZN (n_4_23), .A (n_5_26), .B (n_3_23), .C1 (n_2_22), .C2 (n_3_20) );
AOI211_X1 g_5_21 (.ZN (n_5_21), .A (n_3_25), .B (n_5_22), .C1 (n_1_24), .C2 (n_5_19) );
AOI211_X1 g_4_19 (.ZN (n_4_19), .A (n_4_23), .B (n_4_24), .C1 (n_3_23), .C2 (n_4_21) );
AOI211_X1 g_5_17 (.ZN (n_5_17), .A (n_5_21), .B (n_5_26), .C1 (n_5_22), .C2 (n_2_22) );
AOI211_X1 g_7_16 (.ZN (n_7_16), .A (n_4_19), .B (n_3_25), .C1 (n_4_24), .C2 (n_1_24) );
AOI211_X1 g_6_18 (.ZN (n_6_18), .A (n_5_17), .B (n_4_23), .C1 (n_5_26), .C2 (n_3_23) );
AOI211_X1 g_5_20 (.ZN (n_5_20), .A (n_7_16), .B (n_5_21), .C1 (n_3_25), .C2 (n_5_22) );
AOI211_X1 g_4_22 (.ZN (n_4_22), .A (n_6_18), .B (n_4_19), .C1 (n_4_23), .C2 (n_4_24) );
AOI211_X1 g_3_24 (.ZN (n_3_24), .A (n_5_20), .B (n_5_17), .C1 (n_5_21), .C2 (n_5_26) );
AOI211_X1 g_2_26 (.ZN (n_2_26), .A (n_4_22), .B (n_7_16), .C1 (n_4_19), .C2 (n_3_25) );
AOI211_X1 g_4_25 (.ZN (n_4_25), .A (n_3_24), .B (n_6_18), .C1 (n_5_17), .C2 (n_4_23) );
AOI211_X1 g_6_24 (.ZN (n_6_24), .A (n_2_26), .B (n_5_20), .C1 (n_7_16), .C2 (n_5_21) );
AOI211_X1 g_7_22 (.ZN (n_7_22), .A (n_4_25), .B (n_4_22), .C1 (n_6_18), .C2 (n_4_19) );
AOI211_X1 g_6_20 (.ZN (n_6_20), .A (n_6_24), .B (n_3_24), .C1 (n_5_20), .C2 (n_5_17) );
AOI211_X1 g_7_18 (.ZN (n_7_18), .A (n_7_22), .B (n_2_26), .C1 (n_4_22), .C2 (n_7_16) );
AOI211_X1 g_6_16 (.ZN (n_6_16), .A (n_6_20), .B (n_4_25), .C1 (n_3_24), .C2 (n_6_18) );
AOI211_X1 g_8_15 (.ZN (n_8_15), .A (n_7_18), .B (n_6_24), .C1 (n_2_26), .C2 (n_5_20) );
AOI211_X1 g_7_17 (.ZN (n_7_17), .A (n_6_16), .B (n_7_22), .C1 (n_4_25), .C2 (n_4_22) );
AOI211_X1 g_6_19 (.ZN (n_6_19), .A (n_8_15), .B (n_6_20), .C1 (n_6_24), .C2 (n_3_24) );
AOI211_X1 g_8_18 (.ZN (n_8_18), .A (n_7_17), .B (n_7_18), .C1 (n_7_22), .C2 (n_2_26) );
AOI211_X1 g_7_20 (.ZN (n_7_20), .A (n_6_19), .B (n_6_16), .C1 (n_6_20), .C2 (n_4_25) );
AOI211_X1 g_6_22 (.ZN (n_6_22), .A (n_8_18), .B (n_8_15), .C1 (n_7_18), .C2 (n_6_24) );
AOI211_X1 g_5_24 (.ZN (n_5_24), .A (n_7_20), .B (n_7_17), .C1 (n_6_16), .C2 (n_7_22) );
AOI211_X1 g_4_26 (.ZN (n_4_26), .A (n_6_22), .B (n_6_19), .C1 (n_8_15), .C2 (n_6_20) );
AOI211_X1 g_3_28 (.ZN (n_3_28), .A (n_5_24), .B (n_8_18), .C1 (n_7_17), .C2 (n_7_18) );
AOI211_X1 g_2_30 (.ZN (n_2_30), .A (n_4_26), .B (n_7_20), .C1 (n_6_19), .C2 (n_6_16) );
AOI211_X1 g_4_29 (.ZN (n_4_29), .A (n_3_28), .B (n_6_22), .C1 (n_8_18), .C2 (n_8_15) );
AOI211_X1 g_5_27 (.ZN (n_5_27), .A (n_2_30), .B (n_5_24), .C1 (n_7_20), .C2 (n_7_17) );
AOI211_X1 g_6_25 (.ZN (n_6_25), .A (n_4_29), .B (n_4_26), .C1 (n_6_22), .C2 (n_6_19) );
AOI211_X1 g_5_23 (.ZN (n_5_23), .A (n_5_27), .B (n_3_28), .C1 (n_5_24), .C2 (n_8_18) );
AOI211_X1 g_6_21 (.ZN (n_6_21), .A (n_6_25), .B (n_2_30), .C1 (n_4_26), .C2 (n_7_20) );
AOI211_X1 g_8_20 (.ZN (n_8_20), .A (n_5_23), .B (n_4_29), .C1 (n_3_28), .C2 (n_6_22) );
AOI211_X1 g_10_19 (.ZN (n_10_19), .A (n_6_21), .B (n_5_27), .C1 (n_2_30), .C2 (n_5_24) );
AOI211_X1 g_9_17 (.ZN (n_9_17), .A (n_8_20), .B (n_6_25), .C1 (n_4_29), .C2 (n_4_26) );
AOI211_X1 g_8_19 (.ZN (n_8_19), .A (n_10_19), .B (n_5_23), .C1 (n_5_27), .C2 (n_3_28) );
AOI211_X1 g_7_21 (.ZN (n_7_21), .A (n_9_17), .B (n_6_21), .C1 (n_6_25), .C2 (n_2_30) );
AOI211_X1 g_6_23 (.ZN (n_6_23), .A (n_8_19), .B (n_8_20), .C1 (n_5_23), .C2 (n_4_29) );
AOI211_X1 g_5_25 (.ZN (n_5_25), .A (n_7_21), .B (n_10_19), .C1 (n_6_21), .C2 (n_5_27) );
AOI211_X1 g_4_27 (.ZN (n_4_27), .A (n_6_23), .B (n_9_17), .C1 (n_8_20), .C2 (n_6_25) );
AOI211_X1 g_6_28 (.ZN (n_6_28), .A (n_5_25), .B (n_8_19), .C1 (n_10_19), .C2 (n_5_23) );
AOI211_X1 g_7_26 (.ZN (n_7_26), .A (n_4_27), .B (n_7_21), .C1 (n_9_17), .C2 (n_6_21) );
AOI211_X1 g_8_24 (.ZN (n_8_24), .A (n_6_28), .B (n_6_23), .C1 (n_8_19), .C2 (n_8_20) );
AOI211_X1 g_9_22 (.ZN (n_9_22), .A (n_7_26), .B (n_5_25), .C1 (n_7_21), .C2 (n_10_19) );
AOI211_X1 g_7_23 (.ZN (n_7_23), .A (n_8_24), .B (n_4_27), .C1 (n_6_23), .C2 (n_9_17) );
AOI211_X1 g_8_21 (.ZN (n_8_21), .A (n_9_22), .B (n_6_28), .C1 (n_5_25), .C2 (n_8_19) );
AOI211_X1 g_7_19 (.ZN (n_7_19), .A (n_7_23), .B (n_7_26), .C1 (n_4_27), .C2 (n_7_21) );
AOI211_X1 g_9_18 (.ZN (n_9_18), .A (n_8_21), .B (n_8_24), .C1 (n_6_28), .C2 (n_6_23) );
AOI211_X1 g_10_16 (.ZN (n_10_16), .A (n_7_19), .B (n_9_22), .C1 (n_7_26), .C2 (n_5_25) );
AOI211_X1 g_8_17 (.ZN (n_8_17), .A (n_9_18), .B (n_7_23), .C1 (n_8_24), .C2 (n_4_27) );
AOI211_X1 g_9_19 (.ZN (n_9_19), .A (n_10_16), .B (n_8_21), .C1 (n_9_22), .C2 (n_6_28) );
AOI211_X1 g_11_18 (.ZN (n_11_18), .A (n_8_17), .B (n_7_19), .C1 (n_7_23), .C2 (n_7_26) );
AOI211_X1 g_10_20 (.ZN (n_10_20), .A (n_9_19), .B (n_9_18), .C1 (n_8_21), .C2 (n_8_24) );
AOI211_X1 g_12_19 (.ZN (n_12_19), .A (n_11_18), .B (n_10_16), .C1 (n_7_19), .C2 (n_9_22) );
AOI211_X1 g_10_18 (.ZN (n_10_18), .A (n_10_20), .B (n_8_17), .C1 (n_9_18), .C2 (n_7_23) );
AOI211_X1 g_12_17 (.ZN (n_12_17), .A (n_12_19), .B (n_9_19), .C1 (n_10_16), .C2 (n_8_21) );
AOI211_X1 g_14_18 (.ZN (n_14_18), .A (n_10_18), .B (n_11_18), .C1 (n_8_17), .C2 (n_7_19) );
AOI211_X1 g_16_19 (.ZN (n_16_19), .A (n_12_17), .B (n_10_20), .C1 (n_9_19), .C2 (n_9_18) );
AOI211_X1 g_14_20 (.ZN (n_14_20), .A (n_14_18), .B (n_12_19), .C1 (n_11_18), .C2 (n_10_16) );
AOI211_X1 g_16_21 (.ZN (n_16_21), .A (n_16_19), .B (n_10_18), .C1 (n_10_20), .C2 (n_8_17) );
AOI211_X1 g_18_20 (.ZN (n_18_20), .A (n_14_20), .B (n_12_17), .C1 (n_12_19), .C2 (n_9_19) );
AOI211_X1 g_20_21 (.ZN (n_20_21), .A (n_16_21), .B (n_14_18), .C1 (n_10_18), .C2 (n_11_18) );
AOI211_X1 g_18_22 (.ZN (n_18_22), .A (n_18_20), .B (n_16_19), .C1 (n_12_17), .C2 (n_10_20) );
AOI211_X1 g_20_23 (.ZN (n_20_23), .A (n_20_21), .B (n_14_20), .C1 (n_14_18), .C2 (n_12_19) );
AOI211_X1 g_22_22 (.ZN (n_22_22), .A (n_18_22), .B (n_16_21), .C1 (n_16_19), .C2 (n_10_18) );
AOI211_X1 g_24_21 (.ZN (n_24_21), .A (n_20_23), .B (n_18_20), .C1 (n_14_20), .C2 (n_12_17) );
AOI211_X1 g_26_20 (.ZN (n_26_20), .A (n_22_22), .B (n_20_21), .C1 (n_16_21), .C2 (n_14_18) );
AOI211_X1 g_28_19 (.ZN (n_28_19), .A (n_24_21), .B (n_18_22), .C1 (n_18_20), .C2 (n_16_19) );
AOI211_X1 g_30_18 (.ZN (n_30_18), .A (n_26_20), .B (n_20_23), .C1 (n_20_21), .C2 (n_14_20) );
AOI211_X1 g_32_17 (.ZN (n_32_17), .A (n_28_19), .B (n_22_22), .C1 (n_18_22), .C2 (n_16_21) );
AOI211_X1 g_34_16 (.ZN (n_34_16), .A (n_30_18), .B (n_24_21), .C1 (n_20_23), .C2 (n_18_20) );
AOI211_X1 g_33_18 (.ZN (n_33_18), .A (n_32_17), .B (n_26_20), .C1 (n_22_22), .C2 (n_20_21) );
AOI211_X1 g_35_17 (.ZN (n_35_17), .A (n_34_16), .B (n_28_19), .C1 (n_24_21), .C2 (n_18_22) );
AOI211_X1 g_37_16 (.ZN (n_37_16), .A (n_33_18), .B (n_30_18), .C1 (n_26_20), .C2 (n_20_23) );
AOI211_X1 g_39_15 (.ZN (n_39_15), .A (n_35_17), .B (n_32_17), .C1 (n_28_19), .C2 (n_22_22) );
AOI211_X1 g_41_14 (.ZN (n_41_14), .A (n_37_16), .B (n_34_16), .C1 (n_30_18), .C2 (n_24_21) );
AOI211_X1 g_40_16 (.ZN (n_40_16), .A (n_39_15), .B (n_33_18), .C1 (n_32_17), .C2 (n_26_20) );
AOI211_X1 g_42_15 (.ZN (n_42_15), .A (n_41_14), .B (n_35_17), .C1 (n_34_16), .C2 (n_28_19) );
AOI211_X1 g_44_14 (.ZN (n_44_14), .A (n_40_16), .B (n_37_16), .C1 (n_33_18), .C2 (n_30_18) );
AOI211_X1 g_46_13 (.ZN (n_46_13), .A (n_42_15), .B (n_39_15), .C1 (n_35_17), .C2 (n_32_17) );
AOI211_X1 g_48_12 (.ZN (n_48_12), .A (n_44_14), .B (n_41_14), .C1 (n_37_16), .C2 (n_34_16) );
AOI211_X1 g_50_11 (.ZN (n_50_11), .A (n_46_13), .B (n_40_16), .C1 (n_39_15), .C2 (n_33_18) );
AOI211_X1 g_52_10 (.ZN (n_52_10), .A (n_48_12), .B (n_42_15), .C1 (n_41_14), .C2 (n_35_17) );
AOI211_X1 g_51_12 (.ZN (n_51_12), .A (n_50_11), .B (n_44_14), .C1 (n_40_16), .C2 (n_37_16) );
AOI211_X1 g_53_11 (.ZN (n_53_11), .A (n_52_10), .B (n_46_13), .C1 (n_42_15), .C2 (n_39_15) );
AOI211_X1 g_55_10 (.ZN (n_55_10), .A (n_51_12), .B (n_48_12), .C1 (n_44_14), .C2 (n_41_14) );
AOI211_X1 g_57_9 (.ZN (n_57_9), .A (n_53_11), .B (n_50_11), .C1 (n_46_13), .C2 (n_40_16) );
AOI211_X1 g_59_8 (.ZN (n_59_8), .A (n_55_10), .B (n_52_10), .C1 (n_48_12), .C2 (n_42_15) );
AOI211_X1 g_61_7 (.ZN (n_61_7), .A (n_57_9), .B (n_51_12), .C1 (n_50_11), .C2 (n_44_14) );
AOI211_X1 g_63_6 (.ZN (n_63_6), .A (n_59_8), .B (n_53_11), .C1 (n_52_10), .C2 (n_46_13) );
AOI211_X1 g_65_5 (.ZN (n_65_5), .A (n_61_7), .B (n_55_10), .C1 (n_51_12), .C2 (n_48_12) );
AOI211_X1 g_67_4 (.ZN (n_67_4), .A (n_63_6), .B (n_57_9), .C1 (n_53_11), .C2 (n_50_11) );
AOI211_X1 g_69_3 (.ZN (n_69_3), .A (n_65_5), .B (n_59_8), .C1 (n_55_10), .C2 (n_52_10) );
AOI211_X1 g_71_2 (.ZN (n_71_2), .A (n_67_4), .B (n_61_7), .C1 (n_57_9), .C2 (n_51_12) );
AOI211_X1 g_73_1 (.ZN (n_73_1), .A (n_69_3), .B (n_63_6), .C1 (n_59_8), .C2 (n_53_11) );
AOI211_X1 g_72_3 (.ZN (n_72_3), .A (n_71_2), .B (n_65_5), .C1 (n_61_7), .C2 (n_55_10) );
AOI211_X1 g_70_4 (.ZN (n_70_4), .A (n_73_1), .B (n_67_4), .C1 (n_63_6), .C2 (n_57_9) );
AOI211_X1 g_68_5 (.ZN (n_68_5), .A (n_72_3), .B (n_69_3), .C1 (n_65_5), .C2 (n_59_8) );
AOI211_X1 g_66_6 (.ZN (n_66_6), .A (n_70_4), .B (n_71_2), .C1 (n_67_4), .C2 (n_61_7) );
AOI211_X1 g_64_7 (.ZN (n_64_7), .A (n_68_5), .B (n_73_1), .C1 (n_69_3), .C2 (n_63_6) );
AOI211_X1 g_62_8 (.ZN (n_62_8), .A (n_66_6), .B (n_72_3), .C1 (n_71_2), .C2 (n_65_5) );
AOI211_X1 g_60_9 (.ZN (n_60_9), .A (n_64_7), .B (n_70_4), .C1 (n_73_1), .C2 (n_67_4) );
AOI211_X1 g_58_10 (.ZN (n_58_10), .A (n_62_8), .B (n_68_5), .C1 (n_72_3), .C2 (n_69_3) );
AOI211_X1 g_56_11 (.ZN (n_56_11), .A (n_60_9), .B (n_66_6), .C1 (n_70_4), .C2 (n_71_2) );
AOI211_X1 g_54_12 (.ZN (n_54_12), .A (n_58_10), .B (n_64_7), .C1 (n_68_5), .C2 (n_73_1) );
AOI211_X1 g_52_13 (.ZN (n_52_13), .A (n_56_11), .B (n_62_8), .C1 (n_66_6), .C2 (n_72_3) );
AOI211_X1 g_50_14 (.ZN (n_50_14), .A (n_54_12), .B (n_60_9), .C1 (n_64_7), .C2 (n_70_4) );
AOI211_X1 g_48_13 (.ZN (n_48_13), .A (n_52_13), .B (n_58_10), .C1 (n_62_8), .C2 (n_68_5) );
AOI211_X1 g_46_14 (.ZN (n_46_14), .A (n_50_14), .B (n_56_11), .C1 (n_60_9), .C2 (n_66_6) );
AOI211_X1 g_44_13 (.ZN (n_44_13), .A (n_48_13), .B (n_54_12), .C1 (n_58_10), .C2 (n_64_7) );
AOI211_X1 g_42_14 (.ZN (n_42_14), .A (n_46_14), .B (n_52_13), .C1 (n_56_11), .C2 (n_62_8) );
AOI211_X1 g_40_15 (.ZN (n_40_15), .A (n_44_13), .B (n_50_14), .C1 (n_54_12), .C2 (n_60_9) );
AOI211_X1 g_38_16 (.ZN (n_38_16), .A (n_42_14), .B (n_48_13), .C1 (n_52_13), .C2 (n_58_10) );
AOI211_X1 g_36_17 (.ZN (n_36_17), .A (n_40_15), .B (n_46_14), .C1 (n_50_14), .C2 (n_56_11) );
AOI211_X1 g_34_18 (.ZN (n_34_18), .A (n_38_16), .B (n_44_13), .C1 (n_48_13), .C2 (n_54_12) );
AOI211_X1 g_35_16 (.ZN (n_35_16), .A (n_36_17), .B (n_42_14), .C1 (n_46_14), .C2 (n_52_13) );
AOI211_X1 g_33_17 (.ZN (n_33_17), .A (n_34_18), .B (n_40_15), .C1 (n_44_13), .C2 (n_50_14) );
AOI211_X1 g_31_18 (.ZN (n_31_18), .A (n_35_16), .B (n_38_16), .C1 (n_42_14), .C2 (n_48_13) );
AOI211_X1 g_29_19 (.ZN (n_29_19), .A (n_33_17), .B (n_36_17), .C1 (n_40_15), .C2 (n_46_14) );
AOI211_X1 g_27_20 (.ZN (n_27_20), .A (n_31_18), .B (n_34_18), .C1 (n_38_16), .C2 (n_44_13) );
AOI211_X1 g_25_21 (.ZN (n_25_21), .A (n_29_19), .B (n_35_16), .C1 (n_36_17), .C2 (n_42_14) );
AOI211_X1 g_23_22 (.ZN (n_23_22), .A (n_27_20), .B (n_33_17), .C1 (n_34_18), .C2 (n_40_15) );
AOI211_X1 g_21_23 (.ZN (n_21_23), .A (n_25_21), .B (n_31_18), .C1 (n_35_16), .C2 (n_38_16) );
AOI211_X1 g_19_22 (.ZN (n_19_22), .A (n_23_22), .B (n_29_19), .C1 (n_33_17), .C2 (n_36_17) );
AOI211_X1 g_17_21 (.ZN (n_17_21), .A (n_21_23), .B (n_27_20), .C1 (n_31_18), .C2 (n_34_18) );
AOI211_X1 g_15_20 (.ZN (n_15_20), .A (n_19_22), .B (n_25_21), .C1 (n_29_19), .C2 (n_35_16) );
AOI211_X1 g_13_19 (.ZN (n_13_19), .A (n_17_21), .B (n_23_22), .C1 (n_27_20), .C2 (n_33_17) );
AOI211_X1 g_11_20 (.ZN (n_11_20), .A (n_15_20), .B (n_21_23), .C1 (n_25_21), .C2 (n_31_18) );
AOI211_X1 g_9_21 (.ZN (n_9_21), .A (n_13_19), .B (n_19_22), .C1 (n_23_22), .C2 (n_29_19) );
AOI211_X1 g_8_23 (.ZN (n_8_23), .A (n_11_20), .B (n_17_21), .C1 (n_21_23), .C2 (n_27_20) );
AOI211_X1 g_7_25 (.ZN (n_7_25), .A (n_9_21), .B (n_15_20), .C1 (n_19_22), .C2 (n_25_21) );
AOI211_X1 g_6_27 (.ZN (n_6_27), .A (n_8_23), .B (n_13_19), .C1 (n_17_21), .C2 (n_23_22) );
AOI211_X1 g_5_29 (.ZN (n_5_29), .A (n_7_25), .B (n_11_20), .C1 (n_15_20), .C2 (n_21_23) );
AOI211_X1 g_4_31 (.ZN (n_4_31), .A (n_6_27), .B (n_9_21), .C1 (n_13_19), .C2 (n_19_22) );
AOI211_X1 g_6_32 (.ZN (n_6_32), .A (n_5_29), .B (n_8_23), .C1 (n_11_20), .C2 (n_17_21) );
AOI211_X1 g_4_33 (.ZN (n_4_33), .A (n_4_31), .B (n_7_25), .C1 (n_9_21), .C2 (n_15_20) );
AOI211_X1 g_2_34 (.ZN (n_2_34), .A (n_6_32), .B (n_6_27), .C1 (n_8_23), .C2 (n_13_19) );
AOI211_X1 g_3_32 (.ZN (n_3_32), .A (n_4_33), .B (n_5_29), .C1 (n_7_25), .C2 (n_11_20) );
AOI211_X1 g_5_31 (.ZN (n_5_31), .A (n_2_34), .B (n_4_31), .C1 (n_6_27), .C2 (n_9_21) );
AOI211_X1 g_7_30 (.ZN (n_7_30), .A (n_3_32), .B (n_6_32), .C1 (n_5_29), .C2 (n_8_23) );
AOI211_X1 g_8_28 (.ZN (n_8_28), .A (n_5_31), .B (n_4_33), .C1 (n_4_31), .C2 (n_7_25) );
AOI211_X1 g_6_29 (.ZN (n_6_29), .A (n_7_30), .B (n_2_34), .C1 (n_6_32), .C2 (n_6_27) );
AOI211_X1 g_4_30 (.ZN (n_4_30), .A (n_8_28), .B (n_3_32), .C1 (n_4_33), .C2 (n_5_29) );
AOI211_X1 g_5_28 (.ZN (n_5_28), .A (n_6_29), .B (n_5_31), .C1 (n_2_34), .C2 (n_4_31) );
AOI211_X1 g_7_27 (.ZN (n_7_27), .A (n_4_30), .B (n_7_30), .C1 (n_3_32), .C2 (n_6_32) );
AOI211_X1 g_9_26 (.ZN (n_9_26), .A (n_5_28), .B (n_8_28), .C1 (n_5_31), .C2 (n_4_33) );
AOI211_X1 g_10_24 (.ZN (n_10_24), .A (n_7_27), .B (n_6_29), .C1 (n_7_30), .C2 (n_2_34) );
AOI211_X1 g_8_25 (.ZN (n_8_25), .A (n_9_26), .B (n_4_30), .C1 (n_8_28), .C2 (n_3_32) );
AOI211_X1 g_6_26 (.ZN (n_6_26), .A (n_10_24), .B (n_5_28), .C1 (n_6_29), .C2 (n_5_31) );
AOI211_X1 g_7_24 (.ZN (n_7_24), .A (n_8_25), .B (n_7_27), .C1 (n_4_30), .C2 (n_7_30) );
AOI211_X1 g_9_23 (.ZN (n_9_23), .A (n_6_26), .B (n_9_26), .C1 (n_5_28), .C2 (n_8_28) );
AOI211_X1 g_11_22 (.ZN (n_11_22), .A (n_7_24), .B (n_10_24), .C1 (n_7_27), .C2 (n_6_29) );
AOI211_X1 g_13_21 (.ZN (n_13_21), .A (n_9_23), .B (n_8_25), .C1 (n_9_26), .C2 (n_4_30) );
AOI211_X1 g_15_22 (.ZN (n_15_22), .A (n_11_22), .B (n_6_26), .C1 (n_10_24), .C2 (n_5_28) );
AOI211_X1 g_17_23 (.ZN (n_17_23), .A (n_13_21), .B (n_7_24), .C1 (n_8_25), .C2 (n_7_27) );
AOI211_X1 g_19_24 (.ZN (n_19_24), .A (n_15_22), .B (n_9_23), .C1 (n_6_26), .C2 (n_9_26) );
AOI211_X1 g_21_25 (.ZN (n_21_25), .A (n_17_23), .B (n_11_22), .C1 (n_7_24), .C2 (n_10_24) );
AOI211_X1 g_23_24 (.ZN (n_23_24), .A (n_19_24), .B (n_13_21), .C1 (n_9_23), .C2 (n_8_25) );
AOI211_X1 g_24_22 (.ZN (n_24_22), .A (n_21_25), .B (n_15_22), .C1 (n_11_22), .C2 (n_6_26) );
AOI211_X1 g_26_21 (.ZN (n_26_21), .A (n_23_24), .B (n_17_23), .C1 (n_13_21), .C2 (n_7_24) );
AOI211_X1 g_25_23 (.ZN (n_25_23), .A (n_24_22), .B (n_19_24), .C1 (n_15_22), .C2 (n_9_23) );
AOI211_X1 g_27_22 (.ZN (n_27_22), .A (n_26_21), .B (n_21_25), .C1 (n_17_23), .C2 (n_11_22) );
AOI211_X1 g_29_21 (.ZN (n_29_21), .A (n_25_23), .B (n_23_24), .C1 (n_19_24), .C2 (n_13_21) );
AOI211_X1 g_30_19 (.ZN (n_30_19), .A (n_27_22), .B (n_24_22), .C1 (n_21_25), .C2 (n_15_22) );
AOI211_X1 g_32_18 (.ZN (n_32_18), .A (n_29_21), .B (n_26_21), .C1 (n_23_24), .C2 (n_17_23) );
AOI211_X1 g_34_17 (.ZN (n_34_17), .A (n_30_19), .B (n_25_23), .C1 (n_24_22), .C2 (n_19_24) );
AOI211_X1 g_36_16 (.ZN (n_36_16), .A (n_32_18), .B (n_27_22), .C1 (n_26_21), .C2 (n_21_25) );
AOI211_X1 g_38_17 (.ZN (n_38_17), .A (n_34_17), .B (n_29_21), .C1 (n_25_23), .C2 (n_23_24) );
AOI211_X1 g_36_18 (.ZN (n_36_18), .A (n_36_16), .B (n_30_19), .C1 (n_27_22), .C2 (n_24_22) );
AOI211_X1 g_34_19 (.ZN (n_34_19), .A (n_38_17), .B (n_32_18), .C1 (n_29_21), .C2 (n_26_21) );
AOI211_X1 g_32_20 (.ZN (n_32_20), .A (n_36_18), .B (n_34_17), .C1 (n_30_19), .C2 (n_25_23) );
AOI211_X1 g_30_21 (.ZN (n_30_21), .A (n_34_19), .B (n_36_16), .C1 (n_32_18), .C2 (n_27_22) );
AOI211_X1 g_31_19 (.ZN (n_31_19), .A (n_32_20), .B (n_38_17), .C1 (n_34_17), .C2 (n_29_21) );
AOI211_X1 g_29_20 (.ZN (n_29_20), .A (n_30_21), .B (n_36_18), .C1 (n_36_16), .C2 (n_30_19) );
AOI211_X1 g_27_21 (.ZN (n_27_21), .A (n_31_19), .B (n_34_19), .C1 (n_38_17), .C2 (n_32_18) );
AOI211_X1 g_25_22 (.ZN (n_25_22), .A (n_29_20), .B (n_32_20), .C1 (n_36_18), .C2 (n_34_17) );
AOI211_X1 g_23_23 (.ZN (n_23_23), .A (n_27_21), .B (n_30_21), .C1 (n_34_19), .C2 (n_36_16) );
AOI211_X1 g_21_24 (.ZN (n_21_24), .A (n_25_22), .B (n_31_19), .C1 (n_32_20), .C2 (n_38_17) );
AOI211_X1 g_19_23 (.ZN (n_19_23), .A (n_23_23), .B (n_29_20), .C1 (n_30_21), .C2 (n_36_18) );
AOI211_X1 g_17_22 (.ZN (n_17_22), .A (n_21_24), .B (n_27_21), .C1 (n_31_19), .C2 (n_34_19) );
AOI211_X1 g_15_21 (.ZN (n_15_21), .A (n_19_23), .B (n_25_22), .C1 (n_29_20), .C2 (n_32_20) );
AOI211_X1 g_13_20 (.ZN (n_13_20), .A (n_17_22), .B (n_23_23), .C1 (n_27_21), .C2 (n_30_21) );
AOI211_X1 g_11_19 (.ZN (n_11_19), .A (n_15_21), .B (n_21_24), .C1 (n_25_22), .C2 (n_31_19) );
AOI211_X1 g_9_20 (.ZN (n_9_20), .A (n_13_20), .B (n_19_23), .C1 (n_23_23), .C2 (n_29_20) );
AOI211_X1 g_8_22 (.ZN (n_8_22), .A (n_11_19), .B (n_17_22), .C1 (n_21_24), .C2 (n_27_21) );
AOI211_X1 g_10_21 (.ZN (n_10_21), .A (n_9_20), .B (n_15_21), .C1 (n_19_23), .C2 (n_25_22) );
AOI211_X1 g_12_20 (.ZN (n_12_20), .A (n_8_22), .B (n_13_20), .C1 (n_17_22), .C2 (n_23_23) );
AOI211_X1 g_14_21 (.ZN (n_14_21), .A (n_10_21), .B (n_11_19), .C1 (n_15_21), .C2 (n_21_24) );
AOI211_X1 g_12_22 (.ZN (n_12_22), .A (n_12_20), .B (n_9_20), .C1 (n_13_20), .C2 (n_19_23) );
AOI211_X1 g_10_23 (.ZN (n_10_23), .A (n_14_21), .B (n_8_22), .C1 (n_11_19), .C2 (n_17_22) );
AOI211_X1 g_11_21 (.ZN (n_11_21), .A (n_12_22), .B (n_10_21), .C1 (n_9_20), .C2 (n_15_21) );
AOI211_X1 g_13_22 (.ZN (n_13_22), .A (n_10_23), .B (n_12_20), .C1 (n_8_22), .C2 (n_13_20) );
AOI211_X1 g_15_23 (.ZN (n_15_23), .A (n_11_21), .B (n_14_21), .C1 (n_10_21), .C2 (n_11_19) );
AOI211_X1 g_17_24 (.ZN (n_17_24), .A (n_13_22), .B (n_12_22), .C1 (n_12_20), .C2 (n_9_20) );
AOI211_X1 g_16_22 (.ZN (n_16_22), .A (n_15_23), .B (n_10_23), .C1 (n_14_21), .C2 (n_8_22) );
AOI211_X1 g_14_23 (.ZN (n_14_23), .A (n_17_24), .B (n_11_21), .C1 (n_12_22), .C2 (n_10_21) );
AOI211_X1 g_12_24 (.ZN (n_12_24), .A (n_16_22), .B (n_13_22), .C1 (n_10_23), .C2 (n_12_20) );
AOI211_X1 g_10_25 (.ZN (n_10_25), .A (n_14_23), .B (n_15_23), .C1 (n_11_21), .C2 (n_14_21) );
AOI211_X1 g_11_23 (.ZN (n_11_23), .A (n_12_24), .B (n_17_24), .C1 (n_13_22), .C2 (n_12_22) );
AOI211_X1 g_12_21 (.ZN (n_12_21), .A (n_10_25), .B (n_16_22), .C1 (n_15_23), .C2 (n_10_23) );
AOI211_X1 g_10_22 (.ZN (n_10_22), .A (n_11_23), .B (n_14_23), .C1 (n_17_24), .C2 (n_11_21) );
AOI211_X1 g_9_24 (.ZN (n_9_24), .A (n_12_21), .B (n_12_24), .C1 (n_16_22), .C2 (n_13_22) );
AOI211_X1 g_8_26 (.ZN (n_8_26), .A (n_10_22), .B (n_10_25), .C1 (n_14_23), .C2 (n_15_23) );
AOI211_X1 g_7_28 (.ZN (n_7_28), .A (n_9_24), .B (n_11_23), .C1 (n_12_24), .C2 (n_17_24) );
AOI211_X1 g_9_27 (.ZN (n_9_27), .A (n_8_26), .B (n_12_21), .C1 (n_10_25), .C2 (n_16_22) );
AOI211_X1 g_11_26 (.ZN (n_11_26), .A (n_7_28), .B (n_10_22), .C1 (n_11_23), .C2 (n_14_23) );
AOI211_X1 g_9_25 (.ZN (n_9_25), .A (n_9_27), .B (n_9_24), .C1 (n_12_21), .C2 (n_12_24) );
AOI211_X1 g_11_24 (.ZN (n_11_24), .A (n_11_26), .B (n_8_26), .C1 (n_10_22), .C2 (n_10_25) );
AOI211_X1 g_13_23 (.ZN (n_13_23), .A (n_9_25), .B (n_7_28), .C1 (n_9_24), .C2 (n_11_23) );
AOI211_X1 g_12_25 (.ZN (n_12_25), .A (n_11_24), .B (n_9_27), .C1 (n_8_26), .C2 (n_12_21) );
AOI211_X1 g_10_26 (.ZN (n_10_26), .A (n_13_23), .B (n_11_26), .C1 (n_7_28), .C2 (n_10_22) );
AOI211_X1 g_8_27 (.ZN (n_8_27), .A (n_12_25), .B (n_9_25), .C1 (n_9_27), .C2 (n_9_24) );
AOI211_X1 g_7_29 (.ZN (n_7_29), .A (n_10_26), .B (n_11_24), .C1 (n_11_26), .C2 (n_8_26) );
AOI211_X1 g_9_28 (.ZN (n_9_28), .A (n_8_27), .B (n_13_23), .C1 (n_9_25), .C2 (n_7_28) );
AOI211_X1 g_11_27 (.ZN (n_11_27), .A (n_7_29), .B (n_12_25), .C1 (n_11_24), .C2 (n_9_27) );
AOI211_X1 g_10_29 (.ZN (n_10_29), .A (n_9_28), .B (n_10_26), .C1 (n_13_23), .C2 (n_11_26) );
AOI211_X1 g_8_30 (.ZN (n_8_30), .A (n_11_27), .B (n_8_27), .C1 (n_12_25), .C2 (n_9_25) );
AOI211_X1 g_6_31 (.ZN (n_6_31), .A (n_10_29), .B (n_7_29), .C1 (n_10_26), .C2 (n_11_24) );
AOI211_X1 g_5_33 (.ZN (n_5_33), .A (n_8_30), .B (n_9_28), .C1 (n_8_27), .C2 (n_13_23) );
AOI211_X1 g_4_35 (.ZN (n_4_35), .A (n_6_31), .B (n_11_27), .C1 (n_7_29), .C2 (n_12_25) );
AOI211_X1 g_6_36 (.ZN (n_6_36), .A (n_5_33), .B (n_10_29), .C1 (n_9_28), .C2 (n_10_26) );
AOI211_X1 g_4_37 (.ZN (n_4_37), .A (n_4_35), .B (n_8_30), .C1 (n_11_27), .C2 (n_8_27) );
AOI211_X1 g_2_38 (.ZN (n_2_38), .A (n_6_36), .B (n_6_31), .C1 (n_10_29), .C2 (n_7_29) );
AOI211_X1 g_3_36 (.ZN (n_3_36), .A (n_4_37), .B (n_5_33), .C1 (n_8_30), .C2 (n_9_28) );
AOI211_X1 g_5_35 (.ZN (n_5_35), .A (n_2_38), .B (n_4_35), .C1 (n_6_31), .C2 (n_11_27) );
AOI211_X1 g_7_34 (.ZN (n_7_34), .A (n_3_36), .B (n_6_36), .C1 (n_5_33), .C2 (n_10_29) );
AOI211_X1 g_8_32 (.ZN (n_8_32), .A (n_5_35), .B (n_4_37), .C1 (n_4_35), .C2 (n_8_30) );
AOI211_X1 g_6_33 (.ZN (n_6_33), .A (n_7_34), .B (n_2_38), .C1 (n_6_36), .C2 (n_6_31) );
AOI211_X1 g_4_34 (.ZN (n_4_34), .A (n_8_32), .B (n_3_36), .C1 (n_4_37), .C2 (n_5_33) );
AOI211_X1 g_5_32 (.ZN (n_5_32), .A (n_6_33), .B (n_5_35), .C1 (n_2_38), .C2 (n_4_35) );
AOI211_X1 g_6_30 (.ZN (n_6_30), .A (n_4_34), .B (n_7_34), .C1 (n_3_36), .C2 (n_6_36) );
AOI211_X1 g_8_29 (.ZN (n_8_29), .A (n_5_32), .B (n_8_32), .C1 (n_5_35), .C2 (n_4_37) );
AOI211_X1 g_7_31 (.ZN (n_7_31), .A (n_6_30), .B (n_6_33), .C1 (n_7_34), .C2 (n_2_38) );
AOI211_X1 g_9_30 (.ZN (n_9_30), .A (n_8_29), .B (n_4_34), .C1 (n_8_32), .C2 (n_3_36) );
AOI211_X1 g_10_28 (.ZN (n_10_28), .A (n_7_31), .B (n_5_32), .C1 (n_6_33), .C2 (n_5_35) );
AOI211_X1 g_12_27 (.ZN (n_12_27), .A (n_9_30), .B (n_6_30), .C1 (n_4_34), .C2 (n_7_34) );
AOI211_X1 g_13_25 (.ZN (n_13_25), .A (n_10_28), .B (n_8_29), .C1 (n_5_32), .C2 (n_8_32) );
AOI211_X1 g_12_23 (.ZN (n_12_23), .A (n_12_27), .B (n_7_31), .C1 (n_6_30), .C2 (n_6_33) );
AOI211_X1 g_14_22 (.ZN (n_14_22), .A (n_13_25), .B (n_9_30), .C1 (n_8_29), .C2 (n_4_34) );
AOI211_X1 g_15_24 (.ZN (n_15_24), .A (n_12_23), .B (n_10_28), .C1 (n_7_31), .C2 (n_5_32) );
AOI211_X1 g_14_26 (.ZN (n_14_26), .A (n_14_22), .B (n_12_27), .C1 (n_9_30), .C2 (n_6_30) );
AOI211_X1 g_13_24 (.ZN (n_13_24), .A (n_15_24), .B (n_13_25), .C1 (n_10_28), .C2 (n_8_29) );
AOI211_X1 g_11_25 (.ZN (n_11_25), .A (n_14_26), .B (n_12_23), .C1 (n_12_27), .C2 (n_7_31) );
AOI211_X1 g_10_27 (.ZN (n_10_27), .A (n_13_24), .B (n_14_22), .C1 (n_13_25), .C2 (n_9_30) );
AOI211_X1 g_12_26 (.ZN (n_12_26), .A (n_11_25), .B (n_15_24), .C1 (n_12_23), .C2 (n_10_28) );
AOI211_X1 g_14_25 (.ZN (n_14_25), .A (n_10_27), .B (n_14_26), .C1 (n_14_22), .C2 (n_12_27) );
AOI211_X1 g_16_24 (.ZN (n_16_24), .A (n_12_26), .B (n_13_24), .C1 (n_15_24), .C2 (n_13_25) );
AOI211_X1 g_18_23 (.ZN (n_18_23), .A (n_14_25), .B (n_11_25), .C1 (n_14_26), .C2 (n_12_23) );
AOI211_X1 g_19_25 (.ZN (n_19_25), .A (n_16_24), .B (n_10_27), .C1 (n_13_24), .C2 (n_14_22) );
AOI211_X1 g_17_26 (.ZN (n_17_26), .A (n_18_23), .B (n_12_26), .C1 (n_11_25), .C2 (n_15_24) );
AOI211_X1 g_18_24 (.ZN (n_18_24), .A (n_19_25), .B (n_14_25), .C1 (n_10_27), .C2 (n_14_26) );
AOI211_X1 g_16_23 (.ZN (n_16_23), .A (n_17_26), .B (n_16_24), .C1 (n_12_26), .C2 (n_13_24) );
AOI211_X1 g_14_24 (.ZN (n_14_24), .A (n_18_24), .B (n_18_23), .C1 (n_14_25), .C2 (n_11_25) );
AOI211_X1 g_16_25 (.ZN (n_16_25), .A (n_16_23), .B (n_19_25), .C1 (n_16_24), .C2 (n_10_27) );
AOI211_X1 g_15_27 (.ZN (n_15_27), .A (n_14_24), .B (n_17_26), .C1 (n_18_23), .C2 (n_12_26) );
AOI211_X1 g_13_26 (.ZN (n_13_26), .A (n_16_25), .B (n_18_24), .C1 (n_19_25), .C2 (n_14_25) );
AOI211_X1 g_15_25 (.ZN (n_15_25), .A (n_15_27), .B (n_16_23), .C1 (n_17_26), .C2 (n_16_24) );
AOI211_X1 g_14_27 (.ZN (n_14_27), .A (n_13_26), .B (n_14_24), .C1 (n_18_24), .C2 (n_18_23) );
AOI211_X1 g_12_28 (.ZN (n_12_28), .A (n_15_25), .B (n_16_25), .C1 (n_16_23), .C2 (n_19_25) );
AOI211_X1 g_11_30 (.ZN (n_11_30), .A (n_14_27), .B (n_15_27), .C1 (n_14_24), .C2 (n_17_26) );
AOI211_X1 g_9_29 (.ZN (n_9_29), .A (n_12_28), .B (n_13_26), .C1 (n_16_25), .C2 (n_18_24) );
AOI211_X1 g_11_28 (.ZN (n_11_28), .A (n_11_30), .B (n_15_25), .C1 (n_15_27), .C2 (n_16_23) );
AOI211_X1 g_13_27 (.ZN (n_13_27), .A (n_9_29), .B (n_14_27), .C1 (n_13_26), .C2 (n_14_24) );
AOI211_X1 g_15_26 (.ZN (n_15_26), .A (n_11_28), .B (n_12_28), .C1 (n_15_25), .C2 (n_16_25) );
AOI211_X1 g_17_25 (.ZN (n_17_25), .A (n_13_27), .B (n_11_30), .C1 (n_14_27), .C2 (n_15_27) );
AOI211_X1 g_16_27 (.ZN (n_16_27), .A (n_15_26), .B (n_9_29), .C1 (n_12_28), .C2 (n_13_26) );
AOI211_X1 g_18_26 (.ZN (n_18_26), .A (n_17_25), .B (n_11_28), .C1 (n_11_30), .C2 (n_15_25) );
AOI211_X1 g_20_25 (.ZN (n_20_25), .A (n_16_27), .B (n_13_27), .C1 (n_9_29), .C2 (n_14_27) );
AOI211_X1 g_22_24 (.ZN (n_22_24), .A (n_18_26), .B (n_15_26), .C1 (n_11_28), .C2 (n_12_28) );
AOI211_X1 g_24_23 (.ZN (n_24_23), .A (n_20_25), .B (n_17_25), .C1 (n_13_27), .C2 (n_11_30) );
AOI211_X1 g_26_22 (.ZN (n_26_22), .A (n_22_24), .B (n_16_27), .C1 (n_15_26), .C2 (n_9_29) );
AOI211_X1 g_28_21 (.ZN (n_28_21), .A (n_24_23), .B (n_18_26), .C1 (n_17_25), .C2 (n_11_28) );
AOI211_X1 g_30_20 (.ZN (n_30_20), .A (n_26_22), .B (n_20_25), .C1 (n_16_27), .C2 (n_13_27) );
AOI211_X1 g_32_19 (.ZN (n_32_19), .A (n_28_21), .B (n_22_24), .C1 (n_18_26), .C2 (n_15_26) );
AOI211_X1 g_31_21 (.ZN (n_31_21), .A (n_30_20), .B (n_24_23), .C1 (n_20_25), .C2 (n_17_25) );
AOI211_X1 g_33_20 (.ZN (n_33_20), .A (n_32_19), .B (n_26_22), .C1 (n_22_24), .C2 (n_16_27) );
AOI211_X1 g_35_19 (.ZN (n_35_19), .A (n_31_21), .B (n_28_21), .C1 (n_24_23), .C2 (n_18_26) );
AOI211_X1 g_37_18 (.ZN (n_37_18), .A (n_33_20), .B (n_30_20), .C1 (n_26_22), .C2 (n_20_25) );
AOI211_X1 g_39_17 (.ZN (n_39_17), .A (n_35_19), .B (n_32_19), .C1 (n_28_21), .C2 (n_22_24) );
AOI211_X1 g_41_16 (.ZN (n_41_16), .A (n_37_18), .B (n_31_21), .C1 (n_30_20), .C2 (n_24_23) );
AOI211_X1 g_43_15 (.ZN (n_43_15), .A (n_39_17), .B (n_33_20), .C1 (n_32_19), .C2 (n_26_22) );
AOI211_X1 g_45_14 (.ZN (n_45_14), .A (n_41_16), .B (n_35_19), .C1 (n_31_21), .C2 (n_28_21) );
AOI211_X1 g_47_13 (.ZN (n_47_13), .A (n_43_15), .B (n_37_18), .C1 (n_33_20), .C2 (n_30_20) );
AOI211_X1 g_46_15 (.ZN (n_46_15), .A (n_45_14), .B (n_39_17), .C1 (n_35_19), .C2 (n_32_19) );
AOI211_X1 g_48_14 (.ZN (n_48_14), .A (n_47_13), .B (n_41_16), .C1 (n_37_18), .C2 (n_31_21) );
AOI211_X1 g_50_13 (.ZN (n_50_13), .A (n_46_15), .B (n_43_15), .C1 (n_39_17), .C2 (n_33_20) );
AOI211_X1 g_52_12 (.ZN (n_52_12), .A (n_48_14), .B (n_45_14), .C1 (n_41_16), .C2 (n_35_19) );
AOI211_X1 g_54_11 (.ZN (n_54_11), .A (n_50_13), .B (n_47_13), .C1 (n_43_15), .C2 (n_37_18) );
AOI211_X1 g_56_10 (.ZN (n_56_10), .A (n_52_12), .B (n_46_15), .C1 (n_45_14), .C2 (n_39_17) );
AOI211_X1 g_58_9 (.ZN (n_58_9), .A (n_54_11), .B (n_48_14), .C1 (n_47_13), .C2 (n_41_16) );
AOI211_X1 g_57_11 (.ZN (n_57_11), .A (n_56_10), .B (n_50_13), .C1 (n_46_15), .C2 (n_43_15) );
AOI211_X1 g_59_10 (.ZN (n_59_10), .A (n_58_9), .B (n_52_12), .C1 (n_48_14), .C2 (n_45_14) );
AOI211_X1 g_61_9 (.ZN (n_61_9), .A (n_57_11), .B (n_54_11), .C1 (n_50_13), .C2 (n_47_13) );
AOI211_X1 g_63_8 (.ZN (n_63_8), .A (n_59_10), .B (n_56_10), .C1 (n_52_12), .C2 (n_46_15) );
AOI211_X1 g_65_7 (.ZN (n_65_7), .A (n_61_9), .B (n_58_9), .C1 (n_54_11), .C2 (n_48_14) );
AOI211_X1 g_67_6 (.ZN (n_67_6), .A (n_63_8), .B (n_57_11), .C1 (n_56_10), .C2 (n_50_13) );
AOI211_X1 g_69_5 (.ZN (n_69_5), .A (n_65_7), .B (n_59_10), .C1 (n_58_9), .C2 (n_52_12) );
AOI211_X1 g_71_4 (.ZN (n_71_4), .A (n_67_6), .B (n_61_9), .C1 (n_57_11), .C2 (n_54_11) );
AOI211_X1 g_73_3 (.ZN (n_73_3), .A (n_69_5), .B (n_63_8), .C1 (n_59_10), .C2 (n_56_10) );
AOI211_X1 g_75_2 (.ZN (n_75_2), .A (n_71_4), .B (n_65_7), .C1 (n_61_9), .C2 (n_58_9) );
AOI211_X1 g_77_1 (.ZN (n_77_1), .A (n_73_3), .B (n_67_6), .C1 (n_63_8), .C2 (n_57_11) );
AOI211_X1 g_76_3 (.ZN (n_76_3), .A (n_75_2), .B (n_69_5), .C1 (n_65_7), .C2 (n_59_10) );
AOI211_X1 g_78_2 (.ZN (n_78_2), .A (n_77_1), .B (n_71_4), .C1 (n_67_6), .C2 (n_61_9) );
AOI211_X1 g_80_1 (.ZN (n_80_1), .A (n_76_3), .B (n_73_3), .C1 (n_69_5), .C2 (n_63_8) );
AOI211_X1 g_79_3 (.ZN (n_79_3), .A (n_78_2), .B (n_75_2), .C1 (n_71_4), .C2 (n_65_7) );
AOI211_X1 g_78_1 (.ZN (n_78_1), .A (n_80_1), .B (n_77_1), .C1 (n_73_3), .C2 (n_67_6) );
AOI211_X1 g_76_2 (.ZN (n_76_2), .A (n_79_3), .B (n_76_3), .C1 (n_75_2), .C2 (n_69_5) );
AOI211_X1 g_74_3 (.ZN (n_74_3), .A (n_78_1), .B (n_78_2), .C1 (n_77_1), .C2 (n_71_4) );
AOI211_X1 g_72_4 (.ZN (n_72_4), .A (n_76_2), .B (n_80_1), .C1 (n_76_3), .C2 (n_73_3) );
AOI211_X1 g_70_5 (.ZN (n_70_5), .A (n_74_3), .B (n_79_3), .C1 (n_78_2), .C2 (n_75_2) );
AOI211_X1 g_68_6 (.ZN (n_68_6), .A (n_72_4), .B (n_78_1), .C1 (n_80_1), .C2 (n_77_1) );
AOI211_X1 g_66_7 (.ZN (n_66_7), .A (n_70_5), .B (n_76_2), .C1 (n_79_3), .C2 (n_76_3) );
AOI211_X1 g_64_8 (.ZN (n_64_8), .A (n_68_6), .B (n_74_3), .C1 (n_78_1), .C2 (n_78_2) );
AOI211_X1 g_62_9 (.ZN (n_62_9), .A (n_66_7), .B (n_72_4), .C1 (n_76_2), .C2 (n_80_1) );
AOI211_X1 g_63_7 (.ZN (n_63_7), .A (n_64_8), .B (n_70_5), .C1 (n_74_3), .C2 (n_79_3) );
AOI211_X1 g_61_8 (.ZN (n_61_8), .A (n_62_9), .B (n_68_6), .C1 (n_72_4), .C2 (n_78_1) );
AOI211_X1 g_59_9 (.ZN (n_59_9), .A (n_63_7), .B (n_66_7), .C1 (n_70_5), .C2 (n_76_2) );
AOI211_X1 g_57_10 (.ZN (n_57_10), .A (n_61_8), .B (n_64_8), .C1 (n_68_6), .C2 (n_74_3) );
AOI211_X1 g_55_11 (.ZN (n_55_11), .A (n_59_9), .B (n_62_9), .C1 (n_66_7), .C2 (n_72_4) );
AOI211_X1 g_53_12 (.ZN (n_53_12), .A (n_57_10), .B (n_63_7), .C1 (n_64_8), .C2 (n_70_5) );
AOI211_X1 g_51_13 (.ZN (n_51_13), .A (n_55_11), .B (n_61_8), .C1 (n_62_9), .C2 (n_68_6) );
AOI211_X1 g_49_14 (.ZN (n_49_14), .A (n_53_12), .B (n_59_9), .C1 (n_63_7), .C2 (n_66_7) );
AOI211_X1 g_47_15 (.ZN (n_47_15), .A (n_51_13), .B (n_57_10), .C1 (n_61_8), .C2 (n_64_8) );
AOI211_X1 g_45_16 (.ZN (n_45_16), .A (n_49_14), .B (n_55_11), .C1 (n_59_9), .C2 (n_62_9) );
AOI211_X1 g_43_17 (.ZN (n_43_17), .A (n_47_15), .B (n_53_12), .C1 (n_57_10), .C2 (n_63_7) );
AOI211_X1 g_44_15 (.ZN (n_44_15), .A (n_45_16), .B (n_51_13), .C1 (n_55_11), .C2 (n_61_8) );
AOI211_X1 g_42_16 (.ZN (n_42_16), .A (n_43_17), .B (n_49_14), .C1 (n_53_12), .C2 (n_59_9) );
AOI211_X1 g_43_14 (.ZN (n_43_14), .A (n_44_15), .B (n_47_15), .C1 (n_51_13), .C2 (n_57_10) );
AOI211_X1 g_41_15 (.ZN (n_41_15), .A (n_42_16), .B (n_45_16), .C1 (n_49_14), .C2 (n_55_11) );
AOI211_X1 g_39_16 (.ZN (n_39_16), .A (n_43_14), .B (n_43_17), .C1 (n_47_15), .C2 (n_53_12) );
AOI211_X1 g_37_17 (.ZN (n_37_17), .A (n_41_15), .B (n_44_15), .C1 (n_45_16), .C2 (n_51_13) );
AOI211_X1 g_35_18 (.ZN (n_35_18), .A (n_39_16), .B (n_42_16), .C1 (n_43_17), .C2 (n_49_14) );
AOI211_X1 g_33_19 (.ZN (n_33_19), .A (n_37_17), .B (n_43_14), .C1 (n_44_15), .C2 (n_47_15) );
AOI211_X1 g_31_20 (.ZN (n_31_20), .A (n_35_18), .B (n_41_15), .C1 (n_42_16), .C2 (n_45_16) );
AOI211_X1 g_30_22 (.ZN (n_30_22), .A (n_33_19), .B (n_39_16), .C1 (n_43_14), .C2 (n_43_17) );
AOI211_X1 g_32_21 (.ZN (n_32_21), .A (n_31_20), .B (n_37_17), .C1 (n_41_15), .C2 (n_44_15) );
AOI211_X1 g_34_20 (.ZN (n_34_20), .A (n_30_22), .B (n_35_18), .C1 (n_39_16), .C2 (n_42_16) );
AOI211_X1 g_36_19 (.ZN (n_36_19), .A (n_32_21), .B (n_33_19), .C1 (n_37_17), .C2 (n_43_14) );
AOI211_X1 g_38_18 (.ZN (n_38_18), .A (n_34_20), .B (n_31_20), .C1 (n_35_18), .C2 (n_41_15) );
AOI211_X1 g_40_17 (.ZN (n_40_17), .A (n_36_19), .B (n_30_22), .C1 (n_33_19), .C2 (n_39_16) );
AOI211_X1 g_39_19 (.ZN (n_39_19), .A (n_38_18), .B (n_32_21), .C1 (n_31_20), .C2 (n_37_17) );
AOI211_X1 g_41_18 (.ZN (n_41_18), .A (n_40_17), .B (n_34_20), .C1 (n_30_22), .C2 (n_35_18) );
AOI211_X1 g_40_20 (.ZN (n_40_20), .A (n_39_19), .B (n_36_19), .C1 (n_32_21), .C2 (n_33_19) );
AOI211_X1 g_39_18 (.ZN (n_39_18), .A (n_41_18), .B (n_38_18), .C1 (n_34_20), .C2 (n_31_20) );
AOI211_X1 g_41_17 (.ZN (n_41_17), .A (n_40_20), .B (n_40_17), .C1 (n_36_19), .C2 (n_30_22) );
AOI211_X1 g_43_16 (.ZN (n_43_16), .A (n_39_18), .B (n_39_19), .C1 (n_38_18), .C2 (n_32_21) );
AOI211_X1 g_45_15 (.ZN (n_45_15), .A (n_41_17), .B (n_41_18), .C1 (n_40_17), .C2 (n_34_20) );
AOI211_X1 g_47_14 (.ZN (n_47_14), .A (n_43_16), .B (n_40_20), .C1 (n_39_19), .C2 (n_36_19) );
AOI211_X1 g_49_13 (.ZN (n_49_13), .A (n_45_15), .B (n_39_18), .C1 (n_41_18), .C2 (n_38_18) );
AOI211_X1 g_48_15 (.ZN (n_48_15), .A (n_47_14), .B (n_41_17), .C1 (n_40_20), .C2 (n_40_17) );
AOI211_X1 g_46_16 (.ZN (n_46_16), .A (n_49_13), .B (n_43_16), .C1 (n_39_18), .C2 (n_39_19) );
AOI211_X1 g_44_17 (.ZN (n_44_17), .A (n_48_15), .B (n_45_15), .C1 (n_41_17), .C2 (n_41_18) );
AOI211_X1 g_42_18 (.ZN (n_42_18), .A (n_46_16), .B (n_47_14), .C1 (n_43_16), .C2 (n_40_20) );
AOI211_X1 g_40_19 (.ZN (n_40_19), .A (n_44_17), .B (n_49_13), .C1 (n_45_15), .C2 (n_39_18) );
AOI211_X1 g_38_20 (.ZN (n_38_20), .A (n_42_18), .B (n_48_15), .C1 (n_47_14), .C2 (n_41_17) );
AOI211_X1 g_36_21 (.ZN (n_36_21), .A (n_40_19), .B (n_46_16), .C1 (n_49_13), .C2 (n_43_16) );
AOI211_X1 g_37_19 (.ZN (n_37_19), .A (n_38_20), .B (n_44_17), .C1 (n_48_15), .C2 (n_45_15) );
AOI211_X1 g_35_20 (.ZN (n_35_20), .A (n_36_21), .B (n_42_18), .C1 (n_46_16), .C2 (n_47_14) );
AOI211_X1 g_33_21 (.ZN (n_33_21), .A (n_37_19), .B (n_40_19), .C1 (n_44_17), .C2 (n_49_13) );
AOI211_X1 g_31_22 (.ZN (n_31_22), .A (n_35_20), .B (n_38_20), .C1 (n_42_18), .C2 (n_48_15) );
AOI211_X1 g_29_23 (.ZN (n_29_23), .A (n_33_21), .B (n_36_21), .C1 (n_40_19), .C2 (n_46_16) );
AOI211_X1 g_27_24 (.ZN (n_27_24), .A (n_31_22), .B (n_37_19), .C1 (n_38_20), .C2 (n_44_17) );
AOI211_X1 g_28_22 (.ZN (n_28_22), .A (n_29_23), .B (n_35_20), .C1 (n_36_21), .C2 (n_42_18) );
AOI211_X1 g_26_23 (.ZN (n_26_23), .A (n_27_24), .B (n_33_21), .C1 (n_37_19), .C2 (n_40_19) );
AOI211_X1 g_24_24 (.ZN (n_24_24), .A (n_28_22), .B (n_31_22), .C1 (n_35_20), .C2 (n_38_20) );
AOI211_X1 g_22_25 (.ZN (n_22_25), .A (n_26_23), .B (n_29_23), .C1 (n_33_21), .C2 (n_36_21) );
AOI211_X1 g_20_24 (.ZN (n_20_24), .A (n_24_24), .B (n_27_24), .C1 (n_31_22), .C2 (n_37_19) );
AOI211_X1 g_18_25 (.ZN (n_18_25), .A (n_22_25), .B (n_28_22), .C1 (n_29_23), .C2 (n_35_20) );
AOI211_X1 g_16_26 (.ZN (n_16_26), .A (n_20_24), .B (n_26_23), .C1 (n_27_24), .C2 (n_33_21) );
AOI211_X1 g_15_28 (.ZN (n_15_28), .A (n_18_25), .B (n_24_24), .C1 (n_28_22), .C2 (n_31_22) );
AOI211_X1 g_13_29 (.ZN (n_13_29), .A (n_16_26), .B (n_22_25), .C1 (n_26_23), .C2 (n_29_23) );
AOI211_X1 g_12_31 (.ZN (n_12_31), .A (n_15_28), .B (n_20_24), .C1 (n_24_24), .C2 (n_27_24) );
AOI211_X1 g_11_29 (.ZN (n_11_29), .A (n_13_29), .B (n_18_25), .C1 (n_22_25), .C2 (n_28_22) );
AOI211_X1 g_13_28 (.ZN (n_13_28), .A (n_12_31), .B (n_16_26), .C1 (n_20_24), .C2 (n_26_23) );
AOI211_X1 g_12_30 (.ZN (n_12_30), .A (n_11_29), .B (n_15_28), .C1 (n_18_25), .C2 (n_24_24) );
AOI211_X1 g_10_31 (.ZN (n_10_31), .A (n_13_28), .B (n_13_29), .C1 (n_16_26), .C2 (n_22_25) );
AOI211_X1 g_9_33 (.ZN (n_9_33), .A (n_12_30), .B (n_12_31), .C1 (n_15_28), .C2 (n_20_24) );
AOI211_X1 g_8_31 (.ZN (n_8_31), .A (n_10_31), .B (n_11_29), .C1 (n_13_29), .C2 (n_18_25) );
AOI211_X1 g_10_30 (.ZN (n_10_30), .A (n_9_33), .B (n_13_28), .C1 (n_12_31), .C2 (n_16_26) );
AOI211_X1 g_12_29 (.ZN (n_12_29), .A (n_8_31), .B (n_12_30), .C1 (n_11_29), .C2 (n_15_28) );
AOI211_X1 g_14_28 (.ZN (n_14_28), .A (n_10_30), .B (n_10_31), .C1 (n_13_28), .C2 (n_13_29) );
AOI211_X1 g_13_30 (.ZN (n_13_30), .A (n_12_29), .B (n_9_33), .C1 (n_12_30), .C2 (n_12_31) );
AOI211_X1 g_15_29 (.ZN (n_15_29), .A (n_14_28), .B (n_8_31), .C1 (n_10_31), .C2 (n_11_29) );
AOI211_X1 g_17_28 (.ZN (n_17_28), .A (n_13_30), .B (n_10_30), .C1 (n_9_33), .C2 (n_13_28) );
AOI211_X1 g_19_27 (.ZN (n_19_27), .A (n_15_29), .B (n_12_29), .C1 (n_8_31), .C2 (n_12_30) );
AOI211_X1 g_21_26 (.ZN (n_21_26), .A (n_17_28), .B (n_14_28), .C1 (n_10_30), .C2 (n_10_31) );
AOI211_X1 g_23_25 (.ZN (n_23_25), .A (n_19_27), .B (n_13_30), .C1 (n_12_29), .C2 (n_9_33) );
AOI211_X1 g_25_24 (.ZN (n_25_24), .A (n_21_26), .B (n_15_29), .C1 (n_14_28), .C2 (n_8_31) );
AOI211_X1 g_27_23 (.ZN (n_27_23), .A (n_23_25), .B (n_17_28), .C1 (n_13_30), .C2 (n_10_30) );
AOI211_X1 g_29_22 (.ZN (n_29_22), .A (n_25_24), .B (n_19_27), .C1 (n_15_29), .C2 (n_12_29) );
AOI211_X1 g_28_24 (.ZN (n_28_24), .A (n_27_23), .B (n_21_26), .C1 (n_17_28), .C2 (n_14_28) );
AOI211_X1 g_30_23 (.ZN (n_30_23), .A (n_29_22), .B (n_23_25), .C1 (n_19_27), .C2 (n_13_30) );
AOI211_X1 g_32_22 (.ZN (n_32_22), .A (n_28_24), .B (n_25_24), .C1 (n_21_26), .C2 (n_15_29) );
AOI211_X1 g_34_21 (.ZN (n_34_21), .A (n_30_23), .B (n_27_23), .C1 (n_23_25), .C2 (n_17_28) );
AOI211_X1 g_36_20 (.ZN (n_36_20), .A (n_32_22), .B (n_29_22), .C1 (n_25_24), .C2 (n_19_27) );
AOI211_X1 g_38_19 (.ZN (n_38_19), .A (n_34_21), .B (n_28_24), .C1 (n_27_23), .C2 (n_21_26) );
AOI211_X1 g_40_18 (.ZN (n_40_18), .A (n_36_20), .B (n_30_23), .C1 (n_29_22), .C2 (n_23_25) );
AOI211_X1 g_42_17 (.ZN (n_42_17), .A (n_38_19), .B (n_32_22), .C1 (n_28_24), .C2 (n_25_24) );
AOI211_X1 g_44_16 (.ZN (n_44_16), .A (n_40_18), .B (n_34_21), .C1 (n_30_23), .C2 (n_27_23) );
AOI211_X1 g_43_18 (.ZN (n_43_18), .A (n_42_17), .B (n_36_20), .C1 (n_32_22), .C2 (n_29_22) );
AOI211_X1 g_45_17 (.ZN (n_45_17), .A (n_44_16), .B (n_38_19), .C1 (n_34_21), .C2 (n_28_24) );
AOI211_X1 g_47_16 (.ZN (n_47_16), .A (n_43_18), .B (n_40_18), .C1 (n_36_20), .C2 (n_30_23) );
AOI211_X1 g_49_15 (.ZN (n_49_15), .A (n_45_17), .B (n_42_17), .C1 (n_38_19), .C2 (n_32_22) );
AOI211_X1 g_51_14 (.ZN (n_51_14), .A (n_47_16), .B (n_44_16), .C1 (n_40_18), .C2 (n_34_21) );
AOI211_X1 g_53_13 (.ZN (n_53_13), .A (n_49_15), .B (n_43_18), .C1 (n_42_17), .C2 (n_36_20) );
AOI211_X1 g_55_12 (.ZN (n_55_12), .A (n_51_14), .B (n_45_17), .C1 (n_44_16), .C2 (n_38_19) );
AOI211_X1 g_54_14 (.ZN (n_54_14), .A (n_53_13), .B (n_47_16), .C1 (n_43_18), .C2 (n_40_18) );
AOI211_X1 g_56_13 (.ZN (n_56_13), .A (n_55_12), .B (n_49_15), .C1 (n_45_17), .C2 (n_42_17) );
AOI211_X1 g_58_12 (.ZN (n_58_12), .A (n_54_14), .B (n_51_14), .C1 (n_47_16), .C2 (n_44_16) );
AOI211_X1 g_60_11 (.ZN (n_60_11), .A (n_56_13), .B (n_53_13), .C1 (n_49_15), .C2 (n_43_18) );
AOI211_X1 g_62_10 (.ZN (n_62_10), .A (n_58_12), .B (n_55_12), .C1 (n_51_14), .C2 (n_45_17) );
AOI211_X1 g_64_9 (.ZN (n_64_9), .A (n_60_11), .B (n_54_14), .C1 (n_53_13), .C2 (n_47_16) );
AOI211_X1 g_66_8 (.ZN (n_66_8), .A (n_62_10), .B (n_56_13), .C1 (n_55_12), .C2 (n_49_15) );
AOI211_X1 g_68_7 (.ZN (n_68_7), .A (n_64_9), .B (n_58_12), .C1 (n_54_14), .C2 (n_51_14) );
AOI211_X1 g_70_6 (.ZN (n_70_6), .A (n_66_8), .B (n_60_11), .C1 (n_56_13), .C2 (n_53_13) );
AOI211_X1 g_72_5 (.ZN (n_72_5), .A (n_68_7), .B (n_62_10), .C1 (n_58_12), .C2 (n_55_12) );
AOI211_X1 g_74_4 (.ZN (n_74_4), .A (n_70_6), .B (n_64_9), .C1 (n_60_11), .C2 (n_54_14) );
AOI211_X1 g_73_6 (.ZN (n_73_6), .A (n_72_5), .B (n_66_8), .C1 (n_62_10), .C2 (n_56_13) );
AOI211_X1 g_75_5 (.ZN (n_75_5), .A (n_74_4), .B (n_68_7), .C1 (n_64_9), .C2 (n_58_12) );
AOI211_X1 g_77_4 (.ZN (n_77_4), .A (n_73_6), .B (n_70_6), .C1 (n_66_8), .C2 (n_60_11) );
AOI211_X1 g_76_6 (.ZN (n_76_6), .A (n_75_5), .B (n_72_5), .C1 (n_68_7), .C2 (n_62_10) );
AOI211_X1 g_75_4 (.ZN (n_75_4), .A (n_77_4), .B (n_74_4), .C1 (n_70_6), .C2 (n_64_9) );
AOI211_X1 g_77_3 (.ZN (n_77_3), .A (n_76_6), .B (n_73_6), .C1 (n_72_5), .C2 (n_66_8) );
AOI211_X1 g_79_2 (.ZN (n_79_2), .A (n_75_4), .B (n_75_5), .C1 (n_74_4), .C2 (n_68_7) );
AOI211_X1 g_81_1 (.ZN (n_81_1), .A (n_77_3), .B (n_77_4), .C1 (n_73_6), .C2 (n_70_6) );
AOI211_X1 g_80_3 (.ZN (n_80_3), .A (n_79_2), .B (n_76_6), .C1 (n_75_5), .C2 (n_72_5) );
AOI211_X1 g_82_2 (.ZN (n_82_2), .A (n_81_1), .B (n_75_4), .C1 (n_77_4), .C2 (n_74_4) );
AOI211_X1 g_84_1 (.ZN (n_84_1), .A (n_80_3), .B (n_77_3), .C1 (n_76_6), .C2 (n_73_6) );
AOI211_X1 g_83_3 (.ZN (n_83_3), .A (n_82_2), .B (n_79_2), .C1 (n_75_4), .C2 (n_75_5) );
AOI211_X1 g_82_1 (.ZN (n_82_1), .A (n_84_1), .B (n_81_1), .C1 (n_77_3), .C2 (n_77_4) );
AOI211_X1 g_80_2 (.ZN (n_80_2), .A (n_83_3), .B (n_80_3), .C1 (n_79_2), .C2 (n_76_6) );
AOI211_X1 g_78_3 (.ZN (n_78_3), .A (n_82_1), .B (n_82_2), .C1 (n_81_1), .C2 (n_75_4) );
AOI211_X1 g_76_4 (.ZN (n_76_4), .A (n_80_2), .B (n_84_1), .C1 (n_80_3), .C2 (n_77_3) );
AOI211_X1 g_74_5 (.ZN (n_74_5), .A (n_78_3), .B (n_83_3), .C1 (n_82_2), .C2 (n_79_2) );
AOI211_X1 g_72_6 (.ZN (n_72_6), .A (n_76_4), .B (n_82_1), .C1 (n_84_1), .C2 (n_81_1) );
AOI211_X1 g_70_7 (.ZN (n_70_7), .A (n_74_5), .B (n_80_2), .C1 (n_83_3), .C2 (n_80_3) );
AOI211_X1 g_68_8 (.ZN (n_68_8), .A (n_72_6), .B (n_78_3), .C1 (n_82_1), .C2 (n_82_2) );
AOI211_X1 g_69_6 (.ZN (n_69_6), .A (n_70_7), .B (n_76_4), .C1 (n_80_2), .C2 (n_84_1) );
AOI211_X1 g_67_7 (.ZN (n_67_7), .A (n_68_8), .B (n_74_5), .C1 (n_78_3), .C2 (n_83_3) );
AOI211_X1 g_65_8 (.ZN (n_65_8), .A (n_69_6), .B (n_72_6), .C1 (n_76_4), .C2 (n_82_1) );
AOI211_X1 g_63_9 (.ZN (n_63_9), .A (n_67_7), .B (n_70_7), .C1 (n_74_5), .C2 (n_80_2) );
AOI211_X1 g_61_10 (.ZN (n_61_10), .A (n_65_8), .B (n_68_8), .C1 (n_72_6), .C2 (n_78_3) );
AOI211_X1 g_59_11 (.ZN (n_59_11), .A (n_63_9), .B (n_69_6), .C1 (n_70_7), .C2 (n_76_4) );
AOI211_X1 g_57_12 (.ZN (n_57_12), .A (n_61_10), .B (n_67_7), .C1 (n_68_8), .C2 (n_74_5) );
AOI211_X1 g_55_13 (.ZN (n_55_13), .A (n_59_11), .B (n_65_8), .C1 (n_69_6), .C2 (n_72_6) );
AOI211_X1 g_53_14 (.ZN (n_53_14), .A (n_57_12), .B (n_63_9), .C1 (n_67_7), .C2 (n_70_7) );
AOI211_X1 g_51_15 (.ZN (n_51_15), .A (n_55_13), .B (n_61_10), .C1 (n_65_8), .C2 (n_68_8) );
AOI211_X1 g_49_16 (.ZN (n_49_16), .A (n_53_14), .B (n_59_11), .C1 (n_63_9), .C2 (n_69_6) );
AOI211_X1 g_47_17 (.ZN (n_47_17), .A (n_51_15), .B (n_57_12), .C1 (n_61_10), .C2 (n_67_7) );
AOI211_X1 g_45_18 (.ZN (n_45_18), .A (n_49_16), .B (n_55_13), .C1 (n_59_11), .C2 (n_65_8) );
AOI211_X1 g_43_19 (.ZN (n_43_19), .A (n_47_17), .B (n_53_14), .C1 (n_57_12), .C2 (n_63_9) );
AOI211_X1 g_41_20 (.ZN (n_41_20), .A (n_45_18), .B (n_51_15), .C1 (n_55_13), .C2 (n_61_10) );
AOI211_X1 g_39_21 (.ZN (n_39_21), .A (n_43_19), .B (n_49_16), .C1 (n_53_14), .C2 (n_59_11) );
AOI211_X1 g_37_20 (.ZN (n_37_20), .A (n_41_20), .B (n_47_17), .C1 (n_51_15), .C2 (n_57_12) );
AOI211_X1 g_35_21 (.ZN (n_35_21), .A (n_39_21), .B (n_45_18), .C1 (n_49_16), .C2 (n_55_13) );
AOI211_X1 g_33_22 (.ZN (n_33_22), .A (n_37_20), .B (n_43_19), .C1 (n_47_17), .C2 (n_53_14) );
AOI211_X1 g_31_23 (.ZN (n_31_23), .A (n_35_21), .B (n_41_20), .C1 (n_45_18), .C2 (n_51_15) );
AOI211_X1 g_29_24 (.ZN (n_29_24), .A (n_33_22), .B (n_39_21), .C1 (n_43_19), .C2 (n_49_16) );
AOI211_X1 g_27_25 (.ZN (n_27_25), .A (n_31_23), .B (n_37_20), .C1 (n_41_20), .C2 (n_47_17) );
AOI211_X1 g_28_23 (.ZN (n_28_23), .A (n_29_24), .B (n_35_21), .C1 (n_39_21), .C2 (n_45_18) );
AOI211_X1 g_26_24 (.ZN (n_26_24), .A (n_27_25), .B (n_33_22), .C1 (n_37_20), .C2 (n_43_19) );
AOI211_X1 g_24_25 (.ZN (n_24_25), .A (n_28_23), .B (n_31_23), .C1 (n_35_21), .C2 (n_41_20) );
AOI211_X1 g_22_26 (.ZN (n_22_26), .A (n_26_24), .B (n_29_24), .C1 (n_33_22), .C2 (n_39_21) );
AOI211_X1 g_20_27 (.ZN (n_20_27), .A (n_24_25), .B (n_27_25), .C1 (n_31_23), .C2 (n_37_20) );
AOI211_X1 g_18_28 (.ZN (n_18_28), .A (n_22_26), .B (n_28_23), .C1 (n_29_24), .C2 (n_35_21) );
AOI211_X1 g_19_26 (.ZN (n_19_26), .A (n_20_27), .B (n_26_24), .C1 (n_27_25), .C2 (n_33_22) );
AOI211_X1 g_17_27 (.ZN (n_17_27), .A (n_18_28), .B (n_24_25), .C1 (n_28_23), .C2 (n_31_23) );
AOI211_X1 g_16_29 (.ZN (n_16_29), .A (n_19_26), .B (n_22_26), .C1 (n_26_24), .C2 (n_29_24) );
AOI211_X1 g_14_30 (.ZN (n_14_30), .A (n_17_27), .B (n_20_27), .C1 (n_24_25), .C2 (n_27_25) );
AOI211_X1 g_13_32 (.ZN (n_13_32), .A (n_16_29), .B (n_18_28), .C1 (n_22_26), .C2 (n_28_23) );
AOI211_X1 g_11_31 (.ZN (n_11_31), .A (n_14_30), .B (n_19_26), .C1 (n_20_27), .C2 (n_26_24) );
AOI211_X1 g_9_32 (.ZN (n_9_32), .A (n_13_32), .B (n_17_27), .C1 (n_18_28), .C2 (n_24_25) );
AOI211_X1 g_7_33 (.ZN (n_7_33), .A (n_11_31), .B (n_16_29), .C1 (n_19_26), .C2 (n_22_26) );
AOI211_X1 g_6_35 (.ZN (n_6_35), .A (n_9_32), .B (n_14_30), .C1 (n_17_27), .C2 (n_20_27) );
AOI211_X1 g_5_37 (.ZN (n_5_37), .A (n_7_33), .B (n_13_32), .C1 (n_16_29), .C2 (n_18_28) );
AOI211_X1 g_4_39 (.ZN (n_4_39), .A (n_6_35), .B (n_11_31), .C1 (n_14_30), .C2 (n_19_26) );
AOI211_X1 g_6_40 (.ZN (n_6_40), .A (n_5_37), .B (n_9_32), .C1 (n_13_32), .C2 (n_17_27) );
AOI211_X1 g_4_41 (.ZN (n_4_41), .A (n_4_39), .B (n_7_33), .C1 (n_11_31), .C2 (n_16_29) );
AOI211_X1 g_2_42 (.ZN (n_2_42), .A (n_6_40), .B (n_6_35), .C1 (n_9_32), .C2 (n_14_30) );
AOI211_X1 g_3_40 (.ZN (n_3_40), .A (n_4_41), .B (n_5_37), .C1 (n_7_33), .C2 (n_13_32) );
AOI211_X1 g_5_39 (.ZN (n_5_39), .A (n_2_42), .B (n_4_39), .C1 (n_6_35), .C2 (n_11_31) );
AOI211_X1 g_7_38 (.ZN (n_7_38), .A (n_3_40), .B (n_6_40), .C1 (n_5_37), .C2 (n_9_32) );
AOI211_X1 g_8_36 (.ZN (n_8_36), .A (n_5_39), .B (n_4_41), .C1 (n_4_39), .C2 (n_7_33) );
AOI211_X1 g_6_37 (.ZN (n_6_37), .A (n_7_38), .B (n_2_42), .C1 (n_6_40), .C2 (n_6_35) );
AOI211_X1 g_4_38 (.ZN (n_4_38), .A (n_8_36), .B (n_3_40), .C1 (n_4_41), .C2 (n_5_37) );
AOI211_X1 g_5_36 (.ZN (n_5_36), .A (n_6_37), .B (n_5_39), .C1 (n_2_42), .C2 (n_4_39) );
AOI211_X1 g_7_35 (.ZN (n_7_35), .A (n_4_38), .B (n_7_38), .C1 (n_3_40), .C2 (n_6_40) );
AOI211_X1 g_9_34 (.ZN (n_9_34), .A (n_5_36), .B (n_8_36), .C1 (n_5_39), .C2 (n_4_41) );
AOI211_X1 g_11_33 (.ZN (n_11_33), .A (n_7_35), .B (n_6_37), .C1 (n_7_38), .C2 (n_2_42) );
AOI211_X1 g_10_35 (.ZN (n_10_35), .A (n_9_34), .B (n_4_38), .C1 (n_8_36), .C2 (n_3_40) );
AOI211_X1 g_8_34 (.ZN (n_8_34), .A (n_11_33), .B (n_5_36), .C1 (n_6_37), .C2 (n_5_39) );
AOI211_X1 g_7_32 (.ZN (n_7_32), .A (n_10_35), .B (n_7_35), .C1 (n_4_38), .C2 (n_7_38) );
AOI211_X1 g_9_31 (.ZN (n_9_31), .A (n_8_34), .B (n_9_34), .C1 (n_5_36), .C2 (n_8_36) );
AOI211_X1 g_8_33 (.ZN (n_8_33), .A (n_7_32), .B (n_11_33), .C1 (n_7_35), .C2 (n_6_37) );
AOI211_X1 g_10_32 (.ZN (n_10_32), .A (n_9_31), .B (n_10_35), .C1 (n_9_34), .C2 (n_4_38) );
AOI211_X1 g_11_34 (.ZN (n_11_34), .A (n_8_33), .B (n_8_34), .C1 (n_11_33), .C2 (n_5_36) );
AOI211_X1 g_12_32 (.ZN (n_12_32), .A (n_10_32), .B (n_7_32), .C1 (n_10_35), .C2 (n_7_35) );
AOI211_X1 g_10_33 (.ZN (n_10_33), .A (n_11_34), .B (n_9_31), .C1 (n_8_34), .C2 (n_9_34) );
AOI211_X1 g_9_35 (.ZN (n_9_35), .A (n_12_32), .B (n_8_33), .C1 (n_7_32), .C2 (n_11_33) );
AOI211_X1 g_7_36 (.ZN (n_7_36), .A (n_10_33), .B (n_10_32), .C1 (n_9_31), .C2 (n_10_35) );
AOI211_X1 g_6_34 (.ZN (n_6_34), .A (n_9_35), .B (n_11_34), .C1 (n_8_33), .C2 (n_8_34) );
AOI211_X1 g_8_35 (.ZN (n_8_35), .A (n_7_36), .B (n_12_32), .C1 (n_10_32), .C2 (n_7_32) );
AOI211_X1 g_7_37 (.ZN (n_7_37), .A (n_6_34), .B (n_10_33), .C1 (n_11_34), .C2 (n_9_31) );
AOI211_X1 g_6_39 (.ZN (n_6_39), .A (n_8_35), .B (n_9_35), .C1 (n_12_32), .C2 (n_8_33) );
AOI211_X1 g_5_41 (.ZN (n_5_41), .A (n_7_37), .B (n_7_36), .C1 (n_10_33), .C2 (n_10_32) );
AOI211_X1 g_4_43 (.ZN (n_4_43), .A (n_6_39), .B (n_6_34), .C1 (n_9_35), .C2 (n_11_34) );
AOI211_X1 g_6_44 (.ZN (n_6_44), .A (n_5_41), .B (n_8_35), .C1 (n_7_36), .C2 (n_12_32) );
AOI211_X1 g_4_45 (.ZN (n_4_45), .A (n_4_43), .B (n_7_37), .C1 (n_6_34), .C2 (n_10_33) );
AOI211_X1 g_2_46 (.ZN (n_2_46), .A (n_6_44), .B (n_6_39), .C1 (n_8_35), .C2 (n_9_35) );
AOI211_X1 g_3_44 (.ZN (n_3_44), .A (n_4_45), .B (n_5_41), .C1 (n_7_37), .C2 (n_7_36) );
AOI211_X1 g_5_43 (.ZN (n_5_43), .A (n_2_46), .B (n_4_43), .C1 (n_6_39), .C2 (n_6_34) );
AOI211_X1 g_7_42 (.ZN (n_7_42), .A (n_3_44), .B (n_6_44), .C1 (n_5_41), .C2 (n_8_35) );
AOI211_X1 g_8_40 (.ZN (n_8_40), .A (n_5_43), .B (n_4_45), .C1 (n_4_43), .C2 (n_7_37) );
AOI211_X1 g_6_41 (.ZN (n_6_41), .A (n_7_42), .B (n_2_46), .C1 (n_6_44), .C2 (n_6_39) );
AOI211_X1 g_4_42 (.ZN (n_4_42), .A (n_8_40), .B (n_3_44), .C1 (n_4_45), .C2 (n_5_41) );
AOI211_X1 g_5_40 (.ZN (n_5_40), .A (n_6_41), .B (n_5_43), .C1 (n_2_46), .C2 (n_4_43) );
AOI211_X1 g_6_38 (.ZN (n_6_38), .A (n_4_42), .B (n_7_42), .C1 (n_3_44), .C2 (n_6_44) );
AOI211_X1 g_8_37 (.ZN (n_8_37), .A (n_5_40), .B (n_8_40), .C1 (n_5_43), .C2 (n_4_45) );
AOI211_X1 g_7_39 (.ZN (n_7_39), .A (n_6_38), .B (n_6_41), .C1 (n_7_42), .C2 (n_2_46) );
AOI211_X1 g_9_38 (.ZN (n_9_38), .A (n_8_37), .B (n_4_42), .C1 (n_8_40), .C2 (n_3_44) );
AOI211_X1 g_10_36 (.ZN (n_10_36), .A (n_7_39), .B (n_5_40), .C1 (n_6_41), .C2 (n_5_43) );
AOI211_X1 g_12_35 (.ZN (n_12_35), .A (n_9_38), .B (n_6_38), .C1 (n_4_42), .C2 (n_7_42) );
AOI211_X1 g_10_34 (.ZN (n_10_34), .A (n_10_36), .B (n_8_37), .C1 (n_5_40), .C2 (n_8_40) );
AOI211_X1 g_11_32 (.ZN (n_11_32), .A (n_12_35), .B (n_7_39), .C1 (n_6_38), .C2 (n_6_41) );
AOI211_X1 g_12_34 (.ZN (n_12_34), .A (n_10_34), .B (n_9_38), .C1 (n_8_37), .C2 (n_4_42) );
AOI211_X1 g_11_36 (.ZN (n_11_36), .A (n_11_32), .B (n_10_36), .C1 (n_7_39), .C2 (n_5_40) );
AOI211_X1 g_9_37 (.ZN (n_9_37), .A (n_12_34), .B (n_12_35), .C1 (n_9_38), .C2 (n_6_38) );
AOI211_X1 g_8_39 (.ZN (n_8_39), .A (n_11_36), .B (n_10_34), .C1 (n_10_36), .C2 (n_8_37) );
AOI211_X1 g_7_41 (.ZN (n_7_41), .A (n_9_37), .B (n_11_32), .C1 (n_12_35), .C2 (n_7_39) );
AOI211_X1 g_6_43 (.ZN (n_6_43), .A (n_8_39), .B (n_12_34), .C1 (n_10_34), .C2 (n_9_38) );
AOI211_X1 g_5_45 (.ZN (n_5_45), .A (n_7_41), .B (n_11_36), .C1 (n_11_32), .C2 (n_10_36) );
AOI211_X1 g_4_47 (.ZN (n_4_47), .A (n_6_43), .B (n_9_37), .C1 (n_12_34), .C2 (n_12_35) );
AOI211_X1 g_6_48 (.ZN (n_6_48), .A (n_5_45), .B (n_8_39), .C1 (n_11_36), .C2 (n_10_34) );
AOI211_X1 g_4_49 (.ZN (n_4_49), .A (n_4_47), .B (n_7_41), .C1 (n_9_37), .C2 (n_11_32) );
AOI211_X1 g_2_50 (.ZN (n_2_50), .A (n_6_48), .B (n_6_43), .C1 (n_8_39), .C2 (n_12_34) );
AOI211_X1 g_3_48 (.ZN (n_3_48), .A (n_4_49), .B (n_5_45), .C1 (n_7_41), .C2 (n_11_36) );
AOI211_X1 g_5_47 (.ZN (n_5_47), .A (n_2_50), .B (n_4_47), .C1 (n_6_43), .C2 (n_9_37) );
AOI211_X1 g_7_46 (.ZN (n_7_46), .A (n_3_48), .B (n_6_48), .C1 (n_5_45), .C2 (n_8_39) );
AOI211_X1 g_8_44 (.ZN (n_8_44), .A (n_5_47), .B (n_4_49), .C1 (n_4_47), .C2 (n_7_41) );
AOI211_X1 g_6_45 (.ZN (n_6_45), .A (n_7_46), .B (n_2_50), .C1 (n_6_48), .C2 (n_6_43) );
AOI211_X1 g_4_46 (.ZN (n_4_46), .A (n_8_44), .B (n_3_48), .C1 (n_4_49), .C2 (n_5_45) );
AOI211_X1 g_5_44 (.ZN (n_5_44), .A (n_6_45), .B (n_5_47), .C1 (n_2_50), .C2 (n_4_47) );
AOI211_X1 g_7_43 (.ZN (n_7_43), .A (n_4_46), .B (n_7_46), .C1 (n_3_48), .C2 (n_6_48) );
AOI211_X1 g_9_42 (.ZN (n_9_42), .A (n_5_44), .B (n_8_44), .C1 (n_5_47), .C2 (n_4_49) );
AOI211_X1 g_10_40 (.ZN (n_10_40), .A (n_7_43), .B (n_6_45), .C1 (n_7_46), .C2 (n_2_50) );
AOI211_X1 g_8_41 (.ZN (n_8_41), .A (n_9_42), .B (n_4_46), .C1 (n_8_44), .C2 (n_3_48) );
AOI211_X1 g_6_42 (.ZN (n_6_42), .A (n_10_40), .B (n_5_44), .C1 (n_6_45), .C2 (n_5_47) );
AOI211_X1 g_7_40 (.ZN (n_7_40), .A (n_8_41), .B (n_7_43), .C1 (n_4_46), .C2 (n_7_46) );
AOI211_X1 g_9_39 (.ZN (n_9_39), .A (n_6_42), .B (n_9_42), .C1 (n_5_44), .C2 (n_8_44) );
AOI211_X1 g_11_38 (.ZN (n_11_38), .A (n_7_40), .B (n_10_40), .C1 (n_7_43), .C2 (n_6_45) );
AOI211_X1 g_13_37 (.ZN (n_13_37), .A (n_9_39), .B (n_8_41), .C1 (n_9_42), .C2 (n_4_46) );
AOI211_X1 g_14_35 (.ZN (n_14_35), .A (n_11_38), .B (n_6_42), .C1 (n_10_40), .C2 (n_5_44) );
AOI211_X1 g_13_33 (.ZN (n_13_33), .A (n_13_37), .B (n_7_40), .C1 (n_8_41), .C2 (n_7_43) );
AOI211_X1 g_14_31 (.ZN (n_14_31), .A (n_14_35), .B (n_9_39), .C1 (n_6_42), .C2 (n_9_42) );
AOI211_X1 g_16_30 (.ZN (n_16_30), .A (n_13_33), .B (n_11_38), .C1 (n_7_40), .C2 (n_10_40) );
AOI211_X1 g_14_29 (.ZN (n_14_29), .A (n_14_31), .B (n_13_37), .C1 (n_9_39), .C2 (n_8_41) );
AOI211_X1 g_16_28 (.ZN (n_16_28), .A (n_16_30), .B (n_14_35), .C1 (n_11_38), .C2 (n_6_42) );
AOI211_X1 g_18_27 (.ZN (n_18_27), .A (n_14_29), .B (n_13_33), .C1 (n_13_37), .C2 (n_7_40) );
AOI211_X1 g_20_26 (.ZN (n_20_26), .A (n_16_28), .B (n_14_31), .C1 (n_14_35), .C2 (n_9_39) );
AOI211_X1 g_19_28 (.ZN (n_19_28), .A (n_18_27), .B (n_16_30), .C1 (n_13_33), .C2 (n_11_38) );
AOI211_X1 g_21_27 (.ZN (n_21_27), .A (n_20_26), .B (n_14_29), .C1 (n_14_31), .C2 (n_13_37) );
AOI211_X1 g_23_26 (.ZN (n_23_26), .A (n_19_28), .B (n_16_28), .C1 (n_16_30), .C2 (n_14_35) );
AOI211_X1 g_25_25 (.ZN (n_25_25), .A (n_21_27), .B (n_18_27), .C1 (n_14_29), .C2 (n_13_33) );
AOI211_X1 g_24_27 (.ZN (n_24_27), .A (n_23_26), .B (n_20_26), .C1 (n_16_28), .C2 (n_14_31) );
AOI211_X1 g_26_26 (.ZN (n_26_26), .A (n_25_25), .B (n_19_28), .C1 (n_18_27), .C2 (n_16_30) );
AOI211_X1 g_28_25 (.ZN (n_28_25), .A (n_24_27), .B (n_21_27), .C1 (n_20_26), .C2 (n_14_29) );
AOI211_X1 g_30_24 (.ZN (n_30_24), .A (n_26_26), .B (n_23_26), .C1 (n_19_28), .C2 (n_16_28) );
AOI211_X1 g_32_23 (.ZN (n_32_23), .A (n_28_25), .B (n_25_25), .C1 (n_21_27), .C2 (n_18_27) );
AOI211_X1 g_34_22 (.ZN (n_34_22), .A (n_30_24), .B (n_24_27), .C1 (n_23_26), .C2 (n_20_26) );
AOI211_X1 g_33_24 (.ZN (n_33_24), .A (n_32_23), .B (n_26_26), .C1 (n_25_25), .C2 (n_19_28) );
AOI211_X1 g_35_23 (.ZN (n_35_23), .A (n_34_22), .B (n_28_25), .C1 (n_24_27), .C2 (n_21_27) );
AOI211_X1 g_37_22 (.ZN (n_37_22), .A (n_33_24), .B (n_30_24), .C1 (n_26_26), .C2 (n_23_26) );
AOI211_X1 g_36_24 (.ZN (n_36_24), .A (n_35_23), .B (n_32_23), .C1 (n_28_25), .C2 (n_25_25) );
AOI211_X1 g_35_22 (.ZN (n_35_22), .A (n_37_22), .B (n_34_22), .C1 (n_30_24), .C2 (n_24_27) );
AOI211_X1 g_37_21 (.ZN (n_37_21), .A (n_36_24), .B (n_33_24), .C1 (n_32_23), .C2 (n_26_26) );
AOI211_X1 g_39_20 (.ZN (n_39_20), .A (n_35_22), .B (n_35_23), .C1 (n_34_22), .C2 (n_28_25) );
AOI211_X1 g_41_19 (.ZN (n_41_19), .A (n_37_21), .B (n_37_22), .C1 (n_33_24), .C2 (n_30_24) );
AOI211_X1 g_40_21 (.ZN (n_40_21), .A (n_39_20), .B (n_36_24), .C1 (n_35_23), .C2 (n_32_23) );
AOI211_X1 g_42_20 (.ZN (n_42_20), .A (n_41_19), .B (n_35_22), .C1 (n_37_22), .C2 (n_34_22) );
AOI211_X1 g_44_19 (.ZN (n_44_19), .A (n_40_21), .B (n_37_21), .C1 (n_36_24), .C2 (n_33_24) );
AOI211_X1 g_46_18 (.ZN (n_46_18), .A (n_42_20), .B (n_39_20), .C1 (n_35_22), .C2 (n_35_23) );
AOI211_X1 g_48_17 (.ZN (n_48_17), .A (n_44_19), .B (n_41_19), .C1 (n_37_21), .C2 (n_37_22) );
AOI211_X1 g_50_16 (.ZN (n_50_16), .A (n_46_18), .B (n_40_21), .C1 (n_39_20), .C2 (n_36_24) );
AOI211_X1 g_52_15 (.ZN (n_52_15), .A (n_48_17), .B (n_42_20), .C1 (n_41_19), .C2 (n_35_22) );
AOI211_X1 g_51_17 (.ZN (n_51_17), .A (n_50_16), .B (n_44_19), .C1 (n_40_21), .C2 (n_37_21) );
AOI211_X1 g_50_15 (.ZN (n_50_15), .A (n_52_15), .B (n_46_18), .C1 (n_42_20), .C2 (n_39_20) );
AOI211_X1 g_52_14 (.ZN (n_52_14), .A (n_51_17), .B (n_48_17), .C1 (n_44_19), .C2 (n_41_19) );
AOI211_X1 g_54_13 (.ZN (n_54_13), .A (n_50_15), .B (n_50_16), .C1 (n_46_18), .C2 (n_40_21) );
AOI211_X1 g_56_12 (.ZN (n_56_12), .A (n_52_14), .B (n_52_15), .C1 (n_48_17), .C2 (n_42_20) );
AOI211_X1 g_58_11 (.ZN (n_58_11), .A (n_54_13), .B (n_51_17), .C1 (n_50_16), .C2 (n_44_19) );
AOI211_X1 g_60_10 (.ZN (n_60_10), .A (n_56_12), .B (n_50_15), .C1 (n_52_15), .C2 (n_46_18) );
AOI211_X1 g_59_12 (.ZN (n_59_12), .A (n_58_11), .B (n_52_14), .C1 (n_51_17), .C2 (n_48_17) );
AOI211_X1 g_61_11 (.ZN (n_61_11), .A (n_60_10), .B (n_54_13), .C1 (n_50_15), .C2 (n_50_16) );
AOI211_X1 g_63_10 (.ZN (n_63_10), .A (n_59_12), .B (n_56_12), .C1 (n_52_14), .C2 (n_52_15) );
AOI211_X1 g_65_9 (.ZN (n_65_9), .A (n_61_11), .B (n_58_11), .C1 (n_54_13), .C2 (n_51_17) );
AOI211_X1 g_67_8 (.ZN (n_67_8), .A (n_63_10), .B (n_60_10), .C1 (n_56_12), .C2 (n_50_15) );
AOI211_X1 g_69_7 (.ZN (n_69_7), .A (n_65_9), .B (n_59_12), .C1 (n_58_11), .C2 (n_52_14) );
AOI211_X1 g_71_6 (.ZN (n_71_6), .A (n_67_8), .B (n_61_11), .C1 (n_60_10), .C2 (n_54_13) );
AOI211_X1 g_73_5 (.ZN (n_73_5), .A (n_69_7), .B (n_63_10), .C1 (n_59_12), .C2 (n_56_12) );
AOI211_X1 g_74_7 (.ZN (n_74_7), .A (n_71_6), .B (n_65_9), .C1 (n_61_11), .C2 (n_58_11) );
AOI211_X1 g_72_8 (.ZN (n_72_8), .A (n_73_5), .B (n_67_8), .C1 (n_63_10), .C2 (n_60_10) );
AOI211_X1 g_70_9 (.ZN (n_70_9), .A (n_74_7), .B (n_69_7), .C1 (n_65_9), .C2 (n_59_12) );
AOI211_X1 g_71_7 (.ZN (n_71_7), .A (n_72_8), .B (n_71_6), .C1 (n_67_8), .C2 (n_61_11) );
AOI211_X1 g_69_8 (.ZN (n_69_8), .A (n_70_9), .B (n_73_5), .C1 (n_69_7), .C2 (n_63_10) );
AOI211_X1 g_67_9 (.ZN (n_67_9), .A (n_71_7), .B (n_74_7), .C1 (n_71_6), .C2 (n_65_9) );
AOI211_X1 g_65_10 (.ZN (n_65_10), .A (n_69_8), .B (n_72_8), .C1 (n_73_5), .C2 (n_67_8) );
AOI211_X1 g_63_11 (.ZN (n_63_11), .A (n_67_9), .B (n_70_9), .C1 (n_74_7), .C2 (n_69_7) );
AOI211_X1 g_61_12 (.ZN (n_61_12), .A (n_65_10), .B (n_71_7), .C1 (n_72_8), .C2 (n_71_6) );
AOI211_X1 g_59_13 (.ZN (n_59_13), .A (n_63_11), .B (n_69_8), .C1 (n_70_9), .C2 (n_73_5) );
AOI211_X1 g_57_14 (.ZN (n_57_14), .A (n_61_12), .B (n_67_9), .C1 (n_71_7), .C2 (n_74_7) );
AOI211_X1 g_55_15 (.ZN (n_55_15), .A (n_59_13), .B (n_65_10), .C1 (n_69_8), .C2 (n_72_8) );
AOI211_X1 g_53_16 (.ZN (n_53_16), .A (n_57_14), .B (n_63_11), .C1 (n_67_9), .C2 (n_70_9) );
AOI211_X1 g_52_18 (.ZN (n_52_18), .A (n_55_15), .B (n_61_12), .C1 (n_65_10), .C2 (n_71_7) );
AOI211_X1 g_51_16 (.ZN (n_51_16), .A (n_53_16), .B (n_59_13), .C1 (n_63_11), .C2 (n_69_8) );
AOI211_X1 g_53_15 (.ZN (n_53_15), .A (n_52_18), .B (n_57_14), .C1 (n_61_12), .C2 (n_67_9) );
AOI211_X1 g_55_14 (.ZN (n_55_14), .A (n_51_16), .B (n_55_15), .C1 (n_59_13), .C2 (n_65_10) );
AOI211_X1 g_57_13 (.ZN (n_57_13), .A (n_53_15), .B (n_53_16), .C1 (n_57_14), .C2 (n_63_11) );
AOI211_X1 g_56_15 (.ZN (n_56_15), .A (n_55_14), .B (n_52_18), .C1 (n_55_15), .C2 (n_61_12) );
AOI211_X1 g_58_14 (.ZN (n_58_14), .A (n_57_13), .B (n_51_16), .C1 (n_53_16), .C2 (n_59_13) );
AOI211_X1 g_60_13 (.ZN (n_60_13), .A (n_56_15), .B (n_53_15), .C1 (n_52_18), .C2 (n_57_14) );
AOI211_X1 g_62_12 (.ZN (n_62_12), .A (n_58_14), .B (n_55_14), .C1 (n_51_16), .C2 (n_55_15) );
AOI211_X1 g_64_11 (.ZN (n_64_11), .A (n_60_13), .B (n_57_13), .C1 (n_53_15), .C2 (n_53_16) );
AOI211_X1 g_66_10 (.ZN (n_66_10), .A (n_62_12), .B (n_56_15), .C1 (n_55_14), .C2 (n_52_18) );
AOI211_X1 g_68_9 (.ZN (n_68_9), .A (n_64_11), .B (n_58_14), .C1 (n_57_13), .C2 (n_51_16) );
AOI211_X1 g_70_8 (.ZN (n_70_8), .A (n_66_10), .B (n_60_13), .C1 (n_56_15), .C2 (n_53_15) );
AOI211_X1 g_72_7 (.ZN (n_72_7), .A (n_68_9), .B (n_62_12), .C1 (n_58_14), .C2 (n_55_14) );
AOI211_X1 g_74_6 (.ZN (n_74_6), .A (n_70_8), .B (n_64_11), .C1 (n_60_13), .C2 (n_57_13) );
AOI211_X1 g_76_5 (.ZN (n_76_5), .A (n_72_7), .B (n_66_10), .C1 (n_62_12), .C2 (n_56_15) );
AOI211_X1 g_78_4 (.ZN (n_78_4), .A (n_74_6), .B (n_68_9), .C1 (n_64_11), .C2 (n_58_14) );
AOI211_X1 g_77_6 (.ZN (n_77_6), .A (n_76_5), .B (n_70_8), .C1 (n_66_10), .C2 (n_60_13) );
AOI211_X1 g_79_5 (.ZN (n_79_5), .A (n_78_4), .B (n_72_7), .C1 (n_68_9), .C2 (n_62_12) );
AOI211_X1 g_81_4 (.ZN (n_81_4), .A (n_77_6), .B (n_74_6), .C1 (n_70_8), .C2 (n_64_11) );
AOI211_X1 g_80_6 (.ZN (n_80_6), .A (n_79_5), .B (n_76_5), .C1 (n_72_7), .C2 (n_66_10) );
AOI211_X1 g_78_5 (.ZN (n_78_5), .A (n_81_4), .B (n_78_4), .C1 (n_74_6), .C2 (n_68_9) );
AOI211_X1 g_80_4 (.ZN (n_80_4), .A (n_80_6), .B (n_77_6), .C1 (n_76_5), .C2 (n_70_8) );
AOI211_X1 g_82_3 (.ZN (n_82_3), .A (n_78_5), .B (n_79_5), .C1 (n_78_4), .C2 (n_72_7) );
AOI211_X1 g_84_2 (.ZN (n_84_2), .A (n_80_4), .B (n_81_4), .C1 (n_77_6), .C2 (n_74_6) );
AOI211_X1 g_86_1 (.ZN (n_86_1), .A (n_82_3), .B (n_80_6), .C1 (n_79_5), .C2 (n_76_5) );
AOI211_X1 g_87_3 (.ZN (n_87_3), .A (n_84_2), .B (n_78_5), .C1 (n_81_4), .C2 (n_78_4) );
AOI211_X1 g_88_1 (.ZN (n_88_1), .A (n_86_1), .B (n_80_4), .C1 (n_80_6), .C2 (n_77_6) );
AOI211_X1 g_86_2 (.ZN (n_86_2), .A (n_87_3), .B (n_82_3), .C1 (n_78_5), .C2 (n_79_5) );
AOI211_X1 g_85_4 (.ZN (n_85_4), .A (n_88_1), .B (n_84_2), .C1 (n_80_4), .C2 (n_81_4) );
AOI211_X1 g_83_5 (.ZN (n_83_5), .A (n_86_2), .B (n_86_1), .C1 (n_82_3), .C2 (n_80_6) );
AOI211_X1 g_84_3 (.ZN (n_84_3), .A (n_85_4), .B (n_87_3), .C1 (n_84_2), .C2 (n_78_5) );
AOI211_X1 g_85_1 (.ZN (n_85_1), .A (n_83_5), .B (n_88_1), .C1 (n_86_1), .C2 (n_80_4) );
AOI211_X1 g_83_2 (.ZN (n_83_2), .A (n_84_3), .B (n_86_2), .C1 (n_87_3), .C2 (n_82_3) );
AOI211_X1 g_81_3 (.ZN (n_81_3), .A (n_85_1), .B (n_85_4), .C1 (n_88_1), .C2 (n_84_2) );
AOI211_X1 g_79_4 (.ZN (n_79_4), .A (n_83_2), .B (n_83_5), .C1 (n_86_2), .C2 (n_86_1) );
AOI211_X1 g_77_5 (.ZN (n_77_5), .A (n_81_3), .B (n_84_3), .C1 (n_85_4), .C2 (n_87_3) );
AOI211_X1 g_75_6 (.ZN (n_75_6), .A (n_79_4), .B (n_85_1), .C1 (n_83_5), .C2 (n_88_1) );
AOI211_X1 g_73_7 (.ZN (n_73_7), .A (n_77_5), .B (n_83_2), .C1 (n_84_3), .C2 (n_86_2) );
AOI211_X1 g_71_8 (.ZN (n_71_8), .A (n_75_6), .B (n_81_3), .C1 (n_85_1), .C2 (n_85_4) );
AOI211_X1 g_69_9 (.ZN (n_69_9), .A (n_73_7), .B (n_79_4), .C1 (n_83_2), .C2 (n_83_5) );
AOI211_X1 g_67_10 (.ZN (n_67_10), .A (n_71_8), .B (n_77_5), .C1 (n_81_3), .C2 (n_84_3) );
AOI211_X1 g_65_11 (.ZN (n_65_11), .A (n_69_9), .B (n_75_6), .C1 (n_79_4), .C2 (n_85_1) );
AOI211_X1 g_66_9 (.ZN (n_66_9), .A (n_67_10), .B (n_73_7), .C1 (n_77_5), .C2 (n_83_2) );
AOI211_X1 g_64_10 (.ZN (n_64_10), .A (n_65_11), .B (n_71_8), .C1 (n_75_6), .C2 (n_81_3) );
AOI211_X1 g_62_11 (.ZN (n_62_11), .A (n_66_9), .B (n_69_9), .C1 (n_73_7), .C2 (n_79_4) );
AOI211_X1 g_60_12 (.ZN (n_60_12), .A (n_64_10), .B (n_67_10), .C1 (n_71_8), .C2 (n_77_5) );
AOI211_X1 g_58_13 (.ZN (n_58_13), .A (n_62_11), .B (n_65_11), .C1 (n_69_9), .C2 (n_75_6) );
AOI211_X1 g_56_14 (.ZN (n_56_14), .A (n_60_12), .B (n_66_9), .C1 (n_67_10), .C2 (n_73_7) );
AOI211_X1 g_54_15 (.ZN (n_54_15), .A (n_58_13), .B (n_64_10), .C1 (n_65_11), .C2 (n_71_8) );
AOI211_X1 g_52_16 (.ZN (n_52_16), .A (n_56_14), .B (n_62_11), .C1 (n_66_9), .C2 (n_69_9) );
AOI211_X1 g_50_17 (.ZN (n_50_17), .A (n_54_15), .B (n_60_12), .C1 (n_64_10), .C2 (n_67_10) );
AOI211_X1 g_48_16 (.ZN (n_48_16), .A (n_52_16), .B (n_58_13), .C1 (n_62_11), .C2 (n_65_11) );
AOI211_X1 g_46_17 (.ZN (n_46_17), .A (n_50_17), .B (n_56_14), .C1 (n_60_12), .C2 (n_66_9) );
AOI211_X1 g_44_18 (.ZN (n_44_18), .A (n_48_16), .B (n_54_15), .C1 (n_58_13), .C2 (n_64_10) );
AOI211_X1 g_42_19 (.ZN (n_42_19), .A (n_46_17), .B (n_52_16), .C1 (n_56_14), .C2 (n_62_11) );
AOI211_X1 g_41_21 (.ZN (n_41_21), .A (n_44_18), .B (n_50_17), .C1 (n_54_15), .C2 (n_60_12) );
AOI211_X1 g_43_20 (.ZN (n_43_20), .A (n_42_19), .B (n_48_16), .C1 (n_52_16), .C2 (n_58_13) );
AOI211_X1 g_45_19 (.ZN (n_45_19), .A (n_41_21), .B (n_46_17), .C1 (n_50_17), .C2 (n_56_14) );
AOI211_X1 g_47_18 (.ZN (n_47_18), .A (n_43_20), .B (n_44_18), .C1 (n_48_16), .C2 (n_54_15) );
AOI211_X1 g_49_17 (.ZN (n_49_17), .A (n_45_19), .B (n_42_19), .C1 (n_46_17), .C2 (n_52_16) );
AOI211_X1 g_48_19 (.ZN (n_48_19), .A (n_47_18), .B (n_41_21), .C1 (n_44_18), .C2 (n_50_17) );
AOI211_X1 g_50_18 (.ZN (n_50_18), .A (n_49_17), .B (n_43_20), .C1 (n_42_19), .C2 (n_48_16) );
AOI211_X1 g_52_17 (.ZN (n_52_17), .A (n_48_19), .B (n_45_19), .C1 (n_41_21), .C2 (n_46_17) );
AOI211_X1 g_54_16 (.ZN (n_54_16), .A (n_50_18), .B (n_47_18), .C1 (n_43_20), .C2 (n_44_18) );
AOI211_X1 g_53_18 (.ZN (n_53_18), .A (n_52_17), .B (n_49_17), .C1 (n_45_19), .C2 (n_42_19) );
AOI211_X1 g_55_17 (.ZN (n_55_17), .A (n_54_16), .B (n_48_19), .C1 (n_47_18), .C2 (n_41_21) );
AOI211_X1 g_57_16 (.ZN (n_57_16), .A (n_53_18), .B (n_50_18), .C1 (n_49_17), .C2 (n_43_20) );
AOI211_X1 g_59_15 (.ZN (n_59_15), .A (n_55_17), .B (n_52_17), .C1 (n_48_19), .C2 (n_45_19) );
AOI211_X1 g_61_14 (.ZN (n_61_14), .A (n_57_16), .B (n_54_16), .C1 (n_50_18), .C2 (n_47_18) );
AOI211_X1 g_63_13 (.ZN (n_63_13), .A (n_59_15), .B (n_53_18), .C1 (n_52_17), .C2 (n_49_17) );
AOI211_X1 g_65_12 (.ZN (n_65_12), .A (n_61_14), .B (n_55_17), .C1 (n_54_16), .C2 (n_48_19) );
AOI211_X1 g_67_11 (.ZN (n_67_11), .A (n_63_13), .B (n_57_16), .C1 (n_53_18), .C2 (n_50_18) );
AOI211_X1 g_69_10 (.ZN (n_69_10), .A (n_65_12), .B (n_59_15), .C1 (n_55_17), .C2 (n_52_17) );
AOI211_X1 g_71_9 (.ZN (n_71_9), .A (n_67_11), .B (n_61_14), .C1 (n_57_16), .C2 (n_54_16) );
AOI211_X1 g_73_8 (.ZN (n_73_8), .A (n_69_10), .B (n_63_13), .C1 (n_59_15), .C2 (n_53_18) );
AOI211_X1 g_75_7 (.ZN (n_75_7), .A (n_71_9), .B (n_65_12), .C1 (n_61_14), .C2 (n_55_17) );
AOI211_X1 g_74_9 (.ZN (n_74_9), .A (n_73_8), .B (n_67_11), .C1 (n_63_13), .C2 (n_57_16) );
AOI211_X1 g_76_8 (.ZN (n_76_8), .A (n_75_7), .B (n_69_10), .C1 (n_65_12), .C2 (n_59_15) );
AOI211_X1 g_78_7 (.ZN (n_78_7), .A (n_74_9), .B (n_71_9), .C1 (n_67_11), .C2 (n_61_14) );
AOI211_X1 g_77_9 (.ZN (n_77_9), .A (n_76_8), .B (n_73_8), .C1 (n_69_10), .C2 (n_63_13) );
AOI211_X1 g_76_7 (.ZN (n_76_7), .A (n_78_7), .B (n_75_7), .C1 (n_71_9), .C2 (n_65_12) );
AOI211_X1 g_78_6 (.ZN (n_78_6), .A (n_77_9), .B (n_74_9), .C1 (n_73_8), .C2 (n_67_11) );
AOI211_X1 g_80_5 (.ZN (n_80_5), .A (n_76_7), .B (n_76_8), .C1 (n_75_7), .C2 (n_69_10) );
AOI211_X1 g_82_4 (.ZN (n_82_4), .A (n_78_6), .B (n_78_7), .C1 (n_74_9), .C2 (n_71_9) );
AOI211_X1 g_81_6 (.ZN (n_81_6), .A (n_80_5), .B (n_77_9), .C1 (n_76_8), .C2 (n_73_8) );
AOI211_X1 g_79_7 (.ZN (n_79_7), .A (n_82_4), .B (n_76_7), .C1 (n_78_7), .C2 (n_75_7) );
AOI211_X1 g_77_8 (.ZN (n_77_8), .A (n_81_6), .B (n_78_6), .C1 (n_77_9), .C2 (n_74_9) );
AOI211_X1 g_75_9 (.ZN (n_75_9), .A (n_79_7), .B (n_80_5), .C1 (n_76_7), .C2 (n_76_8) );
AOI211_X1 g_73_10 (.ZN (n_73_10), .A (n_77_8), .B (n_82_4), .C1 (n_78_6), .C2 (n_78_7) );
AOI211_X1 g_74_8 (.ZN (n_74_8), .A (n_75_9), .B (n_81_6), .C1 (n_80_5), .C2 (n_77_9) );
AOI211_X1 g_72_9 (.ZN (n_72_9), .A (n_73_10), .B (n_79_7), .C1 (n_82_4), .C2 (n_76_7) );
AOI211_X1 g_70_10 (.ZN (n_70_10), .A (n_74_8), .B (n_77_8), .C1 (n_81_6), .C2 (n_78_6) );
AOI211_X1 g_68_11 (.ZN (n_68_11), .A (n_72_9), .B (n_75_9), .C1 (n_79_7), .C2 (n_80_5) );
AOI211_X1 g_66_12 (.ZN (n_66_12), .A (n_70_10), .B (n_73_10), .C1 (n_77_8), .C2 (n_82_4) );
AOI211_X1 g_64_13 (.ZN (n_64_13), .A (n_68_11), .B (n_74_8), .C1 (n_75_9), .C2 (n_81_6) );
AOI211_X1 g_62_14 (.ZN (n_62_14), .A (n_66_12), .B (n_72_9), .C1 (n_73_10), .C2 (n_79_7) );
AOI211_X1 g_63_12 (.ZN (n_63_12), .A (n_64_13), .B (n_70_10), .C1 (n_74_8), .C2 (n_77_8) );
AOI211_X1 g_61_13 (.ZN (n_61_13), .A (n_62_14), .B (n_68_11), .C1 (n_72_9), .C2 (n_75_9) );
AOI211_X1 g_59_14 (.ZN (n_59_14), .A (n_63_12), .B (n_66_12), .C1 (n_70_10), .C2 (n_73_10) );
AOI211_X1 g_57_15 (.ZN (n_57_15), .A (n_61_13), .B (n_64_13), .C1 (n_68_11), .C2 (n_74_8) );
AOI211_X1 g_55_16 (.ZN (n_55_16), .A (n_59_14), .B (n_62_14), .C1 (n_66_12), .C2 (n_72_9) );
AOI211_X1 g_53_17 (.ZN (n_53_17), .A (n_57_15), .B (n_63_12), .C1 (n_64_13), .C2 (n_70_10) );
AOI211_X1 g_51_18 (.ZN (n_51_18), .A (n_55_16), .B (n_61_13), .C1 (n_62_14), .C2 (n_68_11) );
AOI211_X1 g_49_19 (.ZN (n_49_19), .A (n_53_17), .B (n_59_14), .C1 (n_63_12), .C2 (n_66_12) );
AOI211_X1 g_47_20 (.ZN (n_47_20), .A (n_51_18), .B (n_57_15), .C1 (n_61_13), .C2 (n_64_13) );
AOI211_X1 g_48_18 (.ZN (n_48_18), .A (n_49_19), .B (n_55_16), .C1 (n_59_14), .C2 (n_62_14) );
AOI211_X1 g_46_19 (.ZN (n_46_19), .A (n_47_20), .B (n_53_17), .C1 (n_57_15), .C2 (n_63_12) );
AOI211_X1 g_44_20 (.ZN (n_44_20), .A (n_48_18), .B (n_51_18), .C1 (n_55_16), .C2 (n_61_13) );
AOI211_X1 g_42_21 (.ZN (n_42_21), .A (n_46_19), .B (n_49_19), .C1 (n_53_17), .C2 (n_59_14) );
AOI211_X1 g_40_22 (.ZN (n_40_22), .A (n_44_20), .B (n_47_20), .C1 (n_51_18), .C2 (n_57_15) );
AOI211_X1 g_38_21 (.ZN (n_38_21), .A (n_42_21), .B (n_48_18), .C1 (n_49_19), .C2 (n_55_16) );
AOI211_X1 g_36_22 (.ZN (n_36_22), .A (n_40_22), .B (n_46_19), .C1 (n_47_20), .C2 (n_53_17) );
AOI211_X1 g_34_23 (.ZN (n_34_23), .A (n_38_21), .B (n_44_20), .C1 (n_48_18), .C2 (n_51_18) );
AOI211_X1 g_32_24 (.ZN (n_32_24), .A (n_36_22), .B (n_42_21), .C1 (n_46_19), .C2 (n_49_19) );
AOI211_X1 g_30_25 (.ZN (n_30_25), .A (n_34_23), .B (n_40_22), .C1 (n_44_20), .C2 (n_47_20) );
AOI211_X1 g_28_26 (.ZN (n_28_26), .A (n_32_24), .B (n_38_21), .C1 (n_42_21), .C2 (n_48_18) );
AOI211_X1 g_26_25 (.ZN (n_26_25), .A (n_30_25), .B (n_36_22), .C1 (n_40_22), .C2 (n_46_19) );
AOI211_X1 g_24_26 (.ZN (n_24_26), .A (n_28_26), .B (n_34_23), .C1 (n_38_21), .C2 (n_44_20) );
AOI211_X1 g_22_27 (.ZN (n_22_27), .A (n_26_25), .B (n_32_24), .C1 (n_36_22), .C2 (n_42_21) );
AOI211_X1 g_20_28 (.ZN (n_20_28), .A (n_24_26), .B (n_30_25), .C1 (n_34_23), .C2 (n_40_22) );
AOI211_X1 g_18_29 (.ZN (n_18_29), .A (n_22_27), .B (n_28_26), .C1 (n_32_24), .C2 (n_38_21) );
AOI211_X1 g_17_31 (.ZN (n_17_31), .A (n_20_28), .B (n_26_25), .C1 (n_30_25), .C2 (n_36_22) );
AOI211_X1 g_15_30 (.ZN (n_15_30), .A (n_18_29), .B (n_24_26), .C1 (n_28_26), .C2 (n_34_23) );
AOI211_X1 g_17_29 (.ZN (n_17_29), .A (n_17_31), .B (n_22_27), .C1 (n_26_25), .C2 (n_32_24) );
AOI211_X1 g_19_30 (.ZN (n_19_30), .A (n_15_30), .B (n_20_28), .C1 (n_24_26), .C2 (n_30_25) );
AOI211_X1 g_21_29 (.ZN (n_21_29), .A (n_17_29), .B (n_18_29), .C1 (n_22_27), .C2 (n_28_26) );
AOI211_X1 g_23_28 (.ZN (n_23_28), .A (n_19_30), .B (n_17_31), .C1 (n_20_28), .C2 (n_26_25) );
AOI211_X1 g_25_27 (.ZN (n_25_27), .A (n_21_29), .B (n_15_30), .C1 (n_18_29), .C2 (n_24_26) );
AOI211_X1 g_27_26 (.ZN (n_27_26), .A (n_23_28), .B (n_17_29), .C1 (n_17_31), .C2 (n_22_27) );
AOI211_X1 g_29_25 (.ZN (n_29_25), .A (n_25_27), .B (n_19_30), .C1 (n_15_30), .C2 (n_20_28) );
AOI211_X1 g_31_24 (.ZN (n_31_24), .A (n_27_26), .B (n_21_29), .C1 (n_17_29), .C2 (n_18_29) );
AOI211_X1 g_33_23 (.ZN (n_33_23), .A (n_29_25), .B (n_23_28), .C1 (n_19_30), .C2 (n_17_31) );
AOI211_X1 g_34_25 (.ZN (n_34_25), .A (n_31_24), .B (n_25_27), .C1 (n_21_29), .C2 (n_15_30) );
AOI211_X1 g_32_26 (.ZN (n_32_26), .A (n_33_23), .B (n_27_26), .C1 (n_23_28), .C2 (n_17_29) );
AOI211_X1 g_30_27 (.ZN (n_30_27), .A (n_34_25), .B (n_29_25), .C1 (n_25_27), .C2 (n_19_30) );
AOI211_X1 g_31_25 (.ZN (n_31_25), .A (n_32_26), .B (n_31_24), .C1 (n_27_26), .C2 (n_21_29) );
AOI211_X1 g_29_26 (.ZN (n_29_26), .A (n_30_27), .B (n_33_23), .C1 (n_29_25), .C2 (n_23_28) );
AOI211_X1 g_27_27 (.ZN (n_27_27), .A (n_31_25), .B (n_34_25), .C1 (n_31_24), .C2 (n_25_27) );
AOI211_X1 g_25_26 (.ZN (n_25_26), .A (n_29_26), .B (n_32_26), .C1 (n_33_23), .C2 (n_27_26) );
AOI211_X1 g_23_27 (.ZN (n_23_27), .A (n_27_27), .B (n_30_27), .C1 (n_34_25), .C2 (n_29_25) );
AOI211_X1 g_21_28 (.ZN (n_21_28), .A (n_25_26), .B (n_31_25), .C1 (n_32_26), .C2 (n_31_24) );
AOI211_X1 g_19_29 (.ZN (n_19_29), .A (n_23_27), .B (n_29_26), .C1 (n_30_27), .C2 (n_33_23) );
AOI211_X1 g_17_30 (.ZN (n_17_30), .A (n_21_28), .B (n_27_27), .C1 (n_31_25), .C2 (n_34_25) );
AOI211_X1 g_15_31 (.ZN (n_15_31), .A (n_19_29), .B (n_25_26), .C1 (n_29_26), .C2 (n_32_26) );
AOI211_X1 g_14_33 (.ZN (n_14_33), .A (n_17_30), .B (n_23_27), .C1 (n_27_27), .C2 (n_30_27) );
AOI211_X1 g_13_31 (.ZN (n_13_31), .A (n_15_31), .B (n_21_28), .C1 (n_25_26), .C2 (n_31_25) );
AOI211_X1 g_15_32 (.ZN (n_15_32), .A (n_14_33), .B (n_19_29), .C1 (n_23_27), .C2 (n_29_26) );
AOI211_X1 g_14_34 (.ZN (n_14_34), .A (n_13_31), .B (n_17_30), .C1 (n_21_28), .C2 (n_27_27) );
AOI211_X1 g_12_33 (.ZN (n_12_33), .A (n_15_32), .B (n_15_31), .C1 (n_19_29), .C2 (n_25_26) );
AOI211_X1 g_14_32 (.ZN (n_14_32), .A (n_14_34), .B (n_14_33), .C1 (n_17_30), .C2 (n_23_27) );
AOI211_X1 g_16_31 (.ZN (n_16_31), .A (n_12_33), .B (n_13_31), .C1 (n_15_31), .C2 (n_21_28) );
AOI211_X1 g_18_30 (.ZN (n_18_30), .A (n_14_32), .B (n_15_32), .C1 (n_14_33), .C2 (n_19_29) );
AOI211_X1 g_20_29 (.ZN (n_20_29), .A (n_16_31), .B (n_14_34), .C1 (n_13_31), .C2 (n_17_30) );
AOI211_X1 g_22_28 (.ZN (n_22_28), .A (n_18_30), .B (n_12_33), .C1 (n_15_32), .C2 (n_15_31) );
AOI211_X1 g_21_30 (.ZN (n_21_30), .A (n_20_29), .B (n_14_32), .C1 (n_14_34), .C2 (n_14_33) );
AOI211_X1 g_23_29 (.ZN (n_23_29), .A (n_22_28), .B (n_16_31), .C1 (n_12_33), .C2 (n_13_31) );
AOI211_X1 g_25_28 (.ZN (n_25_28), .A (n_21_30), .B (n_18_30), .C1 (n_14_32), .C2 (n_15_32) );
AOI211_X1 g_24_30 (.ZN (n_24_30), .A (n_23_29), .B (n_20_29), .C1 (n_16_31), .C2 (n_14_34) );
AOI211_X1 g_22_29 (.ZN (n_22_29), .A (n_25_28), .B (n_22_28), .C1 (n_18_30), .C2 (n_12_33) );
AOI211_X1 g_24_28 (.ZN (n_24_28), .A (n_24_30), .B (n_21_30), .C1 (n_20_29), .C2 (n_14_32) );
AOI211_X1 g_26_27 (.ZN (n_26_27), .A (n_22_29), .B (n_23_29), .C1 (n_22_28), .C2 (n_16_31) );
AOI211_X1 g_28_28 (.ZN (n_28_28), .A (n_24_28), .B (n_25_28), .C1 (n_21_30), .C2 (n_18_30) );
AOI211_X1 g_26_29 (.ZN (n_26_29), .A (n_26_27), .B (n_24_30), .C1 (n_23_29), .C2 (n_20_29) );
AOI211_X1 g_25_31 (.ZN (n_25_31), .A (n_28_28), .B (n_22_29), .C1 (n_25_28), .C2 (n_22_28) );
AOI211_X1 g_24_29 (.ZN (n_24_29), .A (n_26_29), .B (n_24_28), .C1 (n_24_30), .C2 (n_21_30) );
AOI211_X1 g_26_28 (.ZN (n_26_28), .A (n_25_31), .B (n_26_27), .C1 (n_22_29), .C2 (n_23_29) );
AOI211_X1 g_28_27 (.ZN (n_28_27), .A (n_24_29), .B (n_28_28), .C1 (n_24_28), .C2 (n_25_28) );
AOI211_X1 g_30_26 (.ZN (n_30_26), .A (n_26_28), .B (n_26_29), .C1 (n_26_27), .C2 (n_24_30) );
AOI211_X1 g_32_25 (.ZN (n_32_25), .A (n_28_27), .B (n_25_31), .C1 (n_28_28), .C2 (n_22_29) );
AOI211_X1 g_34_24 (.ZN (n_34_24), .A (n_30_26), .B (n_24_29), .C1 (n_26_29), .C2 (n_24_28) );
AOI211_X1 g_36_23 (.ZN (n_36_23), .A (n_32_25), .B (n_26_28), .C1 (n_25_31), .C2 (n_26_27) );
AOI211_X1 g_38_22 (.ZN (n_38_22), .A (n_34_24), .B (n_28_27), .C1 (n_24_29), .C2 (n_28_28) );
AOI211_X1 g_37_24 (.ZN (n_37_24), .A (n_36_23), .B (n_30_26), .C1 (n_26_28), .C2 (n_26_29) );
AOI211_X1 g_39_23 (.ZN (n_39_23), .A (n_38_22), .B (n_32_25), .C1 (n_28_27), .C2 (n_25_31) );
AOI211_X1 g_41_22 (.ZN (n_41_22), .A (n_37_24), .B (n_34_24), .C1 (n_30_26), .C2 (n_24_29) );
AOI211_X1 g_43_21 (.ZN (n_43_21), .A (n_39_23), .B (n_36_23), .C1 (n_32_25), .C2 (n_26_28) );
AOI211_X1 g_45_20 (.ZN (n_45_20), .A (n_41_22), .B (n_38_22), .C1 (n_34_24), .C2 (n_28_27) );
AOI211_X1 g_47_19 (.ZN (n_47_19), .A (n_43_21), .B (n_37_24), .C1 (n_36_23), .C2 (n_30_26) );
AOI211_X1 g_49_18 (.ZN (n_49_18), .A (n_45_20), .B (n_39_23), .C1 (n_38_22), .C2 (n_32_25) );
AOI211_X1 g_51_19 (.ZN (n_51_19), .A (n_47_19), .B (n_41_22), .C1 (n_37_24), .C2 (n_34_24) );
AOI211_X1 g_49_20 (.ZN (n_49_20), .A (n_49_18), .B (n_43_21), .C1 (n_39_23), .C2 (n_36_23) );
AOI211_X1 g_47_21 (.ZN (n_47_21), .A (n_51_19), .B (n_45_20), .C1 (n_41_22), .C2 (n_38_22) );
AOI211_X1 g_45_22 (.ZN (n_45_22), .A (n_49_20), .B (n_47_19), .C1 (n_43_21), .C2 (n_37_24) );
AOI211_X1 g_46_20 (.ZN (n_46_20), .A (n_47_21), .B (n_49_18), .C1 (n_45_20), .C2 (n_39_23) );
AOI211_X1 g_44_21 (.ZN (n_44_21), .A (n_45_22), .B (n_51_19), .C1 (n_47_19), .C2 (n_41_22) );
AOI211_X1 g_42_22 (.ZN (n_42_22), .A (n_46_20), .B (n_49_20), .C1 (n_49_18), .C2 (n_43_21) );
AOI211_X1 g_40_23 (.ZN (n_40_23), .A (n_44_21), .B (n_47_21), .C1 (n_51_19), .C2 (n_45_20) );
AOI211_X1 g_38_24 (.ZN (n_38_24), .A (n_42_22), .B (n_45_22), .C1 (n_49_20), .C2 (n_47_19) );
AOI211_X1 g_39_22 (.ZN (n_39_22), .A (n_40_23), .B (n_46_20), .C1 (n_47_21), .C2 (n_49_18) );
AOI211_X1 g_37_23 (.ZN (n_37_23), .A (n_38_24), .B (n_44_21), .C1 (n_45_22), .C2 (n_51_19) );
AOI211_X1 g_35_24 (.ZN (n_35_24), .A (n_39_22), .B (n_42_22), .C1 (n_46_20), .C2 (n_49_20) );
AOI211_X1 g_33_25 (.ZN (n_33_25), .A (n_37_23), .B (n_40_23), .C1 (n_44_21), .C2 (n_47_21) );
AOI211_X1 g_31_26 (.ZN (n_31_26), .A (n_35_24), .B (n_38_24), .C1 (n_42_22), .C2 (n_45_22) );
AOI211_X1 g_29_27 (.ZN (n_29_27), .A (n_33_25), .B (n_39_22), .C1 (n_40_23), .C2 (n_46_20) );
AOI211_X1 g_27_28 (.ZN (n_27_28), .A (n_31_26), .B (n_37_23), .C1 (n_38_24), .C2 (n_44_21) );
AOI211_X1 g_25_29 (.ZN (n_25_29), .A (n_29_27), .B (n_35_24), .C1 (n_39_22), .C2 (n_42_22) );
AOI211_X1 g_23_30 (.ZN (n_23_30), .A (n_27_28), .B (n_33_25), .C1 (n_37_23), .C2 (n_40_23) );
AOI211_X1 g_21_31 (.ZN (n_21_31), .A (n_25_29), .B (n_31_26), .C1 (n_35_24), .C2 (n_38_24) );
AOI211_X1 g_19_32 (.ZN (n_19_32), .A (n_23_30), .B (n_29_27), .C1 (n_33_25), .C2 (n_39_22) );
AOI211_X1 g_20_30 (.ZN (n_20_30), .A (n_21_31), .B (n_27_28), .C1 (n_31_26), .C2 (n_37_23) );
AOI211_X1 g_18_31 (.ZN (n_18_31), .A (n_19_32), .B (n_25_29), .C1 (n_29_27), .C2 (n_35_24) );
AOI211_X1 g_16_32 (.ZN (n_16_32), .A (n_20_30), .B (n_23_30), .C1 (n_27_28), .C2 (n_33_25) );
AOI211_X1 g_15_34 (.ZN (n_15_34), .A (n_18_31), .B (n_21_31), .C1 (n_25_29), .C2 (n_31_26) );
AOI211_X1 g_17_33 (.ZN (n_17_33), .A (n_16_32), .B (n_19_32), .C1 (n_23_30), .C2 (n_29_27) );
AOI211_X1 g_16_35 (.ZN (n_16_35), .A (n_15_34), .B (n_20_30), .C1 (n_21_31), .C2 (n_27_28) );
AOI211_X1 g_15_33 (.ZN (n_15_33), .A (n_17_33), .B (n_18_31), .C1 (n_19_32), .C2 (n_25_29) );
AOI211_X1 g_17_32 (.ZN (n_17_32), .A (n_16_35), .B (n_16_32), .C1 (n_20_30), .C2 (n_23_30) );
AOI211_X1 g_19_31 (.ZN (n_19_31), .A (n_15_33), .B (n_15_34), .C1 (n_18_31), .C2 (n_21_31) );
AOI211_X1 g_18_33 (.ZN (n_18_33), .A (n_17_32), .B (n_17_33), .C1 (n_16_32), .C2 (n_19_32) );
AOI211_X1 g_16_34 (.ZN (n_16_34), .A (n_19_31), .B (n_16_35), .C1 (n_15_34), .C2 (n_20_30) );
AOI211_X1 g_15_36 (.ZN (n_15_36), .A (n_18_33), .B (n_15_33), .C1 (n_17_33), .C2 (n_18_31) );
AOI211_X1 g_13_35 (.ZN (n_13_35), .A (n_16_34), .B (n_17_32), .C1 (n_16_35), .C2 (n_16_32) );
AOI211_X1 g_12_37 (.ZN (n_12_37), .A (n_15_36), .B (n_19_31), .C1 (n_15_33), .C2 (n_15_34) );
AOI211_X1 g_14_36 (.ZN (n_14_36), .A (n_13_35), .B (n_18_33), .C1 (n_17_32), .C2 (n_17_33) );
AOI211_X1 g_13_34 (.ZN (n_13_34), .A (n_12_37), .B (n_16_34), .C1 (n_19_31), .C2 (n_16_35) );
AOI211_X1 g_11_35 (.ZN (n_11_35), .A (n_14_36), .B (n_15_36), .C1 (n_18_33), .C2 (n_15_33) );
AOI211_X1 g_9_36 (.ZN (n_9_36), .A (n_13_34), .B (n_13_35), .C1 (n_16_34), .C2 (n_17_32) );
AOI211_X1 g_8_38 (.ZN (n_8_38), .A (n_11_35), .B (n_12_37), .C1 (n_15_36), .C2 (n_19_31) );
AOI211_X1 g_10_37 (.ZN (n_10_37), .A (n_9_36), .B (n_14_36), .C1 (n_13_35), .C2 (n_18_33) );
AOI211_X1 g_12_36 (.ZN (n_12_36), .A (n_8_38), .B (n_13_34), .C1 (n_12_37), .C2 (n_16_34) );
AOI211_X1 g_13_38 (.ZN (n_13_38), .A (n_10_37), .B (n_11_35), .C1 (n_14_36), .C2 (n_15_36) );
AOI211_X1 g_11_37 (.ZN (n_11_37), .A (n_12_36), .B (n_9_36), .C1 (n_13_34), .C2 (n_13_35) );
AOI211_X1 g_13_36 (.ZN (n_13_36), .A (n_13_38), .B (n_8_38), .C1 (n_11_35), .C2 (n_12_37) );
AOI211_X1 g_15_37 (.ZN (n_15_37), .A (n_11_37), .B (n_10_37), .C1 (n_9_36), .C2 (n_14_36) );
AOI211_X1 g_17_36 (.ZN (n_17_36), .A (n_13_36), .B (n_12_36), .C1 (n_8_38), .C2 (n_13_34) );
AOI211_X1 g_18_34 (.ZN (n_18_34), .A (n_15_37), .B (n_13_38), .C1 (n_10_37), .C2 (n_11_35) );
AOI211_X1 g_16_33 (.ZN (n_16_33), .A (n_17_36), .B (n_11_37), .C1 (n_12_36), .C2 (n_9_36) );
AOI211_X1 g_15_35 (.ZN (n_15_35), .A (n_18_34), .B (n_13_36), .C1 (n_13_38), .C2 (n_8_38) );
AOI211_X1 g_17_34 (.ZN (n_17_34), .A (n_16_33), .B (n_15_37), .C1 (n_11_37), .C2 (n_10_37) );
AOI211_X1 g_18_32 (.ZN (n_18_32), .A (n_15_35), .B (n_17_36), .C1 (n_13_36), .C2 (n_12_36) );
AOI211_X1 g_20_31 (.ZN (n_20_31), .A (n_17_34), .B (n_18_34), .C1 (n_15_37), .C2 (n_13_38) );
AOI211_X1 g_22_30 (.ZN (n_22_30), .A (n_18_32), .B (n_16_33), .C1 (n_17_36), .C2 (n_11_37) );
AOI211_X1 g_23_32 (.ZN (n_23_32), .A (n_20_31), .B (n_15_35), .C1 (n_18_34), .C2 (n_13_36) );
AOI211_X1 g_21_33 (.ZN (n_21_33), .A (n_22_30), .B (n_17_34), .C1 (n_16_33), .C2 (n_15_37) );
AOI211_X1 g_22_31 (.ZN (n_22_31), .A (n_23_32), .B (n_18_32), .C1 (n_15_35), .C2 (n_17_36) );
AOI211_X1 g_20_32 (.ZN (n_20_32), .A (n_21_33), .B (n_20_31), .C1 (n_17_34), .C2 (n_18_34) );
AOI211_X1 g_19_34 (.ZN (n_19_34), .A (n_22_31), .B (n_22_30), .C1 (n_18_32), .C2 (n_16_33) );
AOI211_X1 g_17_35 (.ZN (n_17_35), .A (n_20_32), .B (n_23_32), .C1 (n_20_31), .C2 (n_15_35) );
AOI211_X1 g_16_37 (.ZN (n_16_37), .A (n_19_34), .B (n_21_33), .C1 (n_22_30), .C2 (n_17_34) );
AOI211_X1 g_18_36 (.ZN (n_18_36), .A (n_17_35), .B (n_22_31), .C1 (n_23_32), .C2 (n_18_32) );
AOI211_X1 g_20_35 (.ZN (n_20_35), .A (n_16_37), .B (n_20_32), .C1 (n_21_33), .C2 (n_20_31) );
AOI211_X1 g_19_33 (.ZN (n_19_33), .A (n_18_36), .B (n_19_34), .C1 (n_22_31), .C2 (n_22_30) );
AOI211_X1 g_21_32 (.ZN (n_21_32), .A (n_20_35), .B (n_17_35), .C1 (n_20_32), .C2 (n_23_32) );
AOI211_X1 g_23_31 (.ZN (n_23_31), .A (n_19_33), .B (n_16_37), .C1 (n_19_34), .C2 (n_21_33) );
AOI211_X1 g_25_30 (.ZN (n_25_30), .A (n_21_32), .B (n_18_36), .C1 (n_17_35), .C2 (n_22_31) );
AOI211_X1 g_27_29 (.ZN (n_27_29), .A (n_23_31), .B (n_20_35), .C1 (n_16_37), .C2 (n_20_32) );
AOI211_X1 g_29_28 (.ZN (n_29_28), .A (n_25_30), .B (n_19_33), .C1 (n_18_36), .C2 (n_19_34) );
AOI211_X1 g_31_27 (.ZN (n_31_27), .A (n_27_29), .B (n_21_32), .C1 (n_20_35), .C2 (n_17_35) );
AOI211_X1 g_33_26 (.ZN (n_33_26), .A (n_29_28), .B (n_23_31), .C1 (n_19_33), .C2 (n_16_37) );
AOI211_X1 g_35_25 (.ZN (n_35_25), .A (n_31_27), .B (n_25_30), .C1 (n_21_32), .C2 (n_18_36) );
AOI211_X1 g_34_27 (.ZN (n_34_27), .A (n_33_26), .B (n_27_29), .C1 (n_23_31), .C2 (n_20_35) );
AOI211_X1 g_36_26 (.ZN (n_36_26), .A (n_35_25), .B (n_29_28), .C1 (n_25_30), .C2 (n_19_33) );
AOI211_X1 g_38_25 (.ZN (n_38_25), .A (n_34_27), .B (n_31_27), .C1 (n_27_29), .C2 (n_21_32) );
AOI211_X1 g_40_24 (.ZN (n_40_24), .A (n_36_26), .B (n_33_26), .C1 (n_29_28), .C2 (n_23_31) );
AOI211_X1 g_38_23 (.ZN (n_38_23), .A (n_38_25), .B (n_35_25), .C1 (n_31_27), .C2 (n_25_30) );
AOI211_X1 g_37_25 (.ZN (n_37_25), .A (n_40_24), .B (n_34_27), .C1 (n_33_26), .C2 (n_27_29) );
AOI211_X1 g_39_24 (.ZN (n_39_24), .A (n_38_23), .B (n_36_26), .C1 (n_35_25), .C2 (n_29_28) );
AOI211_X1 g_41_23 (.ZN (n_41_23), .A (n_37_25), .B (n_38_25), .C1 (n_34_27), .C2 (n_31_27) );
AOI211_X1 g_43_22 (.ZN (n_43_22), .A (n_39_24), .B (n_40_24), .C1 (n_36_26), .C2 (n_33_26) );
AOI211_X1 g_45_21 (.ZN (n_45_21), .A (n_41_23), .B (n_38_23), .C1 (n_38_25), .C2 (n_35_25) );
AOI211_X1 g_44_23 (.ZN (n_44_23), .A (n_43_22), .B (n_37_25), .C1 (n_40_24), .C2 (n_34_27) );
AOI211_X1 g_46_22 (.ZN (n_46_22), .A (n_45_21), .B (n_39_24), .C1 (n_38_23), .C2 (n_36_26) );
AOI211_X1 g_48_21 (.ZN (n_48_21), .A (n_44_23), .B (n_41_23), .C1 (n_37_25), .C2 (n_38_25) );
AOI211_X1 g_50_20 (.ZN (n_50_20), .A (n_46_22), .B (n_43_22), .C1 (n_39_24), .C2 (n_40_24) );
AOI211_X1 g_52_19 (.ZN (n_52_19), .A (n_48_21), .B (n_45_21), .C1 (n_41_23), .C2 (n_38_23) );
AOI211_X1 g_54_18 (.ZN (n_54_18), .A (n_50_20), .B (n_44_23), .C1 (n_43_22), .C2 (n_37_25) );
AOI211_X1 g_56_17 (.ZN (n_56_17), .A (n_52_19), .B (n_46_22), .C1 (n_45_21), .C2 (n_39_24) );
AOI211_X1 g_58_16 (.ZN (n_58_16), .A (n_54_18), .B (n_48_21), .C1 (n_44_23), .C2 (n_41_23) );
AOI211_X1 g_60_15 (.ZN (n_60_15), .A (n_56_17), .B (n_50_20), .C1 (n_46_22), .C2 (n_43_22) );
AOI211_X1 g_59_17 (.ZN (n_59_17), .A (n_58_16), .B (n_52_19), .C1 (n_48_21), .C2 (n_45_21) );
AOI211_X1 g_58_15 (.ZN (n_58_15), .A (n_60_15), .B (n_54_18), .C1 (n_50_20), .C2 (n_44_23) );
AOI211_X1 g_60_14 (.ZN (n_60_14), .A (n_59_17), .B (n_56_17), .C1 (n_52_19), .C2 (n_46_22) );
AOI211_X1 g_62_13 (.ZN (n_62_13), .A (n_58_15), .B (n_58_16), .C1 (n_54_18), .C2 (n_48_21) );
AOI211_X1 g_64_12 (.ZN (n_64_12), .A (n_60_14), .B (n_60_15), .C1 (n_56_17), .C2 (n_50_20) );
AOI211_X1 g_66_11 (.ZN (n_66_11), .A (n_62_13), .B (n_59_17), .C1 (n_58_16), .C2 (n_52_19) );
AOI211_X1 g_68_10 (.ZN (n_68_10), .A (n_64_12), .B (n_58_15), .C1 (n_60_15), .C2 (n_54_18) );
AOI211_X1 g_67_12 (.ZN (n_67_12), .A (n_66_11), .B (n_60_14), .C1 (n_59_17), .C2 (n_56_17) );
AOI211_X1 g_69_11 (.ZN (n_69_11), .A (n_68_10), .B (n_62_13), .C1 (n_58_15), .C2 (n_58_16) );
AOI211_X1 g_71_10 (.ZN (n_71_10), .A (n_67_12), .B (n_64_12), .C1 (n_60_14), .C2 (n_60_15) );
AOI211_X1 g_73_9 (.ZN (n_73_9), .A (n_69_11), .B (n_66_11), .C1 (n_62_13), .C2 (n_59_17) );
AOI211_X1 g_75_8 (.ZN (n_75_8), .A (n_71_10), .B (n_68_10), .C1 (n_64_12), .C2 (n_58_15) );
AOI211_X1 g_77_7 (.ZN (n_77_7), .A (n_73_9), .B (n_67_12), .C1 (n_66_11), .C2 (n_60_14) );
AOI211_X1 g_79_6 (.ZN (n_79_6), .A (n_75_8), .B (n_69_11), .C1 (n_68_10), .C2 (n_62_13) );
AOI211_X1 g_81_5 (.ZN (n_81_5), .A (n_77_7), .B (n_71_10), .C1 (n_67_12), .C2 (n_64_12) );
AOI211_X1 g_83_4 (.ZN (n_83_4), .A (n_79_6), .B (n_73_9), .C1 (n_69_11), .C2 (n_66_11) );
AOI211_X1 g_85_3 (.ZN (n_85_3), .A (n_81_5), .B (n_75_8), .C1 (n_71_10), .C2 (n_68_10) );
AOI211_X1 g_87_2 (.ZN (n_87_2), .A (n_83_4), .B (n_77_7), .C1 (n_73_9), .C2 (n_67_12) );
AOI211_X1 g_89_1 (.ZN (n_89_1), .A (n_85_3), .B (n_79_6), .C1 (n_75_8), .C2 (n_69_11) );
AOI211_X1 g_88_3 (.ZN (n_88_3), .A (n_87_2), .B (n_81_5), .C1 (n_77_7), .C2 (n_71_10) );
AOI211_X1 g_90_2 (.ZN (n_90_2), .A (n_89_1), .B (n_83_4), .C1 (n_79_6), .C2 (n_73_9) );
AOI211_X1 g_92_1 (.ZN (n_92_1), .A (n_88_3), .B (n_85_3), .C1 (n_81_5), .C2 (n_75_8) );
AOI211_X1 g_91_3 (.ZN (n_91_3), .A (n_90_2), .B (n_87_2), .C1 (n_83_4), .C2 (n_77_7) );
AOI211_X1 g_90_1 (.ZN (n_90_1), .A (n_92_1), .B (n_89_1), .C1 (n_85_3), .C2 (n_79_6) );
AOI211_X1 g_88_2 (.ZN (n_88_2), .A (n_91_3), .B (n_88_3), .C1 (n_87_2), .C2 (n_81_5) );
AOI211_X1 g_86_3 (.ZN (n_86_3), .A (n_90_1), .B (n_90_2), .C1 (n_89_1), .C2 (n_83_4) );
AOI211_X1 g_84_4 (.ZN (n_84_4), .A (n_88_2), .B (n_92_1), .C1 (n_88_3), .C2 (n_85_3) );
AOI211_X1 g_82_5 (.ZN (n_82_5), .A (n_86_3), .B (n_91_3), .C1 (n_90_2), .C2 (n_87_2) );
AOI211_X1 g_81_7 (.ZN (n_81_7), .A (n_84_4), .B (n_90_1), .C1 (n_92_1), .C2 (n_89_1) );
AOI211_X1 g_79_8 (.ZN (n_79_8), .A (n_82_5), .B (n_88_2), .C1 (n_91_3), .C2 (n_88_3) );
AOI211_X1 g_78_10 (.ZN (n_78_10), .A (n_81_7), .B (n_86_3), .C1 (n_90_1), .C2 (n_90_2) );
AOI211_X1 g_76_9 (.ZN (n_76_9), .A (n_79_8), .B (n_84_4), .C1 (n_88_2), .C2 (n_92_1) );
AOI211_X1 g_78_8 (.ZN (n_78_8), .A (n_78_10), .B (n_82_5), .C1 (n_86_3), .C2 (n_91_3) );
AOI211_X1 g_80_7 (.ZN (n_80_7), .A (n_76_9), .B (n_81_7), .C1 (n_84_4), .C2 (n_90_1) );
AOI211_X1 g_82_6 (.ZN (n_82_6), .A (n_78_8), .B (n_79_8), .C1 (n_82_5), .C2 (n_88_2) );
AOI211_X1 g_84_5 (.ZN (n_84_5), .A (n_80_7), .B (n_78_10), .C1 (n_81_7), .C2 (n_86_3) );
AOI211_X1 g_86_4 (.ZN (n_86_4), .A (n_82_6), .B (n_76_9), .C1 (n_79_8), .C2 (n_84_4) );
AOI211_X1 g_85_6 (.ZN (n_85_6), .A (n_84_5), .B (n_78_8), .C1 (n_78_10), .C2 (n_82_5) );
AOI211_X1 g_87_5 (.ZN (n_87_5), .A (n_86_4), .B (n_80_7), .C1 (n_76_9), .C2 (n_81_7) );
AOI211_X1 g_89_4 (.ZN (n_89_4), .A (n_85_6), .B (n_82_6), .C1 (n_78_8), .C2 (n_79_8) );
AOI211_X1 g_88_6 (.ZN (n_88_6), .A (n_87_5), .B (n_84_5), .C1 (n_80_7), .C2 (n_78_10) );
AOI211_X1 g_87_4 (.ZN (n_87_4), .A (n_89_4), .B (n_86_4), .C1 (n_82_6), .C2 (n_76_9) );
AOI211_X1 g_89_3 (.ZN (n_89_3), .A (n_88_6), .B (n_85_6), .C1 (n_84_5), .C2 (n_78_8) );
AOI211_X1 g_91_2 (.ZN (n_91_2), .A (n_87_4), .B (n_87_5), .C1 (n_86_4), .C2 (n_80_7) );
AOI211_X1 g_93_1 (.ZN (n_93_1), .A (n_89_3), .B (n_89_4), .C1 (n_85_6), .C2 (n_82_6) );
AOI211_X1 g_92_3 (.ZN (n_92_3), .A (n_91_2), .B (n_88_6), .C1 (n_87_5), .C2 (n_84_5) );
AOI211_X1 g_94_2 (.ZN (n_94_2), .A (n_93_1), .B (n_87_4), .C1 (n_89_4), .C2 (n_86_4) );
AOI211_X1 g_96_1 (.ZN (n_96_1), .A (n_92_3), .B (n_89_3), .C1 (n_88_6), .C2 (n_85_6) );
AOI211_X1 g_95_3 (.ZN (n_95_3), .A (n_94_2), .B (n_91_2), .C1 (n_87_4), .C2 (n_87_5) );
AOI211_X1 g_94_1 (.ZN (n_94_1), .A (n_96_1), .B (n_93_1), .C1 (n_89_3), .C2 (n_89_4) );
AOI211_X1 g_92_2 (.ZN (n_92_2), .A (n_95_3), .B (n_92_3), .C1 (n_91_2), .C2 (n_88_6) );
AOI211_X1 g_90_3 (.ZN (n_90_3), .A (n_94_1), .B (n_94_2), .C1 (n_93_1), .C2 (n_87_4) );
AOI211_X1 g_88_4 (.ZN (n_88_4), .A (n_92_2), .B (n_96_1), .C1 (n_92_3), .C2 (n_89_3) );
AOI211_X1 g_86_5 (.ZN (n_86_5), .A (n_90_3), .B (n_95_3), .C1 (n_94_2), .C2 (n_91_2) );
AOI211_X1 g_84_6 (.ZN (n_84_6), .A (n_88_4), .B (n_94_1), .C1 (n_96_1), .C2 (n_93_1) );
AOI211_X1 g_82_7 (.ZN (n_82_7), .A (n_86_5), .B (n_92_2), .C1 (n_95_3), .C2 (n_92_3) );
AOI211_X1 g_80_8 (.ZN (n_80_8), .A (n_84_6), .B (n_90_3), .C1 (n_94_1), .C2 (n_94_2) );
AOI211_X1 g_78_9 (.ZN (n_78_9), .A (n_82_7), .B (n_88_4), .C1 (n_92_2), .C2 (n_96_1) );
AOI211_X1 g_76_10 (.ZN (n_76_10), .A (n_80_8), .B (n_86_5), .C1 (n_90_3), .C2 (n_95_3) );
AOI211_X1 g_74_11 (.ZN (n_74_11), .A (n_78_9), .B (n_84_6), .C1 (n_88_4), .C2 (n_94_1) );
AOI211_X1 g_72_10 (.ZN (n_72_10), .A (n_76_10), .B (n_82_7), .C1 (n_86_5), .C2 (n_92_2) );
AOI211_X1 g_70_11 (.ZN (n_70_11), .A (n_74_11), .B (n_80_8), .C1 (n_84_6), .C2 (n_90_3) );
AOI211_X1 g_68_12 (.ZN (n_68_12), .A (n_72_10), .B (n_78_9), .C1 (n_82_7), .C2 (n_88_4) );
AOI211_X1 g_66_13 (.ZN (n_66_13), .A (n_70_11), .B (n_76_10), .C1 (n_80_8), .C2 (n_86_5) );
AOI211_X1 g_64_14 (.ZN (n_64_14), .A (n_68_12), .B (n_74_11), .C1 (n_78_9), .C2 (n_84_6) );
AOI211_X1 g_62_15 (.ZN (n_62_15), .A (n_66_13), .B (n_72_10), .C1 (n_76_10), .C2 (n_82_7) );
AOI211_X1 g_60_16 (.ZN (n_60_16), .A (n_64_14), .B (n_70_11), .C1 (n_74_11), .C2 (n_80_8) );
AOI211_X1 g_58_17 (.ZN (n_58_17), .A (n_62_15), .B (n_68_12), .C1 (n_72_10), .C2 (n_78_9) );
AOI211_X1 g_56_16 (.ZN (n_56_16), .A (n_60_16), .B (n_66_13), .C1 (n_70_11), .C2 (n_76_10) );
AOI211_X1 g_54_17 (.ZN (n_54_17), .A (n_58_17), .B (n_64_14), .C1 (n_68_12), .C2 (n_74_11) );
AOI211_X1 g_56_18 (.ZN (n_56_18), .A (n_56_16), .B (n_62_15), .C1 (n_66_13), .C2 (n_72_10) );
AOI211_X1 g_54_19 (.ZN (n_54_19), .A (n_54_17), .B (n_60_16), .C1 (n_64_14), .C2 (n_70_11) );
AOI211_X1 g_52_20 (.ZN (n_52_20), .A (n_56_18), .B (n_58_17), .C1 (n_62_15), .C2 (n_68_12) );
AOI211_X1 g_50_19 (.ZN (n_50_19), .A (n_54_19), .B (n_56_16), .C1 (n_60_16), .C2 (n_66_13) );
AOI211_X1 g_48_20 (.ZN (n_48_20), .A (n_52_20), .B (n_54_17), .C1 (n_58_17), .C2 (n_64_14) );
AOI211_X1 g_46_21 (.ZN (n_46_21), .A (n_50_19), .B (n_56_18), .C1 (n_56_16), .C2 (n_62_15) );
AOI211_X1 g_44_22 (.ZN (n_44_22), .A (n_48_20), .B (n_54_19), .C1 (n_54_17), .C2 (n_60_16) );
AOI211_X1 g_42_23 (.ZN (n_42_23), .A (n_46_21), .B (n_52_20), .C1 (n_56_18), .C2 (n_58_17) );
AOI211_X1 g_41_25 (.ZN (n_41_25), .A (n_44_22), .B (n_50_19), .C1 (n_54_19), .C2 (n_56_16) );
AOI211_X1 g_43_24 (.ZN (n_43_24), .A (n_42_23), .B (n_48_20), .C1 (n_52_20), .C2 (n_54_17) );
AOI211_X1 g_45_23 (.ZN (n_45_23), .A (n_41_25), .B (n_46_21), .C1 (n_50_19), .C2 (n_56_18) );
AOI211_X1 g_47_22 (.ZN (n_47_22), .A (n_43_24), .B (n_44_22), .C1 (n_48_20), .C2 (n_54_19) );
AOI211_X1 g_49_21 (.ZN (n_49_21), .A (n_45_23), .B (n_42_23), .C1 (n_46_21), .C2 (n_52_20) );
AOI211_X1 g_51_20 (.ZN (n_51_20), .A (n_47_22), .B (n_41_25), .C1 (n_44_22), .C2 (n_50_19) );
AOI211_X1 g_53_19 (.ZN (n_53_19), .A (n_49_21), .B (n_43_24), .C1 (n_42_23), .C2 (n_48_20) );
AOI211_X1 g_55_18 (.ZN (n_55_18), .A (n_51_20), .B (n_45_23), .C1 (n_41_25), .C2 (n_46_21) );
AOI211_X1 g_57_17 (.ZN (n_57_17), .A (n_53_19), .B (n_47_22), .C1 (n_43_24), .C2 (n_44_22) );
AOI211_X1 g_59_16 (.ZN (n_59_16), .A (n_55_18), .B (n_49_21), .C1 (n_45_23), .C2 (n_42_23) );
AOI211_X1 g_61_15 (.ZN (n_61_15), .A (n_57_17), .B (n_51_20), .C1 (n_47_22), .C2 (n_41_25) );
AOI211_X1 g_63_14 (.ZN (n_63_14), .A (n_59_16), .B (n_53_19), .C1 (n_49_21), .C2 (n_43_24) );
AOI211_X1 g_65_13 (.ZN (n_65_13), .A (n_61_15), .B (n_55_18), .C1 (n_51_20), .C2 (n_45_23) );
AOI211_X1 g_64_15 (.ZN (n_64_15), .A (n_63_14), .B (n_57_17), .C1 (n_53_19), .C2 (n_47_22) );
AOI211_X1 g_66_14 (.ZN (n_66_14), .A (n_65_13), .B (n_59_16), .C1 (n_55_18), .C2 (n_49_21) );
AOI211_X1 g_68_13 (.ZN (n_68_13), .A (n_64_15), .B (n_61_15), .C1 (n_57_17), .C2 (n_51_20) );
AOI211_X1 g_70_12 (.ZN (n_70_12), .A (n_66_14), .B (n_63_14), .C1 (n_59_16), .C2 (n_53_19) );
AOI211_X1 g_72_11 (.ZN (n_72_11), .A (n_68_13), .B (n_65_13), .C1 (n_61_15), .C2 (n_55_18) );
AOI211_X1 g_74_10 (.ZN (n_74_10), .A (n_70_12), .B (n_64_15), .C1 (n_63_14), .C2 (n_57_17) );
AOI211_X1 g_76_11 (.ZN (n_76_11), .A (n_72_11), .B (n_66_14), .C1 (n_65_13), .C2 (n_59_16) );
AOI211_X1 g_74_12 (.ZN (n_74_12), .A (n_74_10), .B (n_68_13), .C1 (n_64_15), .C2 (n_61_15) );
AOI211_X1 g_75_10 (.ZN (n_75_10), .A (n_76_11), .B (n_70_12), .C1 (n_66_14), .C2 (n_63_14) );
AOI211_X1 g_73_11 (.ZN (n_73_11), .A (n_74_12), .B (n_72_11), .C1 (n_68_13), .C2 (n_65_13) );
AOI211_X1 g_71_12 (.ZN (n_71_12), .A (n_75_10), .B (n_74_10), .C1 (n_70_12), .C2 (n_64_15) );
AOI211_X1 g_69_13 (.ZN (n_69_13), .A (n_73_11), .B (n_76_11), .C1 (n_72_11), .C2 (n_66_14) );
AOI211_X1 g_67_14 (.ZN (n_67_14), .A (n_71_12), .B (n_74_12), .C1 (n_74_10), .C2 (n_68_13) );
AOI211_X1 g_65_15 (.ZN (n_65_15), .A (n_69_13), .B (n_75_10), .C1 (n_76_11), .C2 (n_70_12) );
AOI211_X1 g_63_16 (.ZN (n_63_16), .A (n_67_14), .B (n_73_11), .C1 (n_74_12), .C2 (n_72_11) );
AOI211_X1 g_61_17 (.ZN (n_61_17), .A (n_65_15), .B (n_71_12), .C1 (n_75_10), .C2 (n_74_10) );
AOI211_X1 g_59_18 (.ZN (n_59_18), .A (n_63_16), .B (n_69_13), .C1 (n_73_11), .C2 (n_76_11) );
AOI211_X1 g_57_19 (.ZN (n_57_19), .A (n_61_17), .B (n_67_14), .C1 (n_71_12), .C2 (n_74_12) );
AOI211_X1 g_55_20 (.ZN (n_55_20), .A (n_59_18), .B (n_65_15), .C1 (n_69_13), .C2 (n_75_10) );
AOI211_X1 g_53_21 (.ZN (n_53_21), .A (n_57_19), .B (n_63_16), .C1 (n_67_14), .C2 (n_73_11) );
AOI211_X1 g_51_22 (.ZN (n_51_22), .A (n_55_20), .B (n_61_17), .C1 (n_65_15), .C2 (n_71_12) );
AOI211_X1 g_49_23 (.ZN (n_49_23), .A (n_53_21), .B (n_59_18), .C1 (n_63_16), .C2 (n_69_13) );
AOI211_X1 g_50_21 (.ZN (n_50_21), .A (n_51_22), .B (n_57_19), .C1 (n_61_17), .C2 (n_67_14) );
AOI211_X1 g_48_22 (.ZN (n_48_22), .A (n_49_23), .B (n_55_20), .C1 (n_59_18), .C2 (n_65_15) );
AOI211_X1 g_46_23 (.ZN (n_46_23), .A (n_50_21), .B (n_53_21), .C1 (n_57_19), .C2 (n_63_16) );
AOI211_X1 g_44_24 (.ZN (n_44_24), .A (n_48_22), .B (n_51_22), .C1 (n_55_20), .C2 (n_61_17) );
AOI211_X1 g_42_25 (.ZN (n_42_25), .A (n_46_23), .B (n_49_23), .C1 (n_53_21), .C2 (n_59_18) );
AOI211_X1 g_43_23 (.ZN (n_43_23), .A (n_44_24), .B (n_50_21), .C1 (n_51_22), .C2 (n_57_19) );
AOI211_X1 g_41_24 (.ZN (n_41_24), .A (n_42_25), .B (n_48_22), .C1 (n_49_23), .C2 (n_55_20) );
AOI211_X1 g_39_25 (.ZN (n_39_25), .A (n_43_23), .B (n_46_23), .C1 (n_50_21), .C2 (n_53_21) );
AOI211_X1 g_37_26 (.ZN (n_37_26), .A (n_41_24), .B (n_44_24), .C1 (n_48_22), .C2 (n_51_22) );
AOI211_X1 g_35_27 (.ZN (n_35_27), .A (n_39_25), .B (n_42_25), .C1 (n_46_23), .C2 (n_49_23) );
AOI211_X1 g_36_25 (.ZN (n_36_25), .A (n_37_26), .B (n_43_23), .C1 (n_44_24), .C2 (n_50_21) );
AOI211_X1 g_34_26 (.ZN (n_34_26), .A (n_35_27), .B (n_41_24), .C1 (n_42_25), .C2 (n_48_22) );
AOI211_X1 g_32_27 (.ZN (n_32_27), .A (n_36_25), .B (n_39_25), .C1 (n_43_23), .C2 (n_46_23) );
AOI211_X1 g_30_28 (.ZN (n_30_28), .A (n_34_26), .B (n_37_26), .C1 (n_41_24), .C2 (n_44_24) );
AOI211_X1 g_28_29 (.ZN (n_28_29), .A (n_32_27), .B (n_35_27), .C1 (n_39_25), .C2 (n_42_25) );
AOI211_X1 g_26_30 (.ZN (n_26_30), .A (n_30_28), .B (n_36_25), .C1 (n_37_26), .C2 (n_43_23) );
AOI211_X1 g_24_31 (.ZN (n_24_31), .A (n_28_29), .B (n_34_26), .C1 (n_35_27), .C2 (n_41_24) );
AOI211_X1 g_22_32 (.ZN (n_22_32), .A (n_26_30), .B (n_32_27), .C1 (n_36_25), .C2 (n_39_25) );
AOI211_X1 g_20_33 (.ZN (n_20_33), .A (n_24_31), .B (n_30_28), .C1 (n_34_26), .C2 (n_37_26) );
AOI211_X1 g_19_35 (.ZN (n_19_35), .A (n_22_32), .B (n_28_29), .C1 (n_32_27), .C2 (n_35_27) );
AOI211_X1 g_21_34 (.ZN (n_21_34), .A (n_20_33), .B (n_26_30), .C1 (n_30_28), .C2 (n_36_25) );
AOI211_X1 g_23_33 (.ZN (n_23_33), .A (n_19_35), .B (n_24_31), .C1 (n_28_29), .C2 (n_34_26) );
AOI211_X1 g_25_32 (.ZN (n_25_32), .A (n_21_34), .B (n_22_32), .C1 (n_26_30), .C2 (n_32_27) );
AOI211_X1 g_27_31 (.ZN (n_27_31), .A (n_23_33), .B (n_20_33), .C1 (n_24_31), .C2 (n_30_28) );
AOI211_X1 g_29_30 (.ZN (n_29_30), .A (n_25_32), .B (n_19_35), .C1 (n_22_32), .C2 (n_28_29) );
AOI211_X1 g_31_29 (.ZN (n_31_29), .A (n_27_31), .B (n_21_34), .C1 (n_20_33), .C2 (n_26_30) );
AOI211_X1 g_33_28 (.ZN (n_33_28), .A (n_29_30), .B (n_23_33), .C1 (n_19_35), .C2 (n_24_31) );
AOI211_X1 g_35_29 (.ZN (n_35_29), .A (n_31_29), .B (n_25_32), .C1 (n_21_34), .C2 (n_22_32) );
AOI211_X1 g_36_27 (.ZN (n_36_27), .A (n_33_28), .B (n_27_31), .C1 (n_23_33), .C2 (n_20_33) );
AOI211_X1 g_38_26 (.ZN (n_38_26), .A (n_35_29), .B (n_29_30), .C1 (n_25_32), .C2 (n_19_35) );
AOI211_X1 g_40_25 (.ZN (n_40_25), .A (n_36_27), .B (n_31_29), .C1 (n_27_31), .C2 (n_21_34) );
AOI211_X1 g_42_24 (.ZN (n_42_24), .A (n_38_26), .B (n_33_28), .C1 (n_29_30), .C2 (n_23_33) );
AOI211_X1 g_41_26 (.ZN (n_41_26), .A (n_40_25), .B (n_35_29), .C1 (n_31_29), .C2 (n_25_32) );
AOI211_X1 g_43_25 (.ZN (n_43_25), .A (n_42_24), .B (n_36_27), .C1 (n_33_28), .C2 (n_27_31) );
AOI211_X1 g_45_24 (.ZN (n_45_24), .A (n_41_26), .B (n_38_26), .C1 (n_35_29), .C2 (n_29_30) );
AOI211_X1 g_47_23 (.ZN (n_47_23), .A (n_43_25), .B (n_40_25), .C1 (n_36_27), .C2 (n_31_29) );
AOI211_X1 g_49_22 (.ZN (n_49_22), .A (n_45_24), .B (n_42_24), .C1 (n_38_26), .C2 (n_33_28) );
AOI211_X1 g_51_21 (.ZN (n_51_21), .A (n_47_23), .B (n_41_26), .C1 (n_40_25), .C2 (n_35_29) );
AOI211_X1 g_53_20 (.ZN (n_53_20), .A (n_49_22), .B (n_43_25), .C1 (n_42_24), .C2 (n_36_27) );
AOI211_X1 g_55_19 (.ZN (n_55_19), .A (n_51_21), .B (n_45_24), .C1 (n_41_26), .C2 (n_38_26) );
AOI211_X1 g_57_18 (.ZN (n_57_18), .A (n_53_20), .B (n_47_23), .C1 (n_43_25), .C2 (n_40_25) );
AOI211_X1 g_56_20 (.ZN (n_56_20), .A (n_55_19), .B (n_49_22), .C1 (n_45_24), .C2 (n_42_24) );
AOI211_X1 g_58_19 (.ZN (n_58_19), .A (n_57_18), .B (n_51_21), .C1 (n_47_23), .C2 (n_41_26) );
AOI211_X1 g_60_18 (.ZN (n_60_18), .A (n_56_20), .B (n_53_20), .C1 (n_49_22), .C2 (n_43_25) );
AOI211_X1 g_61_16 (.ZN (n_61_16), .A (n_58_19), .B (n_55_19), .C1 (n_51_21), .C2 (n_45_24) );
AOI211_X1 g_63_15 (.ZN (n_63_15), .A (n_60_18), .B (n_57_18), .C1 (n_53_20), .C2 (n_47_23) );
AOI211_X1 g_65_14 (.ZN (n_65_14), .A (n_61_16), .B (n_56_20), .C1 (n_55_19), .C2 (n_49_22) );
AOI211_X1 g_67_13 (.ZN (n_67_13), .A (n_63_15), .B (n_58_19), .C1 (n_57_18), .C2 (n_51_21) );
AOI211_X1 g_69_12 (.ZN (n_69_12), .A (n_65_14), .B (n_60_18), .C1 (n_56_20), .C2 (n_53_20) );
AOI211_X1 g_71_11 (.ZN (n_71_11), .A (n_67_13), .B (n_61_16), .C1 (n_58_19), .C2 (n_55_19) );
AOI211_X1 g_72_13 (.ZN (n_72_13), .A (n_69_12), .B (n_63_15), .C1 (n_60_18), .C2 (n_57_18) );
AOI211_X1 g_70_14 (.ZN (n_70_14), .A (n_71_11), .B (n_65_14), .C1 (n_61_16), .C2 (n_56_20) );
AOI211_X1 g_68_15 (.ZN (n_68_15), .A (n_72_13), .B (n_67_13), .C1 (n_63_15), .C2 (n_58_19) );
AOI211_X1 g_66_16 (.ZN (n_66_16), .A (n_70_14), .B (n_69_12), .C1 (n_65_14), .C2 (n_60_18) );
AOI211_X1 g_64_17 (.ZN (n_64_17), .A (n_68_15), .B (n_71_11), .C1 (n_67_13), .C2 (n_61_16) );
AOI211_X1 g_62_16 (.ZN (n_62_16), .A (n_66_16), .B (n_72_13), .C1 (n_69_12), .C2 (n_63_15) );
AOI211_X1 g_60_17 (.ZN (n_60_17), .A (n_64_17), .B (n_70_14), .C1 (n_71_11), .C2 (n_65_14) );
AOI211_X1 g_58_18 (.ZN (n_58_18), .A (n_62_16), .B (n_68_15), .C1 (n_72_13), .C2 (n_67_13) );
AOI211_X1 g_56_19 (.ZN (n_56_19), .A (n_60_17), .B (n_66_16), .C1 (n_70_14), .C2 (n_69_12) );
AOI211_X1 g_54_20 (.ZN (n_54_20), .A (n_58_18), .B (n_64_17), .C1 (n_68_15), .C2 (n_71_11) );
AOI211_X1 g_52_21 (.ZN (n_52_21), .A (n_56_19), .B (n_62_16), .C1 (n_66_16), .C2 (n_72_13) );
AOI211_X1 g_50_22 (.ZN (n_50_22), .A (n_54_20), .B (n_60_17), .C1 (n_64_17), .C2 (n_70_14) );
AOI211_X1 g_48_23 (.ZN (n_48_23), .A (n_52_21), .B (n_58_18), .C1 (n_62_16), .C2 (n_68_15) );
AOI211_X1 g_46_24 (.ZN (n_46_24), .A (n_50_22), .B (n_56_19), .C1 (n_60_17), .C2 (n_66_16) );
AOI211_X1 g_44_25 (.ZN (n_44_25), .A (n_48_23), .B (n_54_20), .C1 (n_58_18), .C2 (n_64_17) );
AOI211_X1 g_42_26 (.ZN (n_42_26), .A (n_46_24), .B (n_52_21), .C1 (n_56_19), .C2 (n_62_16) );
AOI211_X1 g_40_27 (.ZN (n_40_27), .A (n_44_25), .B (n_50_22), .C1 (n_54_20), .C2 (n_60_17) );
AOI211_X1 g_38_28 (.ZN (n_38_28), .A (n_42_26), .B (n_48_23), .C1 (n_52_21), .C2 (n_58_18) );
AOI211_X1 g_39_26 (.ZN (n_39_26), .A (n_40_27), .B (n_46_24), .C1 (n_50_22), .C2 (n_56_19) );
AOI211_X1 g_37_27 (.ZN (n_37_27), .A (n_38_28), .B (n_44_25), .C1 (n_48_23), .C2 (n_54_20) );
AOI211_X1 g_35_26 (.ZN (n_35_26), .A (n_39_26), .B (n_42_26), .C1 (n_46_24), .C2 (n_52_21) );
AOI211_X1 g_33_27 (.ZN (n_33_27), .A (n_37_27), .B (n_40_27), .C1 (n_44_25), .C2 (n_50_22) );
AOI211_X1 g_31_28 (.ZN (n_31_28), .A (n_35_26), .B (n_38_28), .C1 (n_42_26), .C2 (n_48_23) );
AOI211_X1 g_29_29 (.ZN (n_29_29), .A (n_33_27), .B (n_39_26), .C1 (n_40_27), .C2 (n_46_24) );
AOI211_X1 g_27_30 (.ZN (n_27_30), .A (n_31_28), .B (n_37_27), .C1 (n_38_28), .C2 (n_44_25) );
AOI211_X1 g_26_32 (.ZN (n_26_32), .A (n_29_29), .B (n_35_26), .C1 (n_39_26), .C2 (n_42_26) );
AOI211_X1 g_28_31 (.ZN (n_28_31), .A (n_27_30), .B (n_33_27), .C1 (n_37_27), .C2 (n_40_27) );
AOI211_X1 g_30_30 (.ZN (n_30_30), .A (n_26_32), .B (n_31_28), .C1 (n_35_26), .C2 (n_38_28) );
AOI211_X1 g_32_29 (.ZN (n_32_29), .A (n_28_31), .B (n_29_29), .C1 (n_33_27), .C2 (n_39_26) );
AOI211_X1 g_34_28 (.ZN (n_34_28), .A (n_30_30), .B (n_27_30), .C1 (n_31_28), .C2 (n_37_27) );
AOI211_X1 g_36_29 (.ZN (n_36_29), .A (n_32_29), .B (n_26_32), .C1 (n_29_29), .C2 (n_35_26) );
AOI211_X1 g_34_30 (.ZN (n_34_30), .A (n_34_28), .B (n_28_31), .C1 (n_27_30), .C2 (n_33_27) );
AOI211_X1 g_35_28 (.ZN (n_35_28), .A (n_36_29), .B (n_30_30), .C1 (n_26_32), .C2 (n_31_28) );
AOI211_X1 g_33_29 (.ZN (n_33_29), .A (n_34_30), .B (n_32_29), .C1 (n_28_31), .C2 (n_29_29) );
AOI211_X1 g_32_31 (.ZN (n_32_31), .A (n_35_28), .B (n_34_28), .C1 (n_30_30), .C2 (n_27_30) );
AOI211_X1 g_30_32 (.ZN (n_30_32), .A (n_33_29), .B (n_36_29), .C1 (n_32_29), .C2 (n_26_32) );
AOI211_X1 g_31_30 (.ZN (n_31_30), .A (n_32_31), .B (n_34_30), .C1 (n_34_28), .C2 (n_28_31) );
AOI211_X1 g_32_28 (.ZN (n_32_28), .A (n_30_32), .B (n_35_28), .C1 (n_36_29), .C2 (n_30_30) );
AOI211_X1 g_30_29 (.ZN (n_30_29), .A (n_31_30), .B (n_33_29), .C1 (n_34_30), .C2 (n_32_29) );
AOI211_X1 g_28_30 (.ZN (n_28_30), .A (n_32_28), .B (n_32_31), .C1 (n_35_28), .C2 (n_34_28) );
AOI211_X1 g_26_31 (.ZN (n_26_31), .A (n_30_29), .B (n_30_32), .C1 (n_33_29), .C2 (n_36_29) );
AOI211_X1 g_24_32 (.ZN (n_24_32), .A (n_28_30), .B (n_31_30), .C1 (n_32_31), .C2 (n_34_30) );
AOI211_X1 g_22_33 (.ZN (n_22_33), .A (n_26_31), .B (n_32_28), .C1 (n_30_32), .C2 (n_35_28) );
AOI211_X1 g_20_34 (.ZN (n_20_34), .A (n_24_32), .B (n_30_29), .C1 (n_31_30), .C2 (n_33_29) );
AOI211_X1 g_18_35 (.ZN (n_18_35), .A (n_22_33), .B (n_28_30), .C1 (n_32_28), .C2 (n_32_31) );
AOI211_X1 g_16_36 (.ZN (n_16_36), .A (n_20_34), .B (n_26_31), .C1 (n_30_29), .C2 (n_30_32) );
AOI211_X1 g_14_37 (.ZN (n_14_37), .A (n_18_35), .B (n_24_32), .C1 (n_28_30), .C2 (n_31_30) );
AOI211_X1 g_12_38 (.ZN (n_12_38), .A (n_16_36), .B (n_22_33), .C1 (n_26_31), .C2 (n_32_28) );
AOI211_X1 g_10_39 (.ZN (n_10_39), .A (n_14_37), .B (n_20_34), .C1 (n_24_32), .C2 (n_30_29) );
AOI211_X1 g_9_41 (.ZN (n_9_41), .A (n_12_38), .B (n_18_35), .C1 (n_22_33), .C2 (n_28_30) );
AOI211_X1 g_8_43 (.ZN (n_8_43), .A (n_10_39), .B (n_16_36), .C1 (n_20_34), .C2 (n_26_31) );
AOI211_X1 g_7_45 (.ZN (n_7_45), .A (n_9_41), .B (n_14_37), .C1 (n_18_35), .C2 (n_24_32) );
AOI211_X1 g_6_47 (.ZN (n_6_47), .A (n_8_43), .B (n_12_38), .C1 (n_16_36), .C2 (n_22_33) );
AOI211_X1 g_5_49 (.ZN (n_5_49), .A (n_7_45), .B (n_10_39), .C1 (n_14_37), .C2 (n_20_34) );
AOI211_X1 g_4_51 (.ZN (n_4_51), .A (n_6_47), .B (n_9_41), .C1 (n_12_38), .C2 (n_18_35) );
AOI211_X1 g_6_52 (.ZN (n_6_52), .A (n_5_49), .B (n_8_43), .C1 (n_10_39), .C2 (n_16_36) );
AOI211_X1 g_4_53 (.ZN (n_4_53), .A (n_4_51), .B (n_7_45), .C1 (n_9_41), .C2 (n_14_37) );
AOI211_X1 g_2_54 (.ZN (n_2_54), .A (n_6_52), .B (n_6_47), .C1 (n_8_43), .C2 (n_12_38) );
AOI211_X1 g_3_52 (.ZN (n_3_52), .A (n_4_53), .B (n_5_49), .C1 (n_7_45), .C2 (n_10_39) );
AOI211_X1 g_5_51 (.ZN (n_5_51), .A (n_2_54), .B (n_4_51), .C1 (n_6_47), .C2 (n_9_41) );
AOI211_X1 g_7_50 (.ZN (n_7_50), .A (n_3_52), .B (n_6_52), .C1 (n_5_49), .C2 (n_8_43) );
AOI211_X1 g_8_48 (.ZN (n_8_48), .A (n_5_51), .B (n_4_53), .C1 (n_4_51), .C2 (n_7_45) );
AOI211_X1 g_6_49 (.ZN (n_6_49), .A (n_7_50), .B (n_2_54), .C1 (n_6_52), .C2 (n_6_47) );
AOI211_X1 g_4_50 (.ZN (n_4_50), .A (n_8_48), .B (n_3_52), .C1 (n_4_53), .C2 (n_5_49) );
AOI211_X1 g_5_48 (.ZN (n_5_48), .A (n_6_49), .B (n_5_51), .C1 (n_2_54), .C2 (n_4_51) );
AOI211_X1 g_7_47 (.ZN (n_7_47), .A (n_4_50), .B (n_7_50), .C1 (n_3_52), .C2 (n_6_52) );
AOI211_X1 g_9_46 (.ZN (n_9_46), .A (n_5_48), .B (n_8_48), .C1 (n_5_51), .C2 (n_4_53) );
AOI211_X1 g_10_44 (.ZN (n_10_44), .A (n_7_47), .B (n_6_49), .C1 (n_7_50), .C2 (n_2_54) );
AOI211_X1 g_8_45 (.ZN (n_8_45), .A (n_9_46), .B (n_4_50), .C1 (n_8_48), .C2 (n_3_52) );
AOI211_X1 g_6_46 (.ZN (n_6_46), .A (n_10_44), .B (n_5_48), .C1 (n_6_49), .C2 (n_5_51) );
AOI211_X1 g_7_44 (.ZN (n_7_44), .A (n_8_45), .B (n_7_47), .C1 (n_4_50), .C2 (n_7_50) );
AOI211_X1 g_9_43 (.ZN (n_9_43), .A (n_6_46), .B (n_9_46), .C1 (n_5_48), .C2 (n_8_48) );
AOI211_X1 g_11_42 (.ZN (n_11_42), .A (n_7_44), .B (n_10_44), .C1 (n_7_47), .C2 (n_6_49) );
AOI211_X1 g_12_40 (.ZN (n_12_40), .A (n_9_43), .B (n_8_45), .C1 (n_9_46), .C2 (n_4_50) );
AOI211_X1 g_14_39 (.ZN (n_14_39), .A (n_11_42), .B (n_6_46), .C1 (n_10_44), .C2 (n_5_48) );
AOI211_X1 g_16_38 (.ZN (n_16_38), .A (n_12_40), .B (n_7_44), .C1 (n_8_45), .C2 (n_7_47) );
AOI211_X1 g_18_37 (.ZN (n_18_37), .A (n_14_39), .B (n_9_43), .C1 (n_6_46), .C2 (n_9_46) );
AOI211_X1 g_20_36 (.ZN (n_20_36), .A (n_16_38), .B (n_11_42), .C1 (n_7_44), .C2 (n_10_44) );
AOI211_X1 g_22_35 (.ZN (n_22_35), .A (n_18_37), .B (n_12_40), .C1 (n_9_43), .C2 (n_8_45) );
AOI211_X1 g_24_34 (.ZN (n_24_34), .A (n_20_36), .B (n_14_39), .C1 (n_11_42), .C2 (n_6_46) );
AOI211_X1 g_26_33 (.ZN (n_26_33), .A (n_22_35), .B (n_16_38), .C1 (n_12_40), .C2 (n_7_44) );
AOI211_X1 g_28_32 (.ZN (n_28_32), .A (n_24_34), .B (n_18_37), .C1 (n_14_39), .C2 (n_9_43) );
AOI211_X1 g_30_31 (.ZN (n_30_31), .A (n_26_33), .B (n_20_36), .C1 (n_16_38), .C2 (n_11_42) );
AOI211_X1 g_32_30 (.ZN (n_32_30), .A (n_28_32), .B (n_22_35), .C1 (n_18_37), .C2 (n_12_40) );
AOI211_X1 g_34_29 (.ZN (n_34_29), .A (n_30_31), .B (n_24_34), .C1 (n_20_36), .C2 (n_14_39) );
AOI211_X1 g_36_28 (.ZN (n_36_28), .A (n_32_30), .B (n_26_33), .C1 (n_22_35), .C2 (n_16_38) );
AOI211_X1 g_38_27 (.ZN (n_38_27), .A (n_34_29), .B (n_28_32), .C1 (n_24_34), .C2 (n_18_37) );
AOI211_X1 g_40_26 (.ZN (n_40_26), .A (n_36_28), .B (n_30_31), .C1 (n_26_33), .C2 (n_20_36) );
AOI211_X1 g_39_28 (.ZN (n_39_28), .A (n_38_27), .B (n_32_30), .C1 (n_28_32), .C2 (n_22_35) );
AOI211_X1 g_41_27 (.ZN (n_41_27), .A (n_40_26), .B (n_34_29), .C1 (n_30_31), .C2 (n_24_34) );
AOI211_X1 g_43_26 (.ZN (n_43_26), .A (n_39_28), .B (n_36_28), .C1 (n_32_30), .C2 (n_26_33) );
AOI211_X1 g_45_25 (.ZN (n_45_25), .A (n_41_27), .B (n_38_27), .C1 (n_34_29), .C2 (n_28_32) );
AOI211_X1 g_47_24 (.ZN (n_47_24), .A (n_43_26), .B (n_40_26), .C1 (n_36_28), .C2 (n_30_31) );
AOI211_X1 g_46_26 (.ZN (n_46_26), .A (n_45_25), .B (n_39_28), .C1 (n_38_27), .C2 (n_32_30) );
AOI211_X1 g_48_25 (.ZN (n_48_25), .A (n_47_24), .B (n_41_27), .C1 (n_40_26), .C2 (n_34_29) );
AOI211_X1 g_50_24 (.ZN (n_50_24), .A (n_46_26), .B (n_43_26), .C1 (n_39_28), .C2 (n_36_28) );
AOI211_X1 g_52_23 (.ZN (n_52_23), .A (n_48_25), .B (n_45_25), .C1 (n_41_27), .C2 (n_38_27) );
AOI211_X1 g_54_22 (.ZN (n_54_22), .A (n_50_24), .B (n_47_24), .C1 (n_43_26), .C2 (n_40_26) );
AOI211_X1 g_56_21 (.ZN (n_56_21), .A (n_52_23), .B (n_46_26), .C1 (n_45_25), .C2 (n_39_28) );
AOI211_X1 g_58_20 (.ZN (n_58_20), .A (n_54_22), .B (n_48_25), .C1 (n_47_24), .C2 (n_41_27) );
AOI211_X1 g_60_19 (.ZN (n_60_19), .A (n_56_21), .B (n_50_24), .C1 (n_46_26), .C2 (n_43_26) );
AOI211_X1 g_62_18 (.ZN (n_62_18), .A (n_58_20), .B (n_52_23), .C1 (n_48_25), .C2 (n_45_25) );
AOI211_X1 g_61_20 (.ZN (n_61_20), .A (n_60_19), .B (n_54_22), .C1 (n_50_24), .C2 (n_47_24) );
AOI211_X1 g_59_19 (.ZN (n_59_19), .A (n_62_18), .B (n_56_21), .C1 (n_52_23), .C2 (n_46_26) );
AOI211_X1 g_61_18 (.ZN (n_61_18), .A (n_61_20), .B (n_58_20), .C1 (n_54_22), .C2 (n_48_25) );
AOI211_X1 g_63_17 (.ZN (n_63_17), .A (n_59_19), .B (n_60_19), .C1 (n_56_21), .C2 (n_50_24) );
AOI211_X1 g_65_16 (.ZN (n_65_16), .A (n_61_18), .B (n_62_18), .C1 (n_58_20), .C2 (n_52_23) );
AOI211_X1 g_67_15 (.ZN (n_67_15), .A (n_63_17), .B (n_61_20), .C1 (n_60_19), .C2 (n_54_22) );
AOI211_X1 g_69_14 (.ZN (n_69_14), .A (n_65_16), .B (n_59_19), .C1 (n_62_18), .C2 (n_56_21) );
AOI211_X1 g_71_13 (.ZN (n_71_13), .A (n_67_15), .B (n_61_18), .C1 (n_61_20), .C2 (n_58_20) );
AOI211_X1 g_73_12 (.ZN (n_73_12), .A (n_69_14), .B (n_63_17), .C1 (n_59_19), .C2 (n_60_19) );
AOI211_X1 g_75_11 (.ZN (n_75_11), .A (n_71_13), .B (n_65_16), .C1 (n_61_18), .C2 (n_62_18) );
AOI211_X1 g_77_10 (.ZN (n_77_10), .A (n_73_12), .B (n_67_15), .C1 (n_63_17), .C2 (n_61_20) );
AOI211_X1 g_79_9 (.ZN (n_79_9), .A (n_75_11), .B (n_69_14), .C1 (n_65_16), .C2 (n_59_19) );
AOI211_X1 g_81_8 (.ZN (n_81_8), .A (n_77_10), .B (n_71_13), .C1 (n_67_15), .C2 (n_61_18) );
AOI211_X1 g_83_7 (.ZN (n_83_7), .A (n_79_9), .B (n_73_12), .C1 (n_69_14), .C2 (n_63_17) );
AOI211_X1 g_82_9 (.ZN (n_82_9), .A (n_81_8), .B (n_75_11), .C1 (n_71_13), .C2 (n_65_16) );
AOI211_X1 g_80_10 (.ZN (n_80_10), .A (n_83_7), .B (n_77_10), .C1 (n_73_12), .C2 (n_67_15) );
AOI211_X1 g_78_11 (.ZN (n_78_11), .A (n_82_9), .B (n_79_9), .C1 (n_75_11), .C2 (n_69_14) );
AOI211_X1 g_76_12 (.ZN (n_76_12), .A (n_80_10), .B (n_81_8), .C1 (n_77_10), .C2 (n_71_13) );
AOI211_X1 g_74_13 (.ZN (n_74_13), .A (n_78_11), .B (n_83_7), .C1 (n_79_9), .C2 (n_73_12) );
AOI211_X1 g_72_12 (.ZN (n_72_12), .A (n_76_12), .B (n_82_9), .C1 (n_81_8), .C2 (n_75_11) );
AOI211_X1 g_70_13 (.ZN (n_70_13), .A (n_74_13), .B (n_80_10), .C1 (n_83_7), .C2 (n_77_10) );
AOI211_X1 g_68_14 (.ZN (n_68_14), .A (n_72_12), .B (n_78_11), .C1 (n_82_9), .C2 (n_79_9) );
AOI211_X1 g_66_15 (.ZN (n_66_15), .A (n_70_13), .B (n_76_12), .C1 (n_80_10), .C2 (n_81_8) );
AOI211_X1 g_64_16 (.ZN (n_64_16), .A (n_68_14), .B (n_74_13), .C1 (n_78_11), .C2 (n_83_7) );
AOI211_X1 g_62_17 (.ZN (n_62_17), .A (n_66_15), .B (n_72_12), .C1 (n_76_12), .C2 (n_82_9) );
AOI211_X1 g_63_19 (.ZN (n_63_19), .A (n_64_16), .B (n_70_13), .C1 (n_74_13), .C2 (n_80_10) );
AOI211_X1 g_65_18 (.ZN (n_65_18), .A (n_62_17), .B (n_68_14), .C1 (n_72_12), .C2 (n_78_11) );
AOI211_X1 g_67_17 (.ZN (n_67_17), .A (n_63_19), .B (n_66_15), .C1 (n_70_13), .C2 (n_76_12) );
AOI211_X1 g_69_16 (.ZN (n_69_16), .A (n_65_18), .B (n_64_16), .C1 (n_68_14), .C2 (n_74_13) );
AOI211_X1 g_71_15 (.ZN (n_71_15), .A (n_67_17), .B (n_62_17), .C1 (n_66_15), .C2 (n_72_12) );
AOI211_X1 g_73_14 (.ZN (n_73_14), .A (n_69_16), .B (n_63_19), .C1 (n_64_16), .C2 (n_70_13) );
AOI211_X1 g_75_13 (.ZN (n_75_13), .A (n_71_15), .B (n_65_18), .C1 (n_62_17), .C2 (n_68_14) );
AOI211_X1 g_77_12 (.ZN (n_77_12), .A (n_73_14), .B (n_67_17), .C1 (n_63_19), .C2 (n_66_15) );
AOI211_X1 g_79_11 (.ZN (n_79_11), .A (n_75_13), .B (n_69_16), .C1 (n_65_18), .C2 (n_64_16) );
AOI211_X1 g_80_9 (.ZN (n_80_9), .A (n_77_12), .B (n_71_15), .C1 (n_67_17), .C2 (n_62_17) );
AOI211_X1 g_82_8 (.ZN (n_82_8), .A (n_79_11), .B (n_73_14), .C1 (n_69_16), .C2 (n_63_19) );
AOI211_X1 g_83_6 (.ZN (n_83_6), .A (n_80_9), .B (n_75_13), .C1 (n_71_15), .C2 (n_65_18) );
AOI211_X1 g_85_5 (.ZN (n_85_5), .A (n_82_8), .B (n_77_12), .C1 (n_73_14), .C2 (n_67_17) );
AOI211_X1 g_84_7 (.ZN (n_84_7), .A (n_83_6), .B (n_79_11), .C1 (n_75_13), .C2 (n_69_16) );
AOI211_X1 g_86_6 (.ZN (n_86_6), .A (n_85_5), .B (n_80_9), .C1 (n_77_12), .C2 (n_71_15) );
AOI211_X1 g_88_5 (.ZN (n_88_5), .A (n_84_7), .B (n_82_8), .C1 (n_79_11), .C2 (n_73_14) );
AOI211_X1 g_90_4 (.ZN (n_90_4), .A (n_86_6), .B (n_83_6), .C1 (n_80_9), .C2 (n_75_13) );
AOI211_X1 g_89_6 (.ZN (n_89_6), .A (n_88_5), .B (n_85_5), .C1 (n_82_8), .C2 (n_77_12) );
AOI211_X1 g_91_5 (.ZN (n_91_5), .A (n_90_4), .B (n_84_7), .C1 (n_83_6), .C2 (n_79_11) );
AOI211_X1 g_93_4 (.ZN (n_93_4), .A (n_89_6), .B (n_86_6), .C1 (n_85_5), .C2 (n_80_9) );
AOI211_X1 g_92_6 (.ZN (n_92_6), .A (n_91_5), .B (n_88_5), .C1 (n_84_7), .C2 (n_82_8) );
AOI211_X1 g_90_5 (.ZN (n_90_5), .A (n_93_4), .B (n_90_4), .C1 (n_86_6), .C2 (n_83_6) );
AOI211_X1 g_92_4 (.ZN (n_92_4), .A (n_92_6), .B (n_89_6), .C1 (n_88_5), .C2 (n_85_5) );
AOI211_X1 g_94_3 (.ZN (n_94_3), .A (n_90_5), .B (n_91_5), .C1 (n_90_4), .C2 (n_84_7) );
AOI211_X1 g_96_2 (.ZN (n_96_2), .A (n_92_4), .B (n_93_4), .C1 (n_89_6), .C2 (n_86_6) );
AOI211_X1 g_97_4 (.ZN (n_97_4), .A (n_94_3), .B (n_92_6), .C1 (n_91_5), .C2 (n_88_5) );
AOI211_X1 g_99_5 (.ZN (n_99_5), .A (n_96_2), .B (n_90_5), .C1 (n_93_4), .C2 (n_90_4) );
AOI211_X1 g_100_7 (.ZN (n_100_7), .A (n_97_4), .B (n_92_4), .C1 (n_92_6), .C2 (n_89_6) );
AOI211_X1 g_98_6 (.ZN (n_98_6), .A (n_99_5), .B (n_94_3), .C1 (n_90_5), .C2 (n_91_5) );
AOI211_X1 g_100_5 (.ZN (n_100_5), .A (n_100_7), .B (n_96_2), .C1 (n_92_4), .C2 (n_93_4) );
AOI211_X1 g_98_4 (.ZN (n_98_4), .A (n_98_6), .B (n_97_4), .C1 (n_94_3), .C2 (n_92_6) );
AOI211_X1 g_99_2 (.ZN (n_99_2), .A (n_100_5), .B (n_99_5), .C1 (n_96_2), .C2 (n_90_5) );
AOI211_X1 g_97_1 (.ZN (n_97_1), .A (n_98_4), .B (n_100_7), .C1 (n_97_4), .C2 (n_92_4) );
AOI211_X1 g_96_3 (.ZN (n_96_3), .A (n_99_2), .B (n_98_6), .C1 (n_99_5), .C2 (n_94_3) );
AOI211_X1 g_95_5 (.ZN (n_95_5), .A (n_97_1), .B (n_100_5), .C1 (n_100_7), .C2 (n_96_2) );
AOI211_X1 g_93_6 (.ZN (n_93_6), .A (n_96_3), .B (n_98_4), .C1 (n_98_6), .C2 (n_97_4) );
AOI211_X1 g_94_4 (.ZN (n_94_4), .A (n_95_5), .B (n_99_2), .C1 (n_100_5), .C2 (n_99_5) );
AOI211_X1 g_95_2 (.ZN (n_95_2), .A (n_93_6), .B (n_97_1), .C1 (n_98_4), .C2 (n_100_7) );
AOI211_X1 g_97_3 (.ZN (n_97_3), .A (n_94_4), .B (n_96_3), .C1 (n_99_2), .C2 (n_98_6) );
AOI211_X1 g_96_5 (.ZN (n_96_5), .A (n_95_2), .B (n_95_5), .C1 (n_97_1), .C2 (n_100_5) );
AOI211_X1 g_94_6 (.ZN (n_94_6), .A (n_97_3), .B (n_93_6), .C1 (n_96_3), .C2 (n_98_4) );
AOI211_X1 g_95_4 (.ZN (n_95_4), .A (n_96_5), .B (n_94_4), .C1 (n_95_5), .C2 (n_99_2) );
AOI211_X1 g_93_3 (.ZN (n_93_3), .A (n_94_6), .B (n_95_2), .C1 (n_93_6), .C2 (n_97_1) );
AOI211_X1 g_91_4 (.ZN (n_91_4), .A (n_95_4), .B (n_97_3), .C1 (n_94_4), .C2 (n_96_3) );
AOI211_X1 g_89_5 (.ZN (n_89_5), .A (n_93_3), .B (n_96_5), .C1 (n_95_2), .C2 (n_95_5) );
AOI211_X1 g_87_6 (.ZN (n_87_6), .A (n_91_4), .B (n_94_6), .C1 (n_97_3), .C2 (n_93_6) );
AOI211_X1 g_85_7 (.ZN (n_85_7), .A (n_89_5), .B (n_95_4), .C1 (n_96_5), .C2 (n_94_4) );
AOI211_X1 g_83_8 (.ZN (n_83_8), .A (n_87_6), .B (n_93_3), .C1 (n_94_6), .C2 (n_95_2) );
AOI211_X1 g_81_9 (.ZN (n_81_9), .A (n_85_7), .B (n_91_4), .C1 (n_95_4), .C2 (n_97_3) );
AOI211_X1 g_79_10 (.ZN (n_79_10), .A (n_83_8), .B (n_89_5), .C1 (n_93_3), .C2 (n_96_5) );
AOI211_X1 g_77_11 (.ZN (n_77_11), .A (n_81_9), .B (n_87_6), .C1 (n_91_4), .C2 (n_94_6) );
AOI211_X1 g_75_12 (.ZN (n_75_12), .A (n_79_10), .B (n_85_7), .C1 (n_89_5), .C2 (n_95_4) );
AOI211_X1 g_73_13 (.ZN (n_73_13), .A (n_77_11), .B (n_83_8), .C1 (n_87_6), .C2 (n_93_3) );
AOI211_X1 g_71_14 (.ZN (n_71_14), .A (n_75_12), .B (n_81_9), .C1 (n_85_7), .C2 (n_91_4) );
AOI211_X1 g_69_15 (.ZN (n_69_15), .A (n_73_13), .B (n_79_10), .C1 (n_83_8), .C2 (n_89_5) );
AOI211_X1 g_67_16 (.ZN (n_67_16), .A (n_71_14), .B (n_77_11), .C1 (n_81_9), .C2 (n_87_6) );
AOI211_X1 g_65_17 (.ZN (n_65_17), .A (n_69_15), .B (n_75_12), .C1 (n_79_10), .C2 (n_85_7) );
AOI211_X1 g_63_18 (.ZN (n_63_18), .A (n_67_16), .B (n_73_13), .C1 (n_77_11), .C2 (n_83_8) );
AOI211_X1 g_61_19 (.ZN (n_61_19), .A (n_65_17), .B (n_71_14), .C1 (n_75_12), .C2 (n_81_9) );
AOI211_X1 g_59_20 (.ZN (n_59_20), .A (n_63_18), .B (n_69_15), .C1 (n_73_13), .C2 (n_79_10) );
AOI211_X1 g_57_21 (.ZN (n_57_21), .A (n_61_19), .B (n_67_16), .C1 (n_71_14), .C2 (n_77_11) );
AOI211_X1 g_55_22 (.ZN (n_55_22), .A (n_59_20), .B (n_65_17), .C1 (n_69_15), .C2 (n_75_12) );
AOI211_X1 g_53_23 (.ZN (n_53_23), .A (n_57_21), .B (n_63_18), .C1 (n_67_16), .C2 (n_73_13) );
AOI211_X1 g_54_21 (.ZN (n_54_21), .A (n_55_22), .B (n_61_19), .C1 (n_65_17), .C2 (n_71_14) );
AOI211_X1 g_52_22 (.ZN (n_52_22), .A (n_53_23), .B (n_59_20), .C1 (n_63_18), .C2 (n_69_15) );
AOI211_X1 g_50_23 (.ZN (n_50_23), .A (n_54_21), .B (n_57_21), .C1 (n_61_19), .C2 (n_67_16) );
AOI211_X1 g_48_24 (.ZN (n_48_24), .A (n_52_22), .B (n_55_22), .C1 (n_59_20), .C2 (n_65_17) );
AOI211_X1 g_46_25 (.ZN (n_46_25), .A (n_50_23), .B (n_53_23), .C1 (n_57_21), .C2 (n_63_18) );
AOI211_X1 g_44_26 (.ZN (n_44_26), .A (n_48_24), .B (n_54_21), .C1 (n_55_22), .C2 (n_61_19) );
AOI211_X1 g_42_27 (.ZN (n_42_27), .A (n_46_25), .B (n_52_22), .C1 (n_53_23), .C2 (n_59_20) );
AOI211_X1 g_40_28 (.ZN (n_40_28), .A (n_44_26), .B (n_50_23), .C1 (n_54_21), .C2 (n_57_21) );
AOI211_X1 g_38_29 (.ZN (n_38_29), .A (n_42_27), .B (n_48_24), .C1 (n_52_22), .C2 (n_55_22) );
AOI211_X1 g_39_27 (.ZN (n_39_27), .A (n_40_28), .B (n_46_25), .C1 (n_50_23), .C2 (n_53_23) );
AOI211_X1 g_37_28 (.ZN (n_37_28), .A (n_38_29), .B (n_44_26), .C1 (n_48_24), .C2 (n_54_21) );
AOI211_X1 g_36_30 (.ZN (n_36_30), .A (n_39_27), .B (n_42_27), .C1 (n_46_25), .C2 (n_52_22) );
AOI211_X1 g_34_31 (.ZN (n_34_31), .A (n_37_28), .B (n_40_28), .C1 (n_44_26), .C2 (n_50_23) );
AOI211_X1 g_32_32 (.ZN (n_32_32), .A (n_36_30), .B (n_38_29), .C1 (n_42_27), .C2 (n_48_24) );
AOI211_X1 g_33_30 (.ZN (n_33_30), .A (n_34_31), .B (n_39_27), .C1 (n_40_28), .C2 (n_46_25) );
AOI211_X1 g_31_31 (.ZN (n_31_31), .A (n_32_32), .B (n_37_28), .C1 (n_38_29), .C2 (n_44_26) );
AOI211_X1 g_29_32 (.ZN (n_29_32), .A (n_33_30), .B (n_36_30), .C1 (n_39_27), .C2 (n_42_27) );
AOI211_X1 g_27_33 (.ZN (n_27_33), .A (n_31_31), .B (n_34_31), .C1 (n_37_28), .C2 (n_40_28) );
AOI211_X1 g_25_34 (.ZN (n_25_34), .A (n_29_32), .B (n_32_32), .C1 (n_36_30), .C2 (n_38_29) );
AOI211_X1 g_23_35 (.ZN (n_23_35), .A (n_27_33), .B (n_33_30), .C1 (n_34_31), .C2 (n_39_27) );
AOI211_X1 g_24_33 (.ZN (n_24_33), .A (n_25_34), .B (n_31_31), .C1 (n_32_32), .C2 (n_37_28) );
AOI211_X1 g_22_34 (.ZN (n_22_34), .A (n_23_35), .B (n_29_32), .C1 (n_33_30), .C2 (n_36_30) );
AOI211_X1 g_21_36 (.ZN (n_21_36), .A (n_24_33), .B (n_27_33), .C1 (n_31_31), .C2 (n_34_31) );
AOI211_X1 g_19_37 (.ZN (n_19_37), .A (n_22_34), .B (n_25_34), .C1 (n_29_32), .C2 (n_32_32) );
AOI211_X1 g_17_38 (.ZN (n_17_38), .A (n_21_36), .B (n_23_35), .C1 (n_27_33), .C2 (n_33_30) );
AOI211_X1 g_15_39 (.ZN (n_15_39), .A (n_19_37), .B (n_24_33), .C1 (n_25_34), .C2 (n_31_31) );
AOI211_X1 g_13_40 (.ZN (n_13_40), .A (n_17_38), .B (n_22_34), .C1 (n_23_35), .C2 (n_29_32) );
AOI211_X1 g_14_38 (.ZN (n_14_38), .A (n_15_39), .B (n_21_36), .C1 (n_24_33), .C2 (n_27_33) );
AOI211_X1 g_12_39 (.ZN (n_12_39), .A (n_13_40), .B (n_19_37), .C1 (n_22_34), .C2 (n_25_34) );
AOI211_X1 g_10_38 (.ZN (n_10_38), .A (n_14_38), .B (n_17_38), .C1 (n_21_36), .C2 (n_23_35) );
AOI211_X1 g_9_40 (.ZN (n_9_40), .A (n_12_39), .B (n_15_39), .C1 (n_19_37), .C2 (n_24_33) );
AOI211_X1 g_11_39 (.ZN (n_11_39), .A (n_10_38), .B (n_13_40), .C1 (n_17_38), .C2 (n_22_34) );
AOI211_X1 g_10_41 (.ZN (n_10_41), .A (n_9_40), .B (n_14_38), .C1 (n_15_39), .C2 (n_21_36) );
AOI211_X1 g_8_42 (.ZN (n_8_42), .A (n_11_39), .B (n_12_39), .C1 (n_13_40), .C2 (n_19_37) );
AOI211_X1 g_9_44 (.ZN (n_9_44), .A (n_10_41), .B (n_10_38), .C1 (n_14_38), .C2 (n_17_38) );
AOI211_X1 g_10_42 (.ZN (n_10_42), .A (n_8_42), .B (n_9_40), .C1 (n_12_39), .C2 (n_15_39) );
AOI211_X1 g_11_40 (.ZN (n_11_40), .A (n_9_44), .B (n_11_39), .C1 (n_10_38), .C2 (n_13_40) );
AOI211_X1 g_13_39 (.ZN (n_13_39), .A (n_10_42), .B (n_10_41), .C1 (n_9_40), .C2 (n_14_38) );
AOI211_X1 g_15_38 (.ZN (n_15_38), .A (n_11_40), .B (n_8_42), .C1 (n_11_39), .C2 (n_12_39) );
AOI211_X1 g_17_37 (.ZN (n_17_37), .A (n_13_39), .B (n_9_44), .C1 (n_10_41), .C2 (n_10_38) );
AOI211_X1 g_19_36 (.ZN (n_19_36), .A (n_15_38), .B (n_10_42), .C1 (n_8_42), .C2 (n_9_40) );
AOI211_X1 g_21_35 (.ZN (n_21_35), .A (n_17_37), .B (n_11_40), .C1 (n_9_44), .C2 (n_11_39) );
AOI211_X1 g_23_34 (.ZN (n_23_34), .A (n_19_36), .B (n_13_39), .C1 (n_10_42), .C2 (n_10_41) );
AOI211_X1 g_25_33 (.ZN (n_25_33), .A (n_21_35), .B (n_15_38), .C1 (n_11_40), .C2 (n_8_42) );
AOI211_X1 g_27_32 (.ZN (n_27_32), .A (n_23_34), .B (n_17_37), .C1 (n_13_39), .C2 (n_9_44) );
AOI211_X1 g_29_31 (.ZN (n_29_31), .A (n_25_33), .B (n_19_36), .C1 (n_15_38), .C2 (n_10_42) );
AOI211_X1 g_28_33 (.ZN (n_28_33), .A (n_27_32), .B (n_21_35), .C1 (n_17_37), .C2 (n_11_40) );
AOI211_X1 g_26_34 (.ZN (n_26_34), .A (n_29_31), .B (n_23_34), .C1 (n_19_36), .C2 (n_13_39) );
AOI211_X1 g_24_35 (.ZN (n_24_35), .A (n_28_33), .B (n_25_33), .C1 (n_21_35), .C2 (n_15_38) );
AOI211_X1 g_22_36 (.ZN (n_22_36), .A (n_26_34), .B (n_27_32), .C1 (n_23_34), .C2 (n_17_37) );
AOI211_X1 g_20_37 (.ZN (n_20_37), .A (n_24_35), .B (n_29_31), .C1 (n_25_33), .C2 (n_19_36) );
AOI211_X1 g_18_38 (.ZN (n_18_38), .A (n_22_36), .B (n_28_33), .C1 (n_27_32), .C2 (n_21_35) );
AOI211_X1 g_16_39 (.ZN (n_16_39), .A (n_20_37), .B (n_26_34), .C1 (n_29_31), .C2 (n_23_34) );
AOI211_X1 g_14_40 (.ZN (n_14_40), .A (n_18_38), .B (n_24_35), .C1 (n_28_33), .C2 (n_25_33) );
AOI211_X1 g_12_41 (.ZN (n_12_41), .A (n_16_39), .B (n_22_36), .C1 (n_26_34), .C2 (n_27_32) );
AOI211_X1 g_11_43 (.ZN (n_11_43), .A (n_14_40), .B (n_20_37), .C1 (n_24_35), .C2 (n_29_31) );
AOI211_X1 g_13_42 (.ZN (n_13_42), .A (n_12_41), .B (n_18_38), .C1 (n_22_36), .C2 (n_28_33) );
AOI211_X1 g_11_41 (.ZN (n_11_41), .A (n_11_43), .B (n_16_39), .C1 (n_20_37), .C2 (n_26_34) );
AOI211_X1 g_10_43 (.ZN (n_10_43), .A (n_13_42), .B (n_14_40), .C1 (n_18_38), .C2 (n_24_35) );
AOI211_X1 g_12_42 (.ZN (n_12_42), .A (n_11_41), .B (n_12_41), .C1 (n_16_39), .C2 (n_22_36) );
AOI211_X1 g_14_41 (.ZN (n_14_41), .A (n_10_43), .B (n_11_43), .C1 (n_14_40), .C2 (n_20_37) );
AOI211_X1 g_16_40 (.ZN (n_16_40), .A (n_12_42), .B (n_13_42), .C1 (n_12_41), .C2 (n_18_38) );
AOI211_X1 g_18_39 (.ZN (n_18_39), .A (n_14_41), .B (n_11_41), .C1 (n_11_43), .C2 (n_16_39) );
AOI211_X1 g_20_38 (.ZN (n_20_38), .A (n_16_40), .B (n_10_43), .C1 (n_13_42), .C2 (n_14_40) );
AOI211_X1 g_22_37 (.ZN (n_22_37), .A (n_18_39), .B (n_12_42), .C1 (n_11_41), .C2 (n_12_41) );
AOI211_X1 g_24_36 (.ZN (n_24_36), .A (n_20_38), .B (n_14_41), .C1 (n_10_43), .C2 (n_11_43) );
AOI211_X1 g_26_35 (.ZN (n_26_35), .A (n_22_37), .B (n_16_40), .C1 (n_12_42), .C2 (n_13_42) );
AOI211_X1 g_28_34 (.ZN (n_28_34), .A (n_24_36), .B (n_18_39), .C1 (n_14_41), .C2 (n_11_41) );
AOI211_X1 g_30_33 (.ZN (n_30_33), .A (n_26_35), .B (n_20_38), .C1 (n_16_40), .C2 (n_10_43) );
AOI211_X1 g_29_35 (.ZN (n_29_35), .A (n_28_34), .B (n_22_37), .C1 (n_18_39), .C2 (n_12_42) );
AOI211_X1 g_27_34 (.ZN (n_27_34), .A (n_30_33), .B (n_24_36), .C1 (n_20_38), .C2 (n_14_41) );
AOI211_X1 g_29_33 (.ZN (n_29_33), .A (n_29_35), .B (n_26_35), .C1 (n_22_37), .C2 (n_16_40) );
AOI211_X1 g_31_32 (.ZN (n_31_32), .A (n_27_34), .B (n_28_34), .C1 (n_24_36), .C2 (n_18_39) );
AOI211_X1 g_33_31 (.ZN (n_33_31), .A (n_29_33), .B (n_30_33), .C1 (n_26_35), .C2 (n_20_38) );
AOI211_X1 g_35_30 (.ZN (n_35_30), .A (n_31_32), .B (n_29_35), .C1 (n_28_34), .C2 (n_22_37) );
AOI211_X1 g_37_29 (.ZN (n_37_29), .A (n_33_31), .B (n_27_34), .C1 (n_30_33), .C2 (n_24_36) );
AOI211_X1 g_36_31 (.ZN (n_36_31), .A (n_35_30), .B (n_29_33), .C1 (n_29_35), .C2 (n_26_35) );
AOI211_X1 g_38_30 (.ZN (n_38_30), .A (n_37_29), .B (n_31_32), .C1 (n_27_34), .C2 (n_28_34) );
AOI211_X1 g_40_29 (.ZN (n_40_29), .A (n_36_31), .B (n_33_31), .C1 (n_29_33), .C2 (n_30_33) );
AOI211_X1 g_42_28 (.ZN (n_42_28), .A (n_38_30), .B (n_35_30), .C1 (n_31_32), .C2 (n_29_35) );
AOI211_X1 g_44_27 (.ZN (n_44_27), .A (n_40_29), .B (n_37_29), .C1 (n_33_31), .C2 (n_27_34) );
AOI211_X1 g_43_29 (.ZN (n_43_29), .A (n_42_28), .B (n_36_31), .C1 (n_35_30), .C2 (n_29_33) );
AOI211_X1 g_41_28 (.ZN (n_41_28), .A (n_44_27), .B (n_38_30), .C1 (n_37_29), .C2 (n_31_32) );
AOI211_X1 g_43_27 (.ZN (n_43_27), .A (n_43_29), .B (n_40_29), .C1 (n_36_31), .C2 (n_33_31) );
AOI211_X1 g_45_26 (.ZN (n_45_26), .A (n_41_28), .B (n_42_28), .C1 (n_38_30), .C2 (n_35_30) );
AOI211_X1 g_47_25 (.ZN (n_47_25), .A (n_43_27), .B (n_44_27), .C1 (n_40_29), .C2 (n_37_29) );
AOI211_X1 g_49_24 (.ZN (n_49_24), .A (n_45_26), .B (n_43_29), .C1 (n_42_28), .C2 (n_36_31) );
AOI211_X1 g_51_23 (.ZN (n_51_23), .A (n_47_25), .B (n_41_28), .C1 (n_44_27), .C2 (n_38_30) );
AOI211_X1 g_53_22 (.ZN (n_53_22), .A (n_49_24), .B (n_43_27), .C1 (n_43_29), .C2 (n_40_29) );
AOI211_X1 g_55_21 (.ZN (n_55_21), .A (n_51_23), .B (n_45_26), .C1 (n_41_28), .C2 (n_42_28) );
AOI211_X1 g_57_20 (.ZN (n_57_20), .A (n_53_22), .B (n_47_25), .C1 (n_43_27), .C2 (n_44_27) );
AOI211_X1 g_59_21 (.ZN (n_59_21), .A (n_55_21), .B (n_49_24), .C1 (n_45_26), .C2 (n_43_29) );
AOI211_X1 g_57_22 (.ZN (n_57_22), .A (n_57_20), .B (n_51_23), .C1 (n_47_25), .C2 (n_41_28) );
AOI211_X1 g_55_23 (.ZN (n_55_23), .A (n_59_21), .B (n_53_22), .C1 (n_49_24), .C2 (n_43_27) );
AOI211_X1 g_53_24 (.ZN (n_53_24), .A (n_57_22), .B (n_55_21), .C1 (n_51_23), .C2 (n_45_26) );
AOI211_X1 g_51_25 (.ZN (n_51_25), .A (n_55_23), .B (n_57_20), .C1 (n_53_22), .C2 (n_47_25) );
AOI211_X1 g_49_26 (.ZN (n_49_26), .A (n_53_24), .B (n_59_21), .C1 (n_55_21), .C2 (n_49_24) );
AOI211_X1 g_47_27 (.ZN (n_47_27), .A (n_51_25), .B (n_57_22), .C1 (n_57_20), .C2 (n_51_23) );
AOI211_X1 g_45_28 (.ZN (n_45_28), .A (n_49_26), .B (n_55_23), .C1 (n_59_21), .C2 (n_53_22) );
AOI211_X1 g_44_30 (.ZN (n_44_30), .A (n_47_27), .B (n_53_24), .C1 (n_57_22), .C2 (n_55_21) );
AOI211_X1 g_43_28 (.ZN (n_43_28), .A (n_45_28), .B (n_51_25), .C1 (n_55_23), .C2 (n_57_20) );
AOI211_X1 g_45_27 (.ZN (n_45_27), .A (n_44_30), .B (n_49_26), .C1 (n_53_24), .C2 (n_59_21) );
AOI211_X1 g_47_26 (.ZN (n_47_26), .A (n_43_28), .B (n_47_27), .C1 (n_51_25), .C2 (n_57_22) );
AOI211_X1 g_49_25 (.ZN (n_49_25), .A (n_45_27), .B (n_45_28), .C1 (n_49_26), .C2 (n_55_23) );
AOI211_X1 g_51_24 (.ZN (n_51_24), .A (n_47_26), .B (n_44_30), .C1 (n_47_27), .C2 (n_53_24) );
AOI211_X1 g_50_26 (.ZN (n_50_26), .A (n_49_25), .B (n_43_28), .C1 (n_45_28), .C2 (n_51_25) );
AOI211_X1 g_52_25 (.ZN (n_52_25), .A (n_51_24), .B (n_45_27), .C1 (n_44_30), .C2 (n_49_26) );
AOI211_X1 g_54_24 (.ZN (n_54_24), .A (n_50_26), .B (n_47_26), .C1 (n_43_28), .C2 (n_47_27) );
AOI211_X1 g_56_23 (.ZN (n_56_23), .A (n_52_25), .B (n_49_25), .C1 (n_45_27), .C2 (n_45_28) );
AOI211_X1 g_58_22 (.ZN (n_58_22), .A (n_54_24), .B (n_51_24), .C1 (n_47_26), .C2 (n_44_30) );
AOI211_X1 g_60_21 (.ZN (n_60_21), .A (n_56_23), .B (n_50_26), .C1 (n_49_25), .C2 (n_43_28) );
AOI211_X1 g_62_20 (.ZN (n_62_20), .A (n_58_22), .B (n_52_25), .C1 (n_51_24), .C2 (n_45_27) );
AOI211_X1 g_64_19 (.ZN (n_64_19), .A (n_60_21), .B (n_54_24), .C1 (n_50_26), .C2 (n_47_26) );
AOI211_X1 g_66_18 (.ZN (n_66_18), .A (n_62_20), .B (n_56_23), .C1 (n_52_25), .C2 (n_49_25) );
AOI211_X1 g_68_17 (.ZN (n_68_17), .A (n_64_19), .B (n_58_22), .C1 (n_54_24), .C2 (n_51_24) );
AOI211_X1 g_70_16 (.ZN (n_70_16), .A (n_66_18), .B (n_60_21), .C1 (n_56_23), .C2 (n_50_26) );
AOI211_X1 g_72_15 (.ZN (n_72_15), .A (n_68_17), .B (n_62_20), .C1 (n_58_22), .C2 (n_52_25) );
AOI211_X1 g_74_14 (.ZN (n_74_14), .A (n_70_16), .B (n_64_19), .C1 (n_60_21), .C2 (n_54_24) );
AOI211_X1 g_76_13 (.ZN (n_76_13), .A (n_72_15), .B (n_66_18), .C1 (n_62_20), .C2 (n_56_23) );
AOI211_X1 g_78_12 (.ZN (n_78_12), .A (n_74_14), .B (n_68_17), .C1 (n_64_19), .C2 (n_58_22) );
AOI211_X1 g_80_11 (.ZN (n_80_11), .A (n_76_13), .B (n_70_16), .C1 (n_66_18), .C2 (n_60_21) );
AOI211_X1 g_82_10 (.ZN (n_82_10), .A (n_78_12), .B (n_72_15), .C1 (n_68_17), .C2 (n_62_20) );
AOI211_X1 g_84_9 (.ZN (n_84_9), .A (n_80_11), .B (n_74_14), .C1 (n_70_16), .C2 (n_64_19) );
AOI211_X1 g_86_8 (.ZN (n_86_8), .A (n_82_10), .B (n_76_13), .C1 (n_72_15), .C2 (n_66_18) );
AOI211_X1 g_88_7 (.ZN (n_88_7), .A (n_84_9), .B (n_78_12), .C1 (n_74_14), .C2 (n_68_17) );
AOI211_X1 g_90_6 (.ZN (n_90_6), .A (n_86_8), .B (n_80_11), .C1 (n_76_13), .C2 (n_70_16) );
AOI211_X1 g_92_5 (.ZN (n_92_5), .A (n_88_7), .B (n_82_10), .C1 (n_78_12), .C2 (n_72_15) );
AOI211_X1 g_91_7 (.ZN (n_91_7), .A (n_90_6), .B (n_84_9), .C1 (n_80_11), .C2 (n_74_14) );
AOI211_X1 g_89_8 (.ZN (n_89_8), .A (n_92_5), .B (n_86_8), .C1 (n_82_10), .C2 (n_76_13) );
AOI211_X1 g_87_7 (.ZN (n_87_7), .A (n_91_7), .B (n_88_7), .C1 (n_84_9), .C2 (n_78_12) );
AOI211_X1 g_85_8 (.ZN (n_85_8), .A (n_89_8), .B (n_90_6), .C1 (n_86_8), .C2 (n_80_11) );
AOI211_X1 g_83_9 (.ZN (n_83_9), .A (n_87_7), .B (n_92_5), .C1 (n_88_7), .C2 (n_82_10) );
AOI211_X1 g_81_10 (.ZN (n_81_10), .A (n_85_8), .B (n_91_7), .C1 (n_90_6), .C2 (n_84_9) );
AOI211_X1 g_80_12 (.ZN (n_80_12), .A (n_83_9), .B (n_89_8), .C1 (n_92_5), .C2 (n_86_8) );
AOI211_X1 g_82_11 (.ZN (n_82_11), .A (n_81_10), .B (n_87_7), .C1 (n_91_7), .C2 (n_88_7) );
AOI211_X1 g_84_10 (.ZN (n_84_10), .A (n_80_12), .B (n_85_8), .C1 (n_89_8), .C2 (n_90_6) );
AOI211_X1 g_86_9 (.ZN (n_86_9), .A (n_82_11), .B (n_83_9), .C1 (n_87_7), .C2 (n_92_5) );
AOI211_X1 g_84_8 (.ZN (n_84_8), .A (n_84_10), .B (n_81_10), .C1 (n_85_8), .C2 (n_91_7) );
AOI211_X1 g_86_7 (.ZN (n_86_7), .A (n_86_9), .B (n_80_12), .C1 (n_83_9), .C2 (n_89_8) );
AOI211_X1 g_87_9 (.ZN (n_87_9), .A (n_84_8), .B (n_82_11), .C1 (n_81_10), .C2 (n_87_7) );
AOI211_X1 g_85_10 (.ZN (n_85_10), .A (n_86_7), .B (n_84_10), .C1 (n_80_12), .C2 (n_85_8) );
AOI211_X1 g_83_11 (.ZN (n_83_11), .A (n_87_9), .B (n_86_9), .C1 (n_82_11), .C2 (n_83_9) );
AOI211_X1 g_81_12 (.ZN (n_81_12), .A (n_85_10), .B (n_84_8), .C1 (n_84_10), .C2 (n_81_10) );
AOI211_X1 g_79_13 (.ZN (n_79_13), .A (n_83_11), .B (n_86_7), .C1 (n_86_9), .C2 (n_80_12) );
AOI211_X1 g_77_14 (.ZN (n_77_14), .A (n_81_12), .B (n_87_9), .C1 (n_84_8), .C2 (n_82_11) );
AOI211_X1 g_75_15 (.ZN (n_75_15), .A (n_79_13), .B (n_85_10), .C1 (n_86_7), .C2 (n_84_10) );
AOI211_X1 g_73_16 (.ZN (n_73_16), .A (n_77_14), .B (n_83_11), .C1 (n_87_9), .C2 (n_86_9) );
AOI211_X1 g_72_14 (.ZN (n_72_14), .A (n_75_15), .B (n_81_12), .C1 (n_85_10), .C2 (n_84_8) );
AOI211_X1 g_70_15 (.ZN (n_70_15), .A (n_73_16), .B (n_79_13), .C1 (n_83_11), .C2 (n_86_7) );
AOI211_X1 g_68_16 (.ZN (n_68_16), .A (n_72_14), .B (n_77_14), .C1 (n_81_12), .C2 (n_87_9) );
AOI211_X1 g_66_17 (.ZN (n_66_17), .A (n_70_15), .B (n_75_15), .C1 (n_79_13), .C2 (n_85_10) );
AOI211_X1 g_64_18 (.ZN (n_64_18), .A (n_68_16), .B (n_73_16), .C1 (n_77_14), .C2 (n_83_11) );
AOI211_X1 g_62_19 (.ZN (n_62_19), .A (n_66_17), .B (n_72_14), .C1 (n_75_15), .C2 (n_81_12) );
AOI211_X1 g_60_20 (.ZN (n_60_20), .A (n_64_18), .B (n_70_15), .C1 (n_73_16), .C2 (n_79_13) );
AOI211_X1 g_58_21 (.ZN (n_58_21), .A (n_62_19), .B (n_68_16), .C1 (n_72_14), .C2 (n_77_14) );
AOI211_X1 g_56_22 (.ZN (n_56_22), .A (n_60_20), .B (n_66_17), .C1 (n_70_15), .C2 (n_75_15) );
AOI211_X1 g_54_23 (.ZN (n_54_23), .A (n_58_21), .B (n_64_18), .C1 (n_68_16), .C2 (n_73_16) );
AOI211_X1 g_52_24 (.ZN (n_52_24), .A (n_56_22), .B (n_62_19), .C1 (n_66_17), .C2 (n_72_14) );
AOI211_X1 g_50_25 (.ZN (n_50_25), .A (n_54_23), .B (n_60_20), .C1 (n_64_18), .C2 (n_70_15) );
AOI211_X1 g_48_26 (.ZN (n_48_26), .A (n_52_24), .B (n_58_21), .C1 (n_62_19), .C2 (n_68_16) );
AOI211_X1 g_46_27 (.ZN (n_46_27), .A (n_50_25), .B (n_56_22), .C1 (n_60_20), .C2 (n_66_17) );
AOI211_X1 g_44_28 (.ZN (n_44_28), .A (n_48_26), .B (n_54_23), .C1 (n_58_21), .C2 (n_64_18) );
AOI211_X1 g_42_29 (.ZN (n_42_29), .A (n_46_27), .B (n_52_24), .C1 (n_56_22), .C2 (n_62_19) );
AOI211_X1 g_40_30 (.ZN (n_40_30), .A (n_44_28), .B (n_50_25), .C1 (n_54_23), .C2 (n_60_20) );
AOI211_X1 g_38_31 (.ZN (n_38_31), .A (n_42_29), .B (n_48_26), .C1 (n_52_24), .C2 (n_58_21) );
AOI211_X1 g_39_29 (.ZN (n_39_29), .A (n_40_30), .B (n_46_27), .C1 (n_50_25), .C2 (n_56_22) );
AOI211_X1 g_37_30 (.ZN (n_37_30), .A (n_38_31), .B (n_44_28), .C1 (n_48_26), .C2 (n_54_23) );
AOI211_X1 g_35_31 (.ZN (n_35_31), .A (n_39_29), .B (n_42_29), .C1 (n_46_27), .C2 (n_52_24) );
AOI211_X1 g_33_32 (.ZN (n_33_32), .A (n_37_30), .B (n_40_30), .C1 (n_44_28), .C2 (n_50_25) );
AOI211_X1 g_31_33 (.ZN (n_31_33), .A (n_35_31), .B (n_38_31), .C1 (n_42_29), .C2 (n_48_26) );
AOI211_X1 g_29_34 (.ZN (n_29_34), .A (n_33_32), .B (n_39_29), .C1 (n_40_30), .C2 (n_46_27) );
AOI211_X1 g_27_35 (.ZN (n_27_35), .A (n_31_33), .B (n_37_30), .C1 (n_38_31), .C2 (n_44_28) );
AOI211_X1 g_25_36 (.ZN (n_25_36), .A (n_29_34), .B (n_35_31), .C1 (n_39_29), .C2 (n_42_29) );
AOI211_X1 g_23_37 (.ZN (n_23_37), .A (n_27_35), .B (n_33_32), .C1 (n_37_30), .C2 (n_40_30) );
AOI211_X1 g_21_38 (.ZN (n_21_38), .A (n_25_36), .B (n_31_33), .C1 (n_35_31), .C2 (n_38_31) );
AOI211_X1 g_19_39 (.ZN (n_19_39), .A (n_23_37), .B (n_29_34), .C1 (n_33_32), .C2 (n_39_29) );
AOI211_X1 g_17_40 (.ZN (n_17_40), .A (n_21_38), .B (n_27_35), .C1 (n_31_33), .C2 (n_37_30) );
AOI211_X1 g_15_41 (.ZN (n_15_41), .A (n_19_39), .B (n_25_36), .C1 (n_29_34), .C2 (n_35_31) );
AOI211_X1 g_14_43 (.ZN (n_14_43), .A (n_17_40), .B (n_23_37), .C1 (n_27_35), .C2 (n_33_32) );
AOI211_X1 g_13_41 (.ZN (n_13_41), .A (n_15_41), .B (n_21_38), .C1 (n_25_36), .C2 (n_31_33) );
AOI211_X1 g_15_40 (.ZN (n_15_40), .A (n_14_43), .B (n_19_39), .C1 (n_23_37), .C2 (n_29_34) );
AOI211_X1 g_17_39 (.ZN (n_17_39), .A (n_13_41), .B (n_17_40), .C1 (n_21_38), .C2 (n_27_35) );
AOI211_X1 g_19_38 (.ZN (n_19_38), .A (n_15_40), .B (n_15_41), .C1 (n_19_39), .C2 (n_25_36) );
AOI211_X1 g_21_37 (.ZN (n_21_37), .A (n_17_39), .B (n_14_43), .C1 (n_17_40), .C2 (n_23_37) );
AOI211_X1 g_23_36 (.ZN (n_23_36), .A (n_19_38), .B (n_13_41), .C1 (n_15_41), .C2 (n_21_38) );
AOI211_X1 g_25_35 (.ZN (n_25_35), .A (n_21_37), .B (n_15_40), .C1 (n_14_43), .C2 (n_19_39) );
AOI211_X1 g_27_36 (.ZN (n_27_36), .A (n_23_36), .B (n_17_39), .C1 (n_13_41), .C2 (n_17_40) );
AOI211_X1 g_25_37 (.ZN (n_25_37), .A (n_25_35), .B (n_19_38), .C1 (n_15_40), .C2 (n_15_41) );
AOI211_X1 g_23_38 (.ZN (n_23_38), .A (n_27_36), .B (n_21_37), .C1 (n_17_39), .C2 (n_14_43) );
AOI211_X1 g_21_39 (.ZN (n_21_39), .A (n_25_37), .B (n_23_36), .C1 (n_19_38), .C2 (n_13_41) );
AOI211_X1 g_19_40 (.ZN (n_19_40), .A (n_23_38), .B (n_25_35), .C1 (n_21_37), .C2 (n_15_40) );
AOI211_X1 g_17_41 (.ZN (n_17_41), .A (n_21_39), .B (n_27_36), .C1 (n_23_36), .C2 (n_17_39) );
AOI211_X1 g_15_42 (.ZN (n_15_42), .A (n_19_40), .B (n_25_37), .C1 (n_25_35), .C2 (n_19_38) );
AOI211_X1 g_13_43 (.ZN (n_13_43), .A (n_17_41), .B (n_23_38), .C1 (n_27_36), .C2 (n_21_37) );
AOI211_X1 g_11_44 (.ZN (n_11_44), .A (n_15_42), .B (n_21_39), .C1 (n_25_37), .C2 (n_23_36) );
AOI211_X1 g_9_45 (.ZN (n_9_45), .A (n_13_43), .B (n_19_40), .C1 (n_23_38), .C2 (n_25_35) );
AOI211_X1 g_8_47 (.ZN (n_8_47), .A (n_11_44), .B (n_17_41), .C1 (n_21_39), .C2 (n_27_36) );
AOI211_X1 g_10_46 (.ZN (n_10_46), .A (n_9_45), .B (n_15_42), .C1 (n_19_40), .C2 (n_25_37) );
AOI211_X1 g_12_45 (.ZN (n_12_45), .A (n_8_47), .B (n_13_43), .C1 (n_17_41), .C2 (n_23_38) );
AOI211_X1 g_14_44 (.ZN (n_14_44), .A (n_10_46), .B (n_11_44), .C1 (n_15_42), .C2 (n_21_39) );
AOI211_X1 g_12_43 (.ZN (n_12_43), .A (n_12_45), .B (n_9_45), .C1 (n_13_43), .C2 (n_19_40) );
AOI211_X1 g_14_42 (.ZN (n_14_42), .A (n_14_44), .B (n_8_47), .C1 (n_11_44), .C2 (n_17_41) );
AOI211_X1 g_16_41 (.ZN (n_16_41), .A (n_12_43), .B (n_10_46), .C1 (n_9_45), .C2 (n_15_42) );
AOI211_X1 g_18_40 (.ZN (n_18_40), .A (n_14_42), .B (n_12_45), .C1 (n_8_47), .C2 (n_13_43) );
AOI211_X1 g_20_39 (.ZN (n_20_39), .A (n_16_41), .B (n_14_44), .C1 (n_10_46), .C2 (n_11_44) );
AOI211_X1 g_22_38 (.ZN (n_22_38), .A (n_18_40), .B (n_12_43), .C1 (n_12_45), .C2 (n_9_45) );
AOI211_X1 g_24_37 (.ZN (n_24_37), .A (n_20_39), .B (n_14_42), .C1 (n_14_44), .C2 (n_8_47) );
AOI211_X1 g_26_36 (.ZN (n_26_36), .A (n_22_38), .B (n_16_41), .C1 (n_12_43), .C2 (n_10_46) );
AOI211_X1 g_28_35 (.ZN (n_28_35), .A (n_24_37), .B (n_18_40), .C1 (n_14_42), .C2 (n_12_45) );
AOI211_X1 g_30_34 (.ZN (n_30_34), .A (n_26_36), .B (n_20_39), .C1 (n_16_41), .C2 (n_14_44) );
AOI211_X1 g_32_33 (.ZN (n_32_33), .A (n_28_35), .B (n_22_38), .C1 (n_18_40), .C2 (n_12_43) );
AOI211_X1 g_34_32 (.ZN (n_34_32), .A (n_30_34), .B (n_24_37), .C1 (n_20_39), .C2 (n_14_42) );
AOI211_X1 g_33_34 (.ZN (n_33_34), .A (n_32_33), .B (n_26_36), .C1 (n_22_38), .C2 (n_16_41) );
AOI211_X1 g_35_33 (.ZN (n_35_33), .A (n_34_32), .B (n_28_35), .C1 (n_24_37), .C2 (n_18_40) );
AOI211_X1 g_37_32 (.ZN (n_37_32), .A (n_33_34), .B (n_30_34), .C1 (n_26_36), .C2 (n_20_39) );
AOI211_X1 g_39_31 (.ZN (n_39_31), .A (n_35_33), .B (n_32_33), .C1 (n_28_35), .C2 (n_22_38) );
AOI211_X1 g_41_30 (.ZN (n_41_30), .A (n_37_32), .B (n_34_32), .C1 (n_30_34), .C2 (n_24_37) );
AOI211_X1 g_40_32 (.ZN (n_40_32), .A (n_39_31), .B (n_33_34), .C1 (n_32_33), .C2 (n_26_36) );
AOI211_X1 g_42_31 (.ZN (n_42_31), .A (n_41_30), .B (n_35_33), .C1 (n_34_32), .C2 (n_28_35) );
AOI211_X1 g_41_29 (.ZN (n_41_29), .A (n_40_32), .B (n_37_32), .C1 (n_33_34), .C2 (n_30_34) );
AOI211_X1 g_39_30 (.ZN (n_39_30), .A (n_42_31), .B (n_39_31), .C1 (n_35_33), .C2 (n_32_33) );
AOI211_X1 g_37_31 (.ZN (n_37_31), .A (n_41_29), .B (n_41_30), .C1 (n_37_32), .C2 (n_34_32) );
AOI211_X1 g_35_32 (.ZN (n_35_32), .A (n_39_30), .B (n_40_32), .C1 (n_39_31), .C2 (n_33_34) );
AOI211_X1 g_33_33 (.ZN (n_33_33), .A (n_37_31), .B (n_42_31), .C1 (n_41_30), .C2 (n_35_33) );
AOI211_X1 g_31_34 (.ZN (n_31_34), .A (n_35_32), .B (n_41_29), .C1 (n_40_32), .C2 (n_37_32) );
AOI211_X1 g_30_36 (.ZN (n_30_36), .A (n_33_33), .B (n_39_30), .C1 (n_42_31), .C2 (n_39_31) );
AOI211_X1 g_32_35 (.ZN (n_32_35), .A (n_31_34), .B (n_37_31), .C1 (n_41_29), .C2 (n_41_30) );
AOI211_X1 g_34_34 (.ZN (n_34_34), .A (n_30_36), .B (n_35_32), .C1 (n_39_30), .C2 (n_40_32) );
AOI211_X1 g_36_33 (.ZN (n_36_33), .A (n_32_35), .B (n_33_33), .C1 (n_37_31), .C2 (n_42_31) );
AOI211_X1 g_38_32 (.ZN (n_38_32), .A (n_34_34), .B (n_31_34), .C1 (n_35_32), .C2 (n_41_29) );
AOI211_X1 g_40_31 (.ZN (n_40_31), .A (n_36_33), .B (n_30_36), .C1 (n_33_33), .C2 (n_39_30) );
AOI211_X1 g_42_30 (.ZN (n_42_30), .A (n_38_32), .B (n_32_35), .C1 (n_31_34), .C2 (n_37_31) );
AOI211_X1 g_44_29 (.ZN (n_44_29), .A (n_40_31), .B (n_34_34), .C1 (n_30_36), .C2 (n_35_32) );
AOI211_X1 g_46_28 (.ZN (n_46_28), .A (n_42_30), .B (n_36_33), .C1 (n_32_35), .C2 (n_33_33) );
AOI211_X1 g_48_27 (.ZN (n_48_27), .A (n_44_29), .B (n_38_32), .C1 (n_34_34), .C2 (n_31_34) );
AOI211_X1 g_47_29 (.ZN (n_47_29), .A (n_46_28), .B (n_40_31), .C1 (n_36_33), .C2 (n_30_36) );
AOI211_X1 g_49_28 (.ZN (n_49_28), .A (n_48_27), .B (n_42_30), .C1 (n_38_32), .C2 (n_32_35) );
AOI211_X1 g_51_27 (.ZN (n_51_27), .A (n_47_29), .B (n_44_29), .C1 (n_40_31), .C2 (n_34_34) );
AOI211_X1 g_53_26 (.ZN (n_53_26), .A (n_49_28), .B (n_46_28), .C1 (n_42_30), .C2 (n_36_33) );
AOI211_X1 g_55_25 (.ZN (n_55_25), .A (n_51_27), .B (n_48_27), .C1 (n_44_29), .C2 (n_38_32) );
AOI211_X1 g_57_24 (.ZN (n_57_24), .A (n_53_26), .B (n_47_29), .C1 (n_46_28), .C2 (n_40_31) );
AOI211_X1 g_59_23 (.ZN (n_59_23), .A (n_55_25), .B (n_49_28), .C1 (n_48_27), .C2 (n_42_30) );
AOI211_X1 g_61_22 (.ZN (n_61_22), .A (n_57_24), .B (n_51_27), .C1 (n_47_29), .C2 (n_44_29) );
AOI211_X1 g_63_21 (.ZN (n_63_21), .A (n_59_23), .B (n_53_26), .C1 (n_49_28), .C2 (n_46_28) );
AOI211_X1 g_65_20 (.ZN (n_65_20), .A (n_61_22), .B (n_55_25), .C1 (n_51_27), .C2 (n_48_27) );
AOI211_X1 g_67_19 (.ZN (n_67_19), .A (n_63_21), .B (n_57_24), .C1 (n_53_26), .C2 (n_47_29) );
AOI211_X1 g_69_18 (.ZN (n_69_18), .A (n_65_20), .B (n_59_23), .C1 (n_55_25), .C2 (n_49_28) );
AOI211_X1 g_71_17 (.ZN (n_71_17), .A (n_67_19), .B (n_61_22), .C1 (n_57_24), .C2 (n_51_27) );
AOI211_X1 g_70_19 (.ZN (n_70_19), .A (n_69_18), .B (n_63_21), .C1 (n_59_23), .C2 (n_53_26) );
AOI211_X1 g_69_17 (.ZN (n_69_17), .A (n_71_17), .B (n_65_20), .C1 (n_61_22), .C2 (n_55_25) );
AOI211_X1 g_71_16 (.ZN (n_71_16), .A (n_70_19), .B (n_67_19), .C1 (n_63_21), .C2 (n_57_24) );
AOI211_X1 g_73_15 (.ZN (n_73_15), .A (n_69_17), .B (n_69_18), .C1 (n_65_20), .C2 (n_59_23) );
AOI211_X1 g_75_14 (.ZN (n_75_14), .A (n_71_16), .B (n_71_17), .C1 (n_67_19), .C2 (n_61_22) );
AOI211_X1 g_77_13 (.ZN (n_77_13), .A (n_73_15), .B (n_70_19), .C1 (n_69_18), .C2 (n_63_21) );
AOI211_X1 g_79_12 (.ZN (n_79_12), .A (n_75_14), .B (n_69_17), .C1 (n_71_17), .C2 (n_65_20) );
AOI211_X1 g_81_11 (.ZN (n_81_11), .A (n_77_13), .B (n_71_16), .C1 (n_70_19), .C2 (n_67_19) );
AOI211_X1 g_83_10 (.ZN (n_83_10), .A (n_79_12), .B (n_73_15), .C1 (n_69_17), .C2 (n_69_18) );
AOI211_X1 g_85_9 (.ZN (n_85_9), .A (n_81_11), .B (n_75_14), .C1 (n_71_16), .C2 (n_71_17) );
AOI211_X1 g_87_8 (.ZN (n_87_8), .A (n_83_10), .B (n_77_13), .C1 (n_73_15), .C2 (n_70_19) );
AOI211_X1 g_89_7 (.ZN (n_89_7), .A (n_85_9), .B (n_79_12), .C1 (n_75_14), .C2 (n_69_17) );
AOI211_X1 g_91_6 (.ZN (n_91_6), .A (n_87_8), .B (n_81_11), .C1 (n_77_13), .C2 (n_71_16) );
AOI211_X1 g_93_5 (.ZN (n_93_5), .A (n_89_7), .B (n_83_10), .C1 (n_79_12), .C2 (n_73_15) );
AOI211_X1 g_92_7 (.ZN (n_92_7), .A (n_91_6), .B (n_85_9), .C1 (n_81_11), .C2 (n_75_14) );
AOI211_X1 g_90_8 (.ZN (n_90_8), .A (n_93_5), .B (n_87_8), .C1 (n_83_10), .C2 (n_77_13) );
AOI211_X1 g_88_9 (.ZN (n_88_9), .A (n_92_7), .B (n_89_7), .C1 (n_85_9), .C2 (n_79_12) );
AOI211_X1 g_86_10 (.ZN (n_86_10), .A (n_90_8), .B (n_91_6), .C1 (n_87_8), .C2 (n_81_11) );
AOI211_X1 g_84_11 (.ZN (n_84_11), .A (n_88_9), .B (n_93_5), .C1 (n_89_7), .C2 (n_83_10) );
AOI211_X1 g_82_12 (.ZN (n_82_12), .A (n_86_10), .B (n_92_7), .C1 (n_91_6), .C2 (n_85_9) );
AOI211_X1 g_80_13 (.ZN (n_80_13), .A (n_84_11), .B (n_90_8), .C1 (n_93_5), .C2 (n_87_8) );
AOI211_X1 g_78_14 (.ZN (n_78_14), .A (n_82_12), .B (n_88_9), .C1 (n_92_7), .C2 (n_89_7) );
AOI211_X1 g_76_15 (.ZN (n_76_15), .A (n_80_13), .B (n_86_10), .C1 (n_90_8), .C2 (n_91_6) );
AOI211_X1 g_74_16 (.ZN (n_74_16), .A (n_78_14), .B (n_84_11), .C1 (n_88_9), .C2 (n_93_5) );
AOI211_X1 g_72_17 (.ZN (n_72_17), .A (n_76_15), .B (n_82_12), .C1 (n_86_10), .C2 (n_92_7) );
AOI211_X1 g_70_18 (.ZN (n_70_18), .A (n_74_16), .B (n_80_13), .C1 (n_84_11), .C2 (n_90_8) );
AOI211_X1 g_68_19 (.ZN (n_68_19), .A (n_72_17), .B (n_78_14), .C1 (n_82_12), .C2 (n_88_9) );
AOI211_X1 g_66_20 (.ZN (n_66_20), .A (n_70_18), .B (n_76_15), .C1 (n_80_13), .C2 (n_86_10) );
AOI211_X1 g_67_18 (.ZN (n_67_18), .A (n_68_19), .B (n_74_16), .C1 (n_78_14), .C2 (n_84_11) );
AOI211_X1 g_65_19 (.ZN (n_65_19), .A (n_66_20), .B (n_72_17), .C1 (n_76_15), .C2 (n_82_12) );
AOI211_X1 g_63_20 (.ZN (n_63_20), .A (n_67_18), .B (n_70_18), .C1 (n_74_16), .C2 (n_80_13) );
AOI211_X1 g_61_21 (.ZN (n_61_21), .A (n_65_19), .B (n_68_19), .C1 (n_72_17), .C2 (n_78_14) );
AOI211_X1 g_59_22 (.ZN (n_59_22), .A (n_63_20), .B (n_66_20), .C1 (n_70_18), .C2 (n_76_15) );
AOI211_X1 g_57_23 (.ZN (n_57_23), .A (n_61_21), .B (n_67_18), .C1 (n_68_19), .C2 (n_74_16) );
AOI211_X1 g_55_24 (.ZN (n_55_24), .A (n_59_22), .B (n_65_19), .C1 (n_66_20), .C2 (n_72_17) );
AOI211_X1 g_53_25 (.ZN (n_53_25), .A (n_57_23), .B (n_63_20), .C1 (n_67_18), .C2 (n_70_18) );
AOI211_X1 g_51_26 (.ZN (n_51_26), .A (n_55_24), .B (n_61_21), .C1 (n_65_19), .C2 (n_68_19) );
AOI211_X1 g_49_27 (.ZN (n_49_27), .A (n_53_25), .B (n_59_22), .C1 (n_63_20), .C2 (n_66_20) );
AOI211_X1 g_47_28 (.ZN (n_47_28), .A (n_51_26), .B (n_57_23), .C1 (n_61_21), .C2 (n_67_18) );
AOI211_X1 g_45_29 (.ZN (n_45_29), .A (n_49_27), .B (n_55_24), .C1 (n_59_22), .C2 (n_65_19) );
AOI211_X1 g_43_30 (.ZN (n_43_30), .A (n_47_28), .B (n_53_25), .C1 (n_57_23), .C2 (n_63_20) );
AOI211_X1 g_41_31 (.ZN (n_41_31), .A (n_45_29), .B (n_51_26), .C1 (n_55_24), .C2 (n_61_21) );
AOI211_X1 g_39_32 (.ZN (n_39_32), .A (n_43_30), .B (n_49_27), .C1 (n_53_25), .C2 (n_59_22) );
AOI211_X1 g_37_33 (.ZN (n_37_33), .A (n_41_31), .B (n_47_28), .C1 (n_51_26), .C2 (n_57_23) );
AOI211_X1 g_35_34 (.ZN (n_35_34), .A (n_39_32), .B (n_45_29), .C1 (n_49_27), .C2 (n_55_24) );
AOI211_X1 g_36_32 (.ZN (n_36_32), .A (n_37_33), .B (n_43_30), .C1 (n_47_28), .C2 (n_53_25) );
AOI211_X1 g_34_33 (.ZN (n_34_33), .A (n_35_34), .B (n_41_31), .C1 (n_45_29), .C2 (n_51_26) );
AOI211_X1 g_32_34 (.ZN (n_32_34), .A (n_36_32), .B (n_39_32), .C1 (n_43_30), .C2 (n_49_27) );
AOI211_X1 g_30_35 (.ZN (n_30_35), .A (n_34_33), .B (n_37_33), .C1 (n_41_31), .C2 (n_47_28) );
AOI211_X1 g_28_36 (.ZN (n_28_36), .A (n_32_34), .B (n_35_34), .C1 (n_39_32), .C2 (n_45_29) );
AOI211_X1 g_26_37 (.ZN (n_26_37), .A (n_30_35), .B (n_36_32), .C1 (n_37_33), .C2 (n_43_30) );
AOI211_X1 g_24_38 (.ZN (n_24_38), .A (n_28_36), .B (n_34_33), .C1 (n_35_34), .C2 (n_41_31) );
AOI211_X1 g_22_39 (.ZN (n_22_39), .A (n_26_37), .B (n_32_34), .C1 (n_36_32), .C2 (n_39_32) );
AOI211_X1 g_20_40 (.ZN (n_20_40), .A (n_24_38), .B (n_30_35), .C1 (n_34_33), .C2 (n_37_33) );
AOI211_X1 g_18_41 (.ZN (n_18_41), .A (n_22_39), .B (n_28_36), .C1 (n_32_34), .C2 (n_35_34) );
AOI211_X1 g_16_42 (.ZN (n_16_42), .A (n_20_40), .B (n_26_37), .C1 (n_30_35), .C2 (n_36_32) );
AOI211_X1 g_15_44 (.ZN (n_15_44), .A (n_18_41), .B (n_24_38), .C1 (n_28_36), .C2 (n_34_33) );
AOI211_X1 g_17_43 (.ZN (n_17_43), .A (n_16_42), .B (n_22_39), .C1 (n_26_37), .C2 (n_32_34) );
AOI211_X1 g_19_42 (.ZN (n_19_42), .A (n_15_44), .B (n_20_40), .C1 (n_24_38), .C2 (n_30_35) );
AOI211_X1 g_21_41 (.ZN (n_21_41), .A (n_17_43), .B (n_18_41), .C1 (n_22_39), .C2 (n_28_36) );
AOI211_X1 g_23_40 (.ZN (n_23_40), .A (n_19_42), .B (n_16_42), .C1 (n_20_40), .C2 (n_26_37) );
AOI211_X1 g_25_39 (.ZN (n_25_39), .A (n_21_41), .B (n_15_44), .C1 (n_18_41), .C2 (n_24_38) );
AOI211_X1 g_27_38 (.ZN (n_27_38), .A (n_23_40), .B (n_17_43), .C1 (n_16_42), .C2 (n_22_39) );
AOI211_X1 g_29_37 (.ZN (n_29_37), .A (n_25_39), .B (n_19_42), .C1 (n_15_44), .C2 (n_20_40) );
AOI211_X1 g_31_36 (.ZN (n_31_36), .A (n_27_38), .B (n_21_41), .C1 (n_17_43), .C2 (n_18_41) );
AOI211_X1 g_33_35 (.ZN (n_33_35), .A (n_29_37), .B (n_23_40), .C1 (n_19_42), .C2 (n_16_42) );
AOI211_X1 g_32_37 (.ZN (n_32_37), .A (n_31_36), .B (n_25_39), .C1 (n_21_41), .C2 (n_15_44) );
AOI211_X1 g_31_35 (.ZN (n_31_35), .A (n_33_35), .B (n_27_38), .C1 (n_23_40), .C2 (n_17_43) );
AOI211_X1 g_29_36 (.ZN (n_29_36), .A (n_32_37), .B (n_29_37), .C1 (n_25_39), .C2 (n_19_42) );
AOI211_X1 g_27_37 (.ZN (n_27_37), .A (n_31_35), .B (n_31_36), .C1 (n_27_38), .C2 (n_21_41) );
AOI211_X1 g_25_38 (.ZN (n_25_38), .A (n_29_36), .B (n_33_35), .C1 (n_29_37), .C2 (n_23_40) );
AOI211_X1 g_23_39 (.ZN (n_23_39), .A (n_27_37), .B (n_32_37), .C1 (n_31_36), .C2 (n_25_39) );
AOI211_X1 g_21_40 (.ZN (n_21_40), .A (n_25_38), .B (n_31_35), .C1 (n_33_35), .C2 (n_27_38) );
AOI211_X1 g_19_41 (.ZN (n_19_41), .A (n_23_39), .B (n_29_36), .C1 (n_32_37), .C2 (n_29_37) );
AOI211_X1 g_17_42 (.ZN (n_17_42), .A (n_21_40), .B (n_27_37), .C1 (n_31_35), .C2 (n_31_36) );
AOI211_X1 g_15_43 (.ZN (n_15_43), .A (n_19_41), .B (n_25_38), .C1 (n_29_36), .C2 (n_33_35) );
AOI211_X1 g_13_44 (.ZN (n_13_44), .A (n_17_42), .B (n_23_39), .C1 (n_27_37), .C2 (n_32_37) );
AOI211_X1 g_11_45 (.ZN (n_11_45), .A (n_15_43), .B (n_21_40), .C1 (n_25_38), .C2 (n_31_35) );
AOI211_X1 g_10_47 (.ZN (n_10_47), .A (n_13_44), .B (n_19_41), .C1 (n_23_39), .C2 (n_29_36) );
AOI211_X1 g_8_46 (.ZN (n_8_46), .A (n_11_45), .B (n_17_42), .C1 (n_21_40), .C2 (n_27_37) );
AOI211_X1 g_10_45 (.ZN (n_10_45), .A (n_10_47), .B (n_15_43), .C1 (n_19_41), .C2 (n_25_38) );
AOI211_X1 g_12_44 (.ZN (n_12_44), .A (n_8_46), .B (n_13_44), .C1 (n_17_42), .C2 (n_23_39) );
AOI211_X1 g_11_46 (.ZN (n_11_46), .A (n_10_45), .B (n_11_45), .C1 (n_15_43), .C2 (n_21_40) );
AOI211_X1 g_13_45 (.ZN (n_13_45), .A (n_12_44), .B (n_10_47), .C1 (n_13_44), .C2 (n_19_41) );
AOI211_X1 g_12_47 (.ZN (n_12_47), .A (n_11_46), .B (n_8_46), .C1 (n_11_45), .C2 (n_17_42) );
AOI211_X1 g_14_46 (.ZN (n_14_46), .A (n_13_45), .B (n_10_45), .C1 (n_10_47), .C2 (n_15_43) );
AOI211_X1 g_16_45 (.ZN (n_16_45), .A (n_12_47), .B (n_12_44), .C1 (n_8_46), .C2 (n_13_44) );
AOI211_X1 g_18_44 (.ZN (n_18_44), .A (n_14_46), .B (n_11_46), .C1 (n_10_45), .C2 (n_11_45) );
AOI211_X1 g_16_43 (.ZN (n_16_43), .A (n_16_45), .B (n_13_45), .C1 (n_12_44), .C2 (n_10_47) );
AOI211_X1 g_18_42 (.ZN (n_18_42), .A (n_18_44), .B (n_12_47), .C1 (n_11_46), .C2 (n_8_46) );
AOI211_X1 g_20_41 (.ZN (n_20_41), .A (n_16_43), .B (n_14_46), .C1 (n_13_45), .C2 (n_10_45) );
AOI211_X1 g_22_40 (.ZN (n_22_40), .A (n_18_42), .B (n_16_45), .C1 (n_12_47), .C2 (n_12_44) );
AOI211_X1 g_24_39 (.ZN (n_24_39), .A (n_20_41), .B (n_18_44), .C1 (n_14_46), .C2 (n_11_46) );
AOI211_X1 g_26_38 (.ZN (n_26_38), .A (n_22_40), .B (n_16_43), .C1 (n_16_45), .C2 (n_13_45) );
AOI211_X1 g_28_37 (.ZN (n_28_37), .A (n_24_39), .B (n_18_42), .C1 (n_18_44), .C2 (n_12_47) );
AOI211_X1 g_30_38 (.ZN (n_30_38), .A (n_26_38), .B (n_20_41), .C1 (n_16_43), .C2 (n_14_46) );
AOI211_X1 g_28_39 (.ZN (n_28_39), .A (n_28_37), .B (n_22_40), .C1 (n_18_42), .C2 (n_16_45) );
AOI211_X1 g_26_40 (.ZN (n_26_40), .A (n_30_38), .B (n_24_39), .C1 (n_20_41), .C2 (n_18_44) );
AOI211_X1 g_24_41 (.ZN (n_24_41), .A (n_28_39), .B (n_26_38), .C1 (n_22_40), .C2 (n_16_43) );
AOI211_X1 g_22_42 (.ZN (n_22_42), .A (n_26_40), .B (n_28_37), .C1 (n_24_39), .C2 (n_18_42) );
AOI211_X1 g_20_43 (.ZN (n_20_43), .A (n_24_41), .B (n_30_38), .C1 (n_26_38), .C2 (n_20_41) );
AOI211_X1 g_19_45 (.ZN (n_19_45), .A (n_22_42), .B (n_28_39), .C1 (n_28_37), .C2 (n_22_40) );
AOI211_X1 g_18_43 (.ZN (n_18_43), .A (n_20_43), .B (n_26_40), .C1 (n_30_38), .C2 (n_24_39) );
AOI211_X1 g_20_42 (.ZN (n_20_42), .A (n_19_45), .B (n_24_41), .C1 (n_28_39), .C2 (n_26_38) );
AOI211_X1 g_22_41 (.ZN (n_22_41), .A (n_18_43), .B (n_22_42), .C1 (n_26_40), .C2 (n_28_37) );
AOI211_X1 g_24_40 (.ZN (n_24_40), .A (n_20_42), .B (n_20_43), .C1 (n_24_41), .C2 (n_30_38) );
AOI211_X1 g_26_39 (.ZN (n_26_39), .A (n_22_41), .B (n_19_45), .C1 (n_22_42), .C2 (n_28_39) );
AOI211_X1 g_28_38 (.ZN (n_28_38), .A (n_24_40), .B (n_18_43), .C1 (n_20_43), .C2 (n_26_40) );
AOI211_X1 g_30_37 (.ZN (n_30_37), .A (n_26_39), .B (n_20_42), .C1 (n_19_45), .C2 (n_24_41) );
AOI211_X1 g_32_36 (.ZN (n_32_36), .A (n_28_38), .B (n_22_41), .C1 (n_18_43), .C2 (n_22_42) );
AOI211_X1 g_34_35 (.ZN (n_34_35), .A (n_30_37), .B (n_24_40), .C1 (n_20_42), .C2 (n_20_43) );
AOI211_X1 g_36_34 (.ZN (n_36_34), .A (n_32_36), .B (n_26_39), .C1 (n_22_41), .C2 (n_19_45) );
AOI211_X1 g_38_33 (.ZN (n_38_33), .A (n_34_35), .B (n_28_38), .C1 (n_24_40), .C2 (n_18_43) );
AOI211_X1 g_37_35 (.ZN (n_37_35), .A (n_36_34), .B (n_30_37), .C1 (n_26_39), .C2 (n_20_42) );
AOI211_X1 g_39_34 (.ZN (n_39_34), .A (n_38_33), .B (n_32_36), .C1 (n_28_38), .C2 (n_22_41) );
AOI211_X1 g_41_33 (.ZN (n_41_33), .A (n_37_35), .B (n_34_35), .C1 (n_30_37), .C2 (n_24_40) );
AOI211_X1 g_43_32 (.ZN (n_43_32), .A (n_39_34), .B (n_36_34), .C1 (n_32_36), .C2 (n_26_39) );
AOI211_X1 g_45_31 (.ZN (n_45_31), .A (n_41_33), .B (n_38_33), .C1 (n_34_35), .C2 (n_28_38) );
AOI211_X1 g_46_29 (.ZN (n_46_29), .A (n_43_32), .B (n_37_35), .C1 (n_36_34), .C2 (n_30_37) );
AOI211_X1 g_48_28 (.ZN (n_48_28), .A (n_45_31), .B (n_39_34), .C1 (n_38_33), .C2 (n_32_36) );
AOI211_X1 g_50_27 (.ZN (n_50_27), .A (n_46_29), .B (n_41_33), .C1 (n_37_35), .C2 (n_34_35) );
AOI211_X1 g_52_26 (.ZN (n_52_26), .A (n_48_28), .B (n_43_32), .C1 (n_39_34), .C2 (n_36_34) );
AOI211_X1 g_54_25 (.ZN (n_54_25), .A (n_50_27), .B (n_45_31), .C1 (n_41_33), .C2 (n_38_33) );
AOI211_X1 g_56_24 (.ZN (n_56_24), .A (n_52_26), .B (n_46_29), .C1 (n_43_32), .C2 (n_37_35) );
AOI211_X1 g_58_23 (.ZN (n_58_23), .A (n_54_25), .B (n_48_28), .C1 (n_45_31), .C2 (n_39_34) );
AOI211_X1 g_60_22 (.ZN (n_60_22), .A (n_56_24), .B (n_50_27), .C1 (n_46_29), .C2 (n_41_33) );
AOI211_X1 g_62_21 (.ZN (n_62_21), .A (n_58_23), .B (n_52_26), .C1 (n_48_28), .C2 (n_43_32) );
AOI211_X1 g_64_20 (.ZN (n_64_20), .A (n_60_22), .B (n_54_25), .C1 (n_50_27), .C2 (n_45_31) );
AOI211_X1 g_66_19 (.ZN (n_66_19), .A (n_62_21), .B (n_56_24), .C1 (n_52_26), .C2 (n_46_29) );
AOI211_X1 g_68_18 (.ZN (n_68_18), .A (n_64_20), .B (n_58_23), .C1 (n_54_25), .C2 (n_48_28) );
AOI211_X1 g_70_17 (.ZN (n_70_17), .A (n_66_19), .B (n_60_22), .C1 (n_56_24), .C2 (n_50_27) );
AOI211_X1 g_72_16 (.ZN (n_72_16), .A (n_68_18), .B (n_62_21), .C1 (n_58_23), .C2 (n_52_26) );
AOI211_X1 g_74_15 (.ZN (n_74_15), .A (n_70_17), .B (n_64_20), .C1 (n_60_22), .C2 (n_54_25) );
AOI211_X1 g_76_14 (.ZN (n_76_14), .A (n_72_16), .B (n_66_19), .C1 (n_62_21), .C2 (n_56_24) );
AOI211_X1 g_78_13 (.ZN (n_78_13), .A (n_74_15), .B (n_68_18), .C1 (n_64_20), .C2 (n_58_23) );
AOI211_X1 g_77_15 (.ZN (n_77_15), .A (n_76_14), .B (n_70_17), .C1 (n_66_19), .C2 (n_60_22) );
AOI211_X1 g_79_14 (.ZN (n_79_14), .A (n_78_13), .B (n_72_16), .C1 (n_68_18), .C2 (n_62_21) );
AOI211_X1 g_81_13 (.ZN (n_81_13), .A (n_77_15), .B (n_74_15), .C1 (n_70_17), .C2 (n_64_20) );
AOI211_X1 g_83_12 (.ZN (n_83_12), .A (n_79_14), .B (n_76_14), .C1 (n_72_16), .C2 (n_66_19) );
AOI211_X1 g_85_11 (.ZN (n_85_11), .A (n_81_13), .B (n_78_13), .C1 (n_74_15), .C2 (n_68_18) );
AOI211_X1 g_87_10 (.ZN (n_87_10), .A (n_83_12), .B (n_77_15), .C1 (n_76_14), .C2 (n_70_17) );
AOI211_X1 g_88_8 (.ZN (n_88_8), .A (n_85_11), .B (n_79_14), .C1 (n_78_13), .C2 (n_72_16) );
AOI211_X1 g_90_7 (.ZN (n_90_7), .A (n_87_10), .B (n_81_13), .C1 (n_77_15), .C2 (n_74_15) );
AOI211_X1 g_89_9 (.ZN (n_89_9), .A (n_88_8), .B (n_83_12), .C1 (n_79_14), .C2 (n_76_14) );
AOI211_X1 g_91_8 (.ZN (n_91_8), .A (n_90_7), .B (n_85_11), .C1 (n_81_13), .C2 (n_78_13) );
AOI211_X1 g_93_7 (.ZN (n_93_7), .A (n_89_9), .B (n_87_10), .C1 (n_83_12), .C2 (n_77_15) );
AOI211_X1 g_94_5 (.ZN (n_94_5), .A (n_91_8), .B (n_88_8), .C1 (n_85_11), .C2 (n_79_14) );
AOI211_X1 g_96_4 (.ZN (n_96_4), .A (n_93_7), .B (n_90_7), .C1 (n_87_10), .C2 (n_81_13) );
AOI211_X1 g_98_3 (.ZN (n_98_3), .A (n_94_5), .B (n_89_9), .C1 (n_88_8), .C2 (n_83_12) );
AOI211_X1 g_100_4 (.ZN (n_100_4), .A (n_96_4), .B (n_91_8), .C1 (n_90_7), .C2 (n_85_11) );
AOI211_X1 g_98_5 (.ZN (n_98_5), .A (n_98_3), .B (n_93_7), .C1 (n_89_9), .C2 (n_87_10) );
AOI211_X1 g_96_6 (.ZN (n_96_6), .A (n_100_4), .B (n_94_5), .C1 (n_91_8), .C2 (n_88_8) );
AOI211_X1 g_94_7 (.ZN (n_94_7), .A (n_98_5), .B (n_96_4), .C1 (n_93_7), .C2 (n_90_7) );
AOI211_X1 g_92_8 (.ZN (n_92_8), .A (n_96_6), .B (n_98_3), .C1 (n_94_5), .C2 (n_89_9) );
AOI211_X1 g_90_9 (.ZN (n_90_9), .A (n_94_7), .B (n_100_4), .C1 (n_96_4), .C2 (n_91_8) );
AOI211_X1 g_88_10 (.ZN (n_88_10), .A (n_92_8), .B (n_98_5), .C1 (n_98_3), .C2 (n_93_7) );
AOI211_X1 g_86_11 (.ZN (n_86_11), .A (n_90_9), .B (n_96_6), .C1 (n_100_4), .C2 (n_94_5) );
AOI211_X1 g_84_12 (.ZN (n_84_12), .A (n_88_10), .B (n_94_7), .C1 (n_98_5), .C2 (n_96_4) );
AOI211_X1 g_82_13 (.ZN (n_82_13), .A (n_86_11), .B (n_92_8), .C1 (n_96_6), .C2 (n_98_3) );
AOI211_X1 g_80_14 (.ZN (n_80_14), .A (n_84_12), .B (n_90_9), .C1 (n_94_7), .C2 (n_100_4) );
AOI211_X1 g_78_15 (.ZN (n_78_15), .A (n_82_13), .B (n_88_10), .C1 (n_92_8), .C2 (n_98_5) );
AOI211_X1 g_76_16 (.ZN (n_76_16), .A (n_80_14), .B (n_86_11), .C1 (n_90_9), .C2 (n_96_6) );
AOI211_X1 g_74_17 (.ZN (n_74_17), .A (n_78_15), .B (n_84_12), .C1 (n_88_10), .C2 (n_94_7) );
AOI211_X1 g_72_18 (.ZN (n_72_18), .A (n_76_16), .B (n_82_13), .C1 (n_86_11), .C2 (n_92_8) );
AOI211_X1 g_71_20 (.ZN (n_71_20), .A (n_74_17), .B (n_80_14), .C1 (n_84_12), .C2 (n_90_9) );
AOI211_X1 g_69_19 (.ZN (n_69_19), .A (n_72_18), .B (n_78_15), .C1 (n_82_13), .C2 (n_88_10) );
AOI211_X1 g_71_18 (.ZN (n_71_18), .A (n_71_20), .B (n_76_16), .C1 (n_80_14), .C2 (n_86_11) );
AOI211_X1 g_73_17 (.ZN (n_73_17), .A (n_69_19), .B (n_74_17), .C1 (n_78_15), .C2 (n_84_12) );
AOI211_X1 g_75_16 (.ZN (n_75_16), .A (n_71_18), .B (n_72_18), .C1 (n_76_16), .C2 (n_82_13) );
AOI211_X1 g_74_18 (.ZN (n_74_18), .A (n_73_17), .B (n_71_20), .C1 (n_74_17), .C2 (n_80_14) );
AOI211_X1 g_76_17 (.ZN (n_76_17), .A (n_75_16), .B (n_69_19), .C1 (n_72_18), .C2 (n_78_15) );
AOI211_X1 g_78_16 (.ZN (n_78_16), .A (n_74_18), .B (n_71_18), .C1 (n_71_20), .C2 (n_76_16) );
AOI211_X1 g_80_15 (.ZN (n_80_15), .A (n_76_17), .B (n_73_17), .C1 (n_69_19), .C2 (n_74_17) );
AOI211_X1 g_82_14 (.ZN (n_82_14), .A (n_78_16), .B (n_75_16), .C1 (n_71_18), .C2 (n_72_18) );
AOI211_X1 g_84_13 (.ZN (n_84_13), .A (n_80_15), .B (n_74_18), .C1 (n_73_17), .C2 (n_71_20) );
AOI211_X1 g_86_12 (.ZN (n_86_12), .A (n_82_14), .B (n_76_17), .C1 (n_75_16), .C2 (n_69_19) );
AOI211_X1 g_88_11 (.ZN (n_88_11), .A (n_84_13), .B (n_78_16), .C1 (n_74_18), .C2 (n_71_18) );
AOI211_X1 g_90_10 (.ZN (n_90_10), .A (n_86_12), .B (n_80_15), .C1 (n_76_17), .C2 (n_73_17) );
AOI211_X1 g_92_9 (.ZN (n_92_9), .A (n_88_11), .B (n_82_14), .C1 (n_78_16), .C2 (n_75_16) );
AOI211_X1 g_94_8 (.ZN (n_94_8), .A (n_90_10), .B (n_84_13), .C1 (n_80_15), .C2 (n_74_18) );
AOI211_X1 g_95_6 (.ZN (n_95_6), .A (n_92_9), .B (n_86_12), .C1 (n_82_14), .C2 (n_76_17) );
AOI211_X1 g_97_5 (.ZN (n_97_5), .A (n_94_8), .B (n_88_11), .C1 (n_84_13), .C2 (n_78_16) );
AOI211_X1 g_96_7 (.ZN (n_96_7), .A (n_95_6), .B (n_90_10), .C1 (n_86_12), .C2 (n_80_15) );
AOI211_X1 g_95_9 (.ZN (n_95_9), .A (n_97_5), .B (n_92_9), .C1 (n_88_11), .C2 (n_82_14) );
AOI211_X1 g_93_8 (.ZN (n_93_8), .A (n_96_7), .B (n_94_8), .C1 (n_90_10), .C2 (n_84_13) );
AOI211_X1 g_95_7 (.ZN (n_95_7), .A (n_95_9), .B (n_95_6), .C1 (n_92_9), .C2 (n_86_12) );
AOI211_X1 g_97_6 (.ZN (n_97_6), .A (n_93_8), .B (n_97_5), .C1 (n_94_8), .C2 (n_88_11) );
AOI211_X1 g_99_7 (.ZN (n_99_7), .A (n_95_7), .B (n_96_7), .C1 (n_95_6), .C2 (n_90_10) );
AOI211_X1 g_97_8 (.ZN (n_97_8), .A (n_97_6), .B (n_95_9), .C1 (n_97_5), .C2 (n_92_9) );
AOI211_X1 g_99_9 (.ZN (n_99_9), .A (n_99_7), .B (n_93_8), .C1 (n_96_7), .C2 (n_94_8) );
AOI211_X1 g_98_7 (.ZN (n_98_7), .A (n_97_8), .B (n_95_7), .C1 (n_95_9), .C2 (n_95_6) );
AOI211_X1 g_100_8 (.ZN (n_100_8), .A (n_99_9), .B (n_97_6), .C1 (n_93_8), .C2 (n_97_5) );
AOI211_X1 g_99_6 (.ZN (n_99_6), .A (n_98_7), .B (n_99_7), .C1 (n_95_7), .C2 (n_96_7) );
AOI211_X1 g_97_7 (.ZN (n_97_7), .A (n_100_8), .B (n_97_8), .C1 (n_97_6), .C2 (n_95_9) );
AOI211_X1 g_95_8 (.ZN (n_95_8), .A (n_99_6), .B (n_99_9), .C1 (n_99_7), .C2 (n_93_8) );
AOI211_X1 g_93_9 (.ZN (n_93_9), .A (n_97_7), .B (n_98_7), .C1 (n_97_8), .C2 (n_95_7) );
AOI211_X1 g_91_10 (.ZN (n_91_10), .A (n_95_8), .B (n_100_8), .C1 (n_99_9), .C2 (n_97_6) );
AOI211_X1 g_89_11 (.ZN (n_89_11), .A (n_93_9), .B (n_99_6), .C1 (n_98_7), .C2 (n_99_7) );
AOI211_X1 g_87_12 (.ZN (n_87_12), .A (n_91_10), .B (n_97_7), .C1 (n_100_8), .C2 (n_97_8) );
AOI211_X1 g_85_13 (.ZN (n_85_13), .A (n_89_11), .B (n_95_8), .C1 (n_99_6), .C2 (n_99_9) );
AOI211_X1 g_83_14 (.ZN (n_83_14), .A (n_87_12), .B (n_93_9), .C1 (n_97_7), .C2 (n_98_7) );
AOI211_X1 g_81_15 (.ZN (n_81_15), .A (n_85_13), .B (n_91_10), .C1 (n_95_8), .C2 (n_100_8) );
AOI211_X1 g_79_16 (.ZN (n_79_16), .A (n_83_14), .B (n_89_11), .C1 (n_93_9), .C2 (n_99_6) );
AOI211_X1 g_77_17 (.ZN (n_77_17), .A (n_81_15), .B (n_87_12), .C1 (n_91_10), .C2 (n_97_7) );
AOI211_X1 g_75_18 (.ZN (n_75_18), .A (n_79_16), .B (n_85_13), .C1 (n_89_11), .C2 (n_95_8) );
AOI211_X1 g_73_19 (.ZN (n_73_19), .A (n_77_17), .B (n_83_14), .C1 (n_87_12), .C2 (n_93_9) );
AOI211_X1 g_75_20 (.ZN (n_75_20), .A (n_75_18), .B (n_81_15), .C1 (n_85_13), .C2 (n_91_10) );
AOI211_X1 g_77_19 (.ZN (n_77_19), .A (n_73_19), .B (n_79_16), .C1 (n_83_14), .C2 (n_89_11) );
AOI211_X1 g_79_18 (.ZN (n_79_18), .A (n_75_20), .B (n_77_17), .C1 (n_81_15), .C2 (n_87_12) );
AOI211_X1 g_81_17 (.ZN (n_81_17), .A (n_77_19), .B (n_75_18), .C1 (n_79_16), .C2 (n_85_13) );
AOI211_X1 g_83_16 (.ZN (n_83_16), .A (n_79_18), .B (n_73_19), .C1 (n_77_17), .C2 (n_83_14) );
AOI211_X1 g_85_15 (.ZN (n_85_15), .A (n_81_17), .B (n_75_20), .C1 (n_75_18), .C2 (n_81_15) );
AOI211_X1 g_87_14 (.ZN (n_87_14), .A (n_83_16), .B (n_77_19), .C1 (n_73_19), .C2 (n_79_16) );
AOI211_X1 g_89_13 (.ZN (n_89_13), .A (n_85_15), .B (n_79_18), .C1 (n_75_20), .C2 (n_77_17) );
AOI211_X1 g_91_12 (.ZN (n_91_12), .A (n_87_14), .B (n_81_17), .C1 (n_77_19), .C2 (n_75_18) );
AOI211_X1 g_92_10 (.ZN (n_92_10), .A (n_89_13), .B (n_83_16), .C1 (n_79_18), .C2 (n_73_19) );
AOI211_X1 g_94_9 (.ZN (n_94_9), .A (n_91_12), .B (n_85_15), .C1 (n_81_17), .C2 (n_75_20) );
AOI211_X1 g_96_8 (.ZN (n_96_8), .A (n_92_10), .B (n_87_14), .C1 (n_83_16), .C2 (n_77_19) );
AOI211_X1 g_98_9 (.ZN (n_98_9), .A (n_94_9), .B (n_89_13), .C1 (n_85_15), .C2 (n_79_18) );
AOI211_X1 g_96_10 (.ZN (n_96_10), .A (n_96_8), .B (n_91_12), .C1 (n_87_14), .C2 (n_81_17) );
AOI211_X1 g_94_11 (.ZN (n_94_11), .A (n_98_9), .B (n_92_10), .C1 (n_89_13), .C2 (n_83_16) );
AOI211_X1 g_92_12 (.ZN (n_92_12), .A (n_96_10), .B (n_94_9), .C1 (n_91_12), .C2 (n_85_15) );
AOI211_X1 g_90_11 (.ZN (n_90_11), .A (n_94_11), .B (n_96_8), .C1 (n_92_10), .C2 (n_87_14) );
AOI211_X1 g_91_9 (.ZN (n_91_9), .A (n_92_12), .B (n_98_9), .C1 (n_94_9), .C2 (n_89_13) );
AOI211_X1 g_93_10 (.ZN (n_93_10), .A (n_90_11), .B (n_96_10), .C1 (n_96_8), .C2 (n_91_12) );
AOI211_X1 g_91_11 (.ZN (n_91_11), .A (n_91_9), .B (n_94_11), .C1 (n_98_9), .C2 (n_92_10) );
AOI211_X1 g_89_10 (.ZN (n_89_10), .A (n_93_10), .B (n_92_12), .C1 (n_96_10), .C2 (n_94_9) );
AOI211_X1 g_88_12 (.ZN (n_88_12), .A (n_91_11), .B (n_90_11), .C1 (n_94_11), .C2 (n_96_8) );
AOI211_X1 g_86_13 (.ZN (n_86_13), .A (n_89_10), .B (n_91_9), .C1 (n_92_12), .C2 (n_98_9) );
AOI211_X1 g_87_11 (.ZN (n_87_11), .A (n_88_12), .B (n_93_10), .C1 (n_90_11), .C2 (n_96_10) );
AOI211_X1 g_85_12 (.ZN (n_85_12), .A (n_86_13), .B (n_91_11), .C1 (n_91_9), .C2 (n_94_11) );
AOI211_X1 g_84_14 (.ZN (n_84_14), .A (n_87_11), .B (n_89_10), .C1 (n_93_10), .C2 (n_92_12) );
AOI211_X1 g_82_15 (.ZN (n_82_15), .A (n_85_12), .B (n_88_12), .C1 (n_91_11), .C2 (n_90_11) );
AOI211_X1 g_83_13 (.ZN (n_83_13), .A (n_84_14), .B (n_86_13), .C1 (n_89_10), .C2 (n_91_9) );
AOI211_X1 g_81_14 (.ZN (n_81_14), .A (n_82_15), .B (n_87_11), .C1 (n_88_12), .C2 (n_93_10) );
AOI211_X1 g_80_16 (.ZN (n_80_16), .A (n_83_13), .B (n_85_12), .C1 (n_86_13), .C2 (n_91_11) );
AOI211_X1 g_78_17 (.ZN (n_78_17), .A (n_81_14), .B (n_84_14), .C1 (n_87_11), .C2 (n_89_10) );
AOI211_X1 g_79_15 (.ZN (n_79_15), .A (n_80_16), .B (n_82_15), .C1 (n_85_12), .C2 (n_88_12) );
AOI211_X1 g_77_16 (.ZN (n_77_16), .A (n_78_17), .B (n_83_13), .C1 (n_84_14), .C2 (n_86_13) );
AOI211_X1 g_76_18 (.ZN (n_76_18), .A (n_79_15), .B (n_81_14), .C1 (n_82_15), .C2 (n_87_11) );
AOI211_X1 g_74_19 (.ZN (n_74_19), .A (n_77_16), .B (n_80_16), .C1 (n_83_13), .C2 (n_85_12) );
AOI211_X1 g_75_17 (.ZN (n_75_17), .A (n_76_18), .B (n_78_17), .C1 (n_81_14), .C2 (n_84_14) );
AOI211_X1 g_73_18 (.ZN (n_73_18), .A (n_74_19), .B (n_79_15), .C1 (n_80_16), .C2 (n_82_15) );
AOI211_X1 g_71_19 (.ZN (n_71_19), .A (n_75_17), .B (n_77_16), .C1 (n_78_17), .C2 (n_83_13) );
AOI211_X1 g_69_20 (.ZN (n_69_20), .A (n_73_18), .B (n_76_18), .C1 (n_79_15), .C2 (n_81_14) );
AOI211_X1 g_67_21 (.ZN (n_67_21), .A (n_71_19), .B (n_74_19), .C1 (n_77_16), .C2 (n_80_16) );
AOI211_X1 g_65_22 (.ZN (n_65_22), .A (n_69_20), .B (n_75_17), .C1 (n_76_18), .C2 (n_78_17) );
AOI211_X1 g_63_23 (.ZN (n_63_23), .A (n_67_21), .B (n_73_18), .C1 (n_74_19), .C2 (n_79_15) );
AOI211_X1 g_64_21 (.ZN (n_64_21), .A (n_65_22), .B (n_71_19), .C1 (n_75_17), .C2 (n_77_16) );
AOI211_X1 g_62_22 (.ZN (n_62_22), .A (n_63_23), .B (n_69_20), .C1 (n_73_18), .C2 (n_76_18) );
AOI211_X1 g_60_23 (.ZN (n_60_23), .A (n_64_21), .B (n_67_21), .C1 (n_71_19), .C2 (n_74_19) );
AOI211_X1 g_58_24 (.ZN (n_58_24), .A (n_62_22), .B (n_65_22), .C1 (n_69_20), .C2 (n_75_17) );
AOI211_X1 g_56_25 (.ZN (n_56_25), .A (n_60_23), .B (n_63_23), .C1 (n_67_21), .C2 (n_73_18) );
AOI211_X1 g_54_26 (.ZN (n_54_26), .A (n_58_24), .B (n_64_21), .C1 (n_65_22), .C2 (n_71_19) );
AOI211_X1 g_52_27 (.ZN (n_52_27), .A (n_56_25), .B (n_62_22), .C1 (n_63_23), .C2 (n_69_20) );
AOI211_X1 g_50_28 (.ZN (n_50_28), .A (n_54_26), .B (n_60_23), .C1 (n_64_21), .C2 (n_67_21) );
AOI211_X1 g_48_29 (.ZN (n_48_29), .A (n_52_27), .B (n_58_24), .C1 (n_62_22), .C2 (n_65_22) );
AOI211_X1 g_46_30 (.ZN (n_46_30), .A (n_50_28), .B (n_56_25), .C1 (n_60_23), .C2 (n_63_23) );
AOI211_X1 g_44_31 (.ZN (n_44_31), .A (n_48_29), .B (n_54_26), .C1 (n_58_24), .C2 (n_64_21) );
AOI211_X1 g_42_32 (.ZN (n_42_32), .A (n_46_30), .B (n_52_27), .C1 (n_56_25), .C2 (n_62_22) );
AOI211_X1 g_40_33 (.ZN (n_40_33), .A (n_44_31), .B (n_50_28), .C1 (n_54_26), .C2 (n_60_23) );
AOI211_X1 g_38_34 (.ZN (n_38_34), .A (n_42_32), .B (n_48_29), .C1 (n_52_27), .C2 (n_58_24) );
AOI211_X1 g_36_35 (.ZN (n_36_35), .A (n_40_33), .B (n_46_30), .C1 (n_50_28), .C2 (n_56_25) );
AOI211_X1 g_34_36 (.ZN (n_34_36), .A (n_38_34), .B (n_44_31), .C1 (n_48_29), .C2 (n_54_26) );
AOI211_X1 g_33_38 (.ZN (n_33_38), .A (n_36_35), .B (n_42_32), .C1 (n_46_30), .C2 (n_52_27) );
AOI211_X1 g_31_37 (.ZN (n_31_37), .A (n_34_36), .B (n_40_33), .C1 (n_44_31), .C2 (n_50_28) );
AOI211_X1 g_33_36 (.ZN (n_33_36), .A (n_33_38), .B (n_38_34), .C1 (n_42_32), .C2 (n_48_29) );
AOI211_X1 g_35_35 (.ZN (n_35_35), .A (n_31_37), .B (n_36_35), .C1 (n_40_33), .C2 (n_46_30) );
AOI211_X1 g_37_34 (.ZN (n_37_34), .A (n_33_36), .B (n_34_36), .C1 (n_38_34), .C2 (n_44_31) );
AOI211_X1 g_39_33 (.ZN (n_39_33), .A (n_35_35), .B (n_33_38), .C1 (n_36_35), .C2 (n_42_32) );
AOI211_X1 g_41_32 (.ZN (n_41_32), .A (n_37_34), .B (n_31_37), .C1 (n_34_36), .C2 (n_40_33) );
AOI211_X1 g_43_31 (.ZN (n_43_31), .A (n_39_33), .B (n_33_36), .C1 (n_33_38), .C2 (n_38_34) );
AOI211_X1 g_45_30 (.ZN (n_45_30), .A (n_41_32), .B (n_35_35), .C1 (n_31_37), .C2 (n_36_35) );
AOI211_X1 g_44_32 (.ZN (n_44_32), .A (n_43_31), .B (n_37_34), .C1 (n_33_36), .C2 (n_34_36) );
AOI211_X1 g_46_31 (.ZN (n_46_31), .A (n_45_30), .B (n_39_33), .C1 (n_35_35), .C2 (n_33_38) );
AOI211_X1 g_48_30 (.ZN (n_48_30), .A (n_44_32), .B (n_41_32), .C1 (n_37_34), .C2 (n_31_37) );
AOI211_X1 g_50_29 (.ZN (n_50_29), .A (n_46_31), .B (n_43_31), .C1 (n_39_33), .C2 (n_33_36) );
AOI211_X1 g_52_28 (.ZN (n_52_28), .A (n_48_30), .B (n_45_30), .C1 (n_41_32), .C2 (n_35_35) );
AOI211_X1 g_54_27 (.ZN (n_54_27), .A (n_50_29), .B (n_44_32), .C1 (n_43_31), .C2 (n_37_34) );
AOI211_X1 g_56_26 (.ZN (n_56_26), .A (n_52_28), .B (n_46_31), .C1 (n_45_30), .C2 (n_39_33) );
AOI211_X1 g_58_25 (.ZN (n_58_25), .A (n_54_27), .B (n_48_30), .C1 (n_44_32), .C2 (n_41_32) );
AOI211_X1 g_60_24 (.ZN (n_60_24), .A (n_56_26), .B (n_50_29), .C1 (n_46_31), .C2 (n_43_31) );
AOI211_X1 g_62_23 (.ZN (n_62_23), .A (n_58_25), .B (n_52_28), .C1 (n_48_30), .C2 (n_45_30) );
AOI211_X1 g_64_22 (.ZN (n_64_22), .A (n_60_24), .B (n_54_27), .C1 (n_50_29), .C2 (n_44_32) );
AOI211_X1 g_66_21 (.ZN (n_66_21), .A (n_62_23), .B (n_56_26), .C1 (n_52_28), .C2 (n_46_31) );
AOI211_X1 g_68_20 (.ZN (n_68_20), .A (n_64_22), .B (n_58_25), .C1 (n_54_27), .C2 (n_48_30) );
AOI211_X1 g_70_21 (.ZN (n_70_21), .A (n_66_21), .B (n_60_24), .C1 (n_56_26), .C2 (n_50_29) );
AOI211_X1 g_72_20 (.ZN (n_72_20), .A (n_68_20), .B (n_62_23), .C1 (n_58_25), .C2 (n_52_28) );
AOI211_X1 g_74_21 (.ZN (n_74_21), .A (n_70_21), .B (n_64_22), .C1 (n_60_24), .C2 (n_54_27) );
AOI211_X1 g_75_19 (.ZN (n_75_19), .A (n_72_20), .B (n_66_21), .C1 (n_62_23), .C2 (n_56_26) );
AOI211_X1 g_77_18 (.ZN (n_77_18), .A (n_74_21), .B (n_68_20), .C1 (n_64_22), .C2 (n_58_25) );
AOI211_X1 g_79_17 (.ZN (n_79_17), .A (n_75_19), .B (n_70_21), .C1 (n_66_21), .C2 (n_60_24) );
AOI211_X1 g_81_16 (.ZN (n_81_16), .A (n_77_18), .B (n_72_20), .C1 (n_68_20), .C2 (n_62_23) );
AOI211_X1 g_83_15 (.ZN (n_83_15), .A (n_79_17), .B (n_74_21), .C1 (n_70_21), .C2 (n_64_22) );
AOI211_X1 g_85_14 (.ZN (n_85_14), .A (n_81_16), .B (n_75_19), .C1 (n_72_20), .C2 (n_66_21) );
AOI211_X1 g_87_13 (.ZN (n_87_13), .A (n_83_15), .B (n_77_18), .C1 (n_74_21), .C2 (n_68_20) );
AOI211_X1 g_89_12 (.ZN (n_89_12), .A (n_85_14), .B (n_79_17), .C1 (n_75_19), .C2 (n_70_21) );
AOI211_X1 g_88_14 (.ZN (n_88_14), .A (n_87_13), .B (n_81_16), .C1 (n_77_18), .C2 (n_72_20) );
AOI211_X1 g_90_13 (.ZN (n_90_13), .A (n_89_12), .B (n_83_15), .C1 (n_79_17), .C2 (n_74_21) );
AOI211_X1 g_89_15 (.ZN (n_89_15), .A (n_88_14), .B (n_85_14), .C1 (n_81_16), .C2 (n_75_19) );
AOI211_X1 g_88_13 (.ZN (n_88_13), .A (n_90_13), .B (n_87_13), .C1 (n_83_15), .C2 (n_77_18) );
AOI211_X1 g_90_12 (.ZN (n_90_12), .A (n_89_15), .B (n_89_12), .C1 (n_85_14), .C2 (n_79_17) );
AOI211_X1 g_92_11 (.ZN (n_92_11), .A (n_88_13), .B (n_88_14), .C1 (n_87_13), .C2 (n_81_16) );
AOI211_X1 g_94_10 (.ZN (n_94_10), .A (n_90_12), .B (n_90_13), .C1 (n_89_12), .C2 (n_83_15) );
AOI211_X1 g_96_9 (.ZN (n_96_9), .A (n_92_11), .B (n_89_15), .C1 (n_88_14), .C2 (n_85_14) );
AOI211_X1 g_98_8 (.ZN (n_98_8), .A (n_94_10), .B (n_88_13), .C1 (n_90_13), .C2 (n_87_13) );
AOI211_X1 g_100_9 (.ZN (n_100_9), .A (n_96_9), .B (n_90_12), .C1 (n_89_15), .C2 (n_89_12) );
AOI211_X1 g_98_10 (.ZN (n_98_10), .A (n_98_8), .B (n_92_11), .C1 (n_88_13), .C2 (n_88_14) );
AOI211_X1 g_100_11 (.ZN (n_100_11), .A (n_100_9), .B (n_94_10), .C1 (n_90_12), .C2 (n_90_13) );
AOI211_X1 g_99_13 (.ZN (n_99_13), .A (n_98_10), .B (n_96_9), .C1 (n_92_11), .C2 (n_89_15) );
AOI211_X1 g_100_15 (.ZN (n_100_15), .A (n_100_11), .B (n_98_8), .C1 (n_94_10), .C2 (n_88_13) );
AOI211_X1 g_98_14 (.ZN (n_98_14), .A (n_99_13), .B (n_100_9), .C1 (n_96_9), .C2 (n_90_12) );
AOI211_X1 g_100_13 (.ZN (n_100_13), .A (n_100_15), .B (n_98_10), .C1 (n_98_8), .C2 (n_92_11) );
AOI211_X1 g_99_11 (.ZN (n_99_11), .A (n_98_14), .B (n_100_11), .C1 (n_100_9), .C2 (n_94_10) );
AOI211_X1 g_97_10 (.ZN (n_97_10), .A (n_100_13), .B (n_99_13), .C1 (n_98_10), .C2 (n_96_9) );
AOI211_X1 g_95_11 (.ZN (n_95_11), .A (n_99_11), .B (n_100_15), .C1 (n_100_11), .C2 (n_98_8) );
AOI211_X1 g_97_12 (.ZN (n_97_12), .A (n_97_10), .B (n_98_14), .C1 (n_99_13), .C2 (n_100_9) );
AOI211_X1 g_95_13 (.ZN (n_95_13), .A (n_95_11), .B (n_100_13), .C1 (n_100_15), .C2 (n_98_10) );
AOI211_X1 g_93_12 (.ZN (n_93_12), .A (n_97_12), .B (n_99_11), .C1 (n_98_14), .C2 (n_100_11) );
AOI211_X1 g_91_13 (.ZN (n_91_13), .A (n_95_13), .B (n_97_10), .C1 (n_100_13), .C2 (n_99_13) );
AOI211_X1 g_89_14 (.ZN (n_89_14), .A (n_93_12), .B (n_95_11), .C1 (n_99_11), .C2 (n_100_15) );
AOI211_X1 g_87_15 (.ZN (n_87_15), .A (n_91_13), .B (n_97_12), .C1 (n_97_10), .C2 (n_98_14) );
AOI211_X1 g_85_16 (.ZN (n_85_16), .A (n_89_14), .B (n_95_13), .C1 (n_95_11), .C2 (n_100_13) );
AOI211_X1 g_86_14 (.ZN (n_86_14), .A (n_87_15), .B (n_93_12), .C1 (n_97_12), .C2 (n_99_11) );
AOI211_X1 g_84_15 (.ZN (n_84_15), .A (n_85_16), .B (n_91_13), .C1 (n_95_13), .C2 (n_97_10) );
AOI211_X1 g_82_16 (.ZN (n_82_16), .A (n_86_14), .B (n_89_14), .C1 (n_93_12), .C2 (n_95_11) );
AOI211_X1 g_80_17 (.ZN (n_80_17), .A (n_84_15), .B (n_87_15), .C1 (n_91_13), .C2 (n_97_12) );
AOI211_X1 g_78_18 (.ZN (n_78_18), .A (n_82_16), .B (n_85_16), .C1 (n_89_14), .C2 (n_95_13) );
AOI211_X1 g_76_19 (.ZN (n_76_19), .A (n_80_17), .B (n_86_14), .C1 (n_87_15), .C2 (n_93_12) );
AOI211_X1 g_74_20 (.ZN (n_74_20), .A (n_78_18), .B (n_84_15), .C1 (n_85_16), .C2 (n_91_13) );
AOI211_X1 g_72_19 (.ZN (n_72_19), .A (n_76_19), .B (n_82_16), .C1 (n_86_14), .C2 (n_89_14) );
AOI211_X1 g_70_20 (.ZN (n_70_20), .A (n_74_20), .B (n_80_17), .C1 (n_84_15), .C2 (n_87_15) );
AOI211_X1 g_68_21 (.ZN (n_68_21), .A (n_72_19), .B (n_78_18), .C1 (n_82_16), .C2 (n_85_16) );
AOI211_X1 g_66_22 (.ZN (n_66_22), .A (n_70_20), .B (n_76_19), .C1 (n_80_17), .C2 (n_86_14) );
AOI211_X1 g_67_20 (.ZN (n_67_20), .A (n_68_21), .B (n_74_20), .C1 (n_78_18), .C2 (n_84_15) );
AOI211_X1 g_65_21 (.ZN (n_65_21), .A (n_66_22), .B (n_72_19), .C1 (n_76_19), .C2 (n_82_16) );
AOI211_X1 g_63_22 (.ZN (n_63_22), .A (n_67_20), .B (n_70_20), .C1 (n_74_20), .C2 (n_80_17) );
AOI211_X1 g_61_23 (.ZN (n_61_23), .A (n_65_21), .B (n_68_21), .C1 (n_72_19), .C2 (n_78_18) );
AOI211_X1 g_59_24 (.ZN (n_59_24), .A (n_63_22), .B (n_66_22), .C1 (n_70_20), .C2 (n_76_19) );
AOI211_X1 g_57_25 (.ZN (n_57_25), .A (n_61_23), .B (n_67_20), .C1 (n_68_21), .C2 (n_74_20) );
AOI211_X1 g_55_26 (.ZN (n_55_26), .A (n_59_24), .B (n_65_21), .C1 (n_66_22), .C2 (n_72_19) );
AOI211_X1 g_53_27 (.ZN (n_53_27), .A (n_57_25), .B (n_63_22), .C1 (n_67_20), .C2 (n_70_20) );
AOI211_X1 g_51_28 (.ZN (n_51_28), .A (n_55_26), .B (n_61_23), .C1 (n_65_21), .C2 (n_68_21) );
AOI211_X1 g_49_29 (.ZN (n_49_29), .A (n_53_27), .B (n_59_24), .C1 (n_63_22), .C2 (n_66_22) );
AOI211_X1 g_47_30 (.ZN (n_47_30), .A (n_51_28), .B (n_57_25), .C1 (n_61_23), .C2 (n_67_20) );
AOI211_X1 g_46_32 (.ZN (n_46_32), .A (n_49_29), .B (n_55_26), .C1 (n_59_24), .C2 (n_65_21) );
AOI211_X1 g_48_31 (.ZN (n_48_31), .A (n_47_30), .B (n_53_27), .C1 (n_57_25), .C2 (n_63_22) );
AOI211_X1 g_50_30 (.ZN (n_50_30), .A (n_46_32), .B (n_51_28), .C1 (n_55_26), .C2 (n_61_23) );
AOI211_X1 g_52_29 (.ZN (n_52_29), .A (n_48_31), .B (n_49_29), .C1 (n_53_27), .C2 (n_59_24) );
AOI211_X1 g_54_28 (.ZN (n_54_28), .A (n_50_30), .B (n_47_30), .C1 (n_51_28), .C2 (n_57_25) );
AOI211_X1 g_56_27 (.ZN (n_56_27), .A (n_52_29), .B (n_46_32), .C1 (n_49_29), .C2 (n_55_26) );
AOI211_X1 g_58_26 (.ZN (n_58_26), .A (n_54_28), .B (n_48_31), .C1 (n_47_30), .C2 (n_53_27) );
AOI211_X1 g_60_25 (.ZN (n_60_25), .A (n_56_27), .B (n_50_30), .C1 (n_46_32), .C2 (n_51_28) );
AOI211_X1 g_62_24 (.ZN (n_62_24), .A (n_58_26), .B (n_52_29), .C1 (n_48_31), .C2 (n_49_29) );
AOI211_X1 g_64_23 (.ZN (n_64_23), .A (n_60_25), .B (n_54_28), .C1 (n_50_30), .C2 (n_47_30) );
AOI211_X1 g_63_25 (.ZN (n_63_25), .A (n_62_24), .B (n_56_27), .C1 (n_52_29), .C2 (n_46_32) );
AOI211_X1 g_61_24 (.ZN (n_61_24), .A (n_64_23), .B (n_58_26), .C1 (n_54_28), .C2 (n_48_31) );
AOI211_X1 g_59_25 (.ZN (n_59_25), .A (n_63_25), .B (n_60_25), .C1 (n_56_27), .C2 (n_50_30) );
AOI211_X1 g_57_26 (.ZN (n_57_26), .A (n_61_24), .B (n_62_24), .C1 (n_58_26), .C2 (n_52_29) );
AOI211_X1 g_55_27 (.ZN (n_55_27), .A (n_59_25), .B (n_64_23), .C1 (n_60_25), .C2 (n_54_28) );
AOI211_X1 g_53_28 (.ZN (n_53_28), .A (n_57_26), .B (n_63_25), .C1 (n_62_24), .C2 (n_56_27) );
AOI211_X1 g_51_29 (.ZN (n_51_29), .A (n_55_27), .B (n_61_24), .C1 (n_64_23), .C2 (n_58_26) );
AOI211_X1 g_49_30 (.ZN (n_49_30), .A (n_53_28), .B (n_59_25), .C1 (n_63_25), .C2 (n_60_25) );
AOI211_X1 g_47_31 (.ZN (n_47_31), .A (n_51_29), .B (n_57_26), .C1 (n_61_24), .C2 (n_62_24) );
AOI211_X1 g_45_32 (.ZN (n_45_32), .A (n_49_30), .B (n_55_27), .C1 (n_59_25), .C2 (n_64_23) );
AOI211_X1 g_43_33 (.ZN (n_43_33), .A (n_47_31), .B (n_53_28), .C1 (n_57_26), .C2 (n_63_25) );
AOI211_X1 g_41_34 (.ZN (n_41_34), .A (n_45_32), .B (n_51_29), .C1 (n_55_27), .C2 (n_61_24) );
AOI211_X1 g_39_35 (.ZN (n_39_35), .A (n_43_33), .B (n_49_30), .C1 (n_53_28), .C2 (n_59_25) );
AOI211_X1 g_37_36 (.ZN (n_37_36), .A (n_41_34), .B (n_47_31), .C1 (n_51_29), .C2 (n_57_26) );
AOI211_X1 g_35_37 (.ZN (n_35_37), .A (n_39_35), .B (n_45_32), .C1 (n_49_30), .C2 (n_55_27) );
AOI211_X1 g_34_39 (.ZN (n_34_39), .A (n_37_36), .B (n_43_33), .C1 (n_47_31), .C2 (n_53_28) );
AOI211_X1 g_33_37 (.ZN (n_33_37), .A (n_35_37), .B (n_41_34), .C1 (n_45_32), .C2 (n_51_29) );
AOI211_X1 g_35_36 (.ZN (n_35_36), .A (n_34_39), .B (n_39_35), .C1 (n_43_33), .C2 (n_49_30) );
AOI211_X1 g_34_38 (.ZN (n_34_38), .A (n_33_37), .B (n_37_36), .C1 (n_41_34), .C2 (n_47_31) );
AOI211_X1 g_36_37 (.ZN (n_36_37), .A (n_35_36), .B (n_35_37), .C1 (n_39_35), .C2 (n_45_32) );
AOI211_X1 g_38_36 (.ZN (n_38_36), .A (n_34_38), .B (n_34_39), .C1 (n_37_36), .C2 (n_43_33) );
AOI211_X1 g_40_35 (.ZN (n_40_35), .A (n_36_37), .B (n_33_37), .C1 (n_35_37), .C2 (n_41_34) );
AOI211_X1 g_42_34 (.ZN (n_42_34), .A (n_38_36), .B (n_35_36), .C1 (n_34_39), .C2 (n_39_35) );
AOI211_X1 g_44_33 (.ZN (n_44_33), .A (n_40_35), .B (n_34_38), .C1 (n_33_37), .C2 (n_37_36) );
AOI211_X1 g_43_35 (.ZN (n_43_35), .A (n_42_34), .B (n_36_37), .C1 (n_35_36), .C2 (n_35_37) );
AOI211_X1 g_42_33 (.ZN (n_42_33), .A (n_44_33), .B (n_38_36), .C1 (n_34_38), .C2 (n_34_39) );
AOI211_X1 g_40_34 (.ZN (n_40_34), .A (n_43_35), .B (n_40_35), .C1 (n_36_37), .C2 (n_33_37) );
AOI211_X1 g_38_35 (.ZN (n_38_35), .A (n_42_33), .B (n_42_34), .C1 (n_38_36), .C2 (n_35_36) );
AOI211_X1 g_36_36 (.ZN (n_36_36), .A (n_40_34), .B (n_44_33), .C1 (n_40_35), .C2 (n_34_38) );
AOI211_X1 g_34_37 (.ZN (n_34_37), .A (n_38_35), .B (n_43_35), .C1 (n_42_34), .C2 (n_36_37) );
AOI211_X1 g_32_38 (.ZN (n_32_38), .A (n_36_36), .B (n_42_33), .C1 (n_44_33), .C2 (n_38_36) );
AOI211_X1 g_30_39 (.ZN (n_30_39), .A (n_34_37), .B (n_40_34), .C1 (n_43_35), .C2 (n_40_35) );
AOI211_X1 g_28_40 (.ZN (n_28_40), .A (n_32_38), .B (n_38_35), .C1 (n_42_33), .C2 (n_42_34) );
AOI211_X1 g_29_38 (.ZN (n_29_38), .A (n_30_39), .B (n_36_36), .C1 (n_40_34), .C2 (n_44_33) );
AOI211_X1 g_27_39 (.ZN (n_27_39), .A (n_28_40), .B (n_34_37), .C1 (n_38_35), .C2 (n_43_35) );
AOI211_X1 g_25_40 (.ZN (n_25_40), .A (n_29_38), .B (n_32_38), .C1 (n_36_36), .C2 (n_42_33) );
AOI211_X1 g_23_41 (.ZN (n_23_41), .A (n_27_39), .B (n_30_39), .C1 (n_34_37), .C2 (n_40_34) );
AOI211_X1 g_21_42 (.ZN (n_21_42), .A (n_25_40), .B (n_28_40), .C1 (n_32_38), .C2 (n_38_35) );
AOI211_X1 g_19_43 (.ZN (n_19_43), .A (n_23_41), .B (n_29_38), .C1 (n_30_39), .C2 (n_36_36) );
AOI211_X1 g_17_44 (.ZN (n_17_44), .A (n_21_42), .B (n_27_39), .C1 (n_28_40), .C2 (n_34_37) );
AOI211_X1 g_15_45 (.ZN (n_15_45), .A (n_19_43), .B (n_25_40), .C1 (n_29_38), .C2 (n_32_38) );
AOI211_X1 g_13_46 (.ZN (n_13_46), .A (n_17_44), .B (n_23_41), .C1 (n_27_39), .C2 (n_30_39) );
AOI211_X1 g_11_47 (.ZN (n_11_47), .A (n_15_45), .B (n_21_42), .C1 (n_25_40), .C2 (n_28_40) );
AOI211_X1 g_9_48 (.ZN (n_9_48), .A (n_13_46), .B (n_19_43), .C1 (n_23_41), .C2 (n_29_38) );
AOI211_X1 g_7_49 (.ZN (n_7_49), .A (n_11_47), .B (n_17_44), .C1 (n_21_42), .C2 (n_27_39) );
AOI211_X1 g_6_51 (.ZN (n_6_51), .A (n_9_48), .B (n_15_45), .C1 (n_19_43), .C2 (n_25_40) );
AOI211_X1 g_5_53 (.ZN (n_5_53), .A (n_7_49), .B (n_13_46), .C1 (n_17_44), .C2 (n_23_41) );
AOI211_X1 g_4_55 (.ZN (n_4_55), .A (n_6_51), .B (n_11_47), .C1 (n_15_45), .C2 (n_21_42) );
AOI211_X1 g_6_56 (.ZN (n_6_56), .A (n_5_53), .B (n_9_48), .C1 (n_13_46), .C2 (n_19_43) );
AOI211_X1 g_4_57 (.ZN (n_4_57), .A (n_4_55), .B (n_7_49), .C1 (n_11_47), .C2 (n_17_44) );
AOI211_X1 g_2_58 (.ZN (n_2_58), .A (n_6_56), .B (n_6_51), .C1 (n_9_48), .C2 (n_15_45) );
AOI211_X1 g_3_56 (.ZN (n_3_56), .A (n_4_57), .B (n_5_53), .C1 (n_7_49), .C2 (n_13_46) );
AOI211_X1 g_5_55 (.ZN (n_5_55), .A (n_2_58), .B (n_4_55), .C1 (n_6_51), .C2 (n_11_47) );
AOI211_X1 g_7_54 (.ZN (n_7_54), .A (n_3_56), .B (n_6_56), .C1 (n_5_53), .C2 (n_9_48) );
AOI211_X1 g_8_52 (.ZN (n_8_52), .A (n_5_55), .B (n_4_57), .C1 (n_4_55), .C2 (n_7_49) );
AOI211_X1 g_6_53 (.ZN (n_6_53), .A (n_7_54), .B (n_2_58), .C1 (n_6_56), .C2 (n_6_51) );
AOI211_X1 g_4_54 (.ZN (n_4_54), .A (n_8_52), .B (n_3_56), .C1 (n_4_57), .C2 (n_5_53) );
AOI211_X1 g_5_52 (.ZN (n_5_52), .A (n_6_53), .B (n_5_55), .C1 (n_2_58), .C2 (n_4_55) );
AOI211_X1 g_7_51 (.ZN (n_7_51), .A (n_4_54), .B (n_7_54), .C1 (n_3_56), .C2 (n_6_56) );
AOI211_X1 g_9_50 (.ZN (n_9_50), .A (n_5_52), .B (n_8_52), .C1 (n_5_55), .C2 (n_4_57) );
AOI211_X1 g_10_48 (.ZN (n_10_48), .A (n_7_51), .B (n_6_53), .C1 (n_7_54), .C2 (n_2_58) );
AOI211_X1 g_8_49 (.ZN (n_8_49), .A (n_9_50), .B (n_4_54), .C1 (n_8_52), .C2 (n_3_56) );
AOI211_X1 g_9_47 (.ZN (n_9_47), .A (n_10_48), .B (n_5_52), .C1 (n_6_53), .C2 (n_5_55) );
AOI211_X1 g_7_48 (.ZN (n_7_48), .A (n_8_49), .B (n_7_51), .C1 (n_4_54), .C2 (n_7_54) );
AOI211_X1 g_6_50 (.ZN (n_6_50), .A (n_9_47), .B (n_9_50), .C1 (n_5_52), .C2 (n_8_52) );
AOI211_X1 g_7_52 (.ZN (n_7_52), .A (n_7_48), .B (n_10_48), .C1 (n_7_51), .C2 (n_6_53) );
AOI211_X1 g_8_50 (.ZN (n_8_50), .A (n_6_50), .B (n_8_49), .C1 (n_9_50), .C2 (n_4_54) );
AOI211_X1 g_10_49 (.ZN (n_10_49), .A (n_7_52), .B (n_9_47), .C1 (n_10_48), .C2 (n_5_52) );
AOI211_X1 g_12_48 (.ZN (n_12_48), .A (n_8_50), .B (n_7_48), .C1 (n_8_49), .C2 (n_7_51) );
AOI211_X1 g_14_47 (.ZN (n_14_47), .A (n_10_49), .B (n_6_50), .C1 (n_9_47), .C2 (n_9_50) );
AOI211_X1 g_12_46 (.ZN (n_12_46), .A (n_12_48), .B (n_7_52), .C1 (n_7_48), .C2 (n_10_48) );
AOI211_X1 g_14_45 (.ZN (n_14_45), .A (n_14_47), .B (n_8_50), .C1 (n_6_50), .C2 (n_8_49) );
AOI211_X1 g_16_44 (.ZN (n_16_44), .A (n_12_46), .B (n_10_49), .C1 (n_7_52), .C2 (n_9_47) );
AOI211_X1 g_17_46 (.ZN (n_17_46), .A (n_14_45), .B (n_12_48), .C1 (n_8_50), .C2 (n_7_48) );
AOI211_X1 g_15_47 (.ZN (n_15_47), .A (n_16_44), .B (n_14_47), .C1 (n_10_49), .C2 (n_6_50) );
AOI211_X1 g_13_48 (.ZN (n_13_48), .A (n_17_46), .B (n_12_46), .C1 (n_12_48), .C2 (n_7_52) );
AOI211_X1 g_11_49 (.ZN (n_11_49), .A (n_15_47), .B (n_14_45), .C1 (n_14_47), .C2 (n_8_50) );
AOI211_X1 g_10_51 (.ZN (n_10_51), .A (n_13_48), .B (n_16_44), .C1 (n_12_46), .C2 (n_10_49) );
AOI211_X1 g_9_49 (.ZN (n_9_49), .A (n_11_49), .B (n_17_46), .C1 (n_14_45), .C2 (n_12_48) );
AOI211_X1 g_11_48 (.ZN (n_11_48), .A (n_10_51), .B (n_15_47), .C1 (n_16_44), .C2 (n_14_47) );
AOI211_X1 g_13_47 (.ZN (n_13_47), .A (n_9_49), .B (n_13_48), .C1 (n_17_46), .C2 (n_12_46) );
AOI211_X1 g_15_46 (.ZN (n_15_46), .A (n_11_48), .B (n_11_49), .C1 (n_15_47), .C2 (n_14_45) );
AOI211_X1 g_17_45 (.ZN (n_17_45), .A (n_13_47), .B (n_10_51), .C1 (n_13_48), .C2 (n_16_44) );
AOI211_X1 g_19_44 (.ZN (n_19_44), .A (n_15_46), .B (n_9_49), .C1 (n_11_49), .C2 (n_17_46) );
AOI211_X1 g_21_43 (.ZN (n_21_43), .A (n_17_45), .B (n_11_48), .C1 (n_10_51), .C2 (n_15_47) );
AOI211_X1 g_23_42 (.ZN (n_23_42), .A (n_19_44), .B (n_13_47), .C1 (n_9_49), .C2 (n_13_48) );
AOI211_X1 g_25_41 (.ZN (n_25_41), .A (n_21_43), .B (n_15_46), .C1 (n_11_48), .C2 (n_11_49) );
AOI211_X1 g_27_40 (.ZN (n_27_40), .A (n_23_42), .B (n_17_45), .C1 (n_13_47), .C2 (n_10_51) );
AOI211_X1 g_29_39 (.ZN (n_29_39), .A (n_25_41), .B (n_19_44), .C1 (n_15_46), .C2 (n_9_49) );
AOI211_X1 g_31_38 (.ZN (n_31_38), .A (n_27_40), .B (n_21_43), .C1 (n_17_45), .C2 (n_11_48) );
AOI211_X1 g_32_40 (.ZN (n_32_40), .A (n_29_39), .B (n_23_42), .C1 (n_19_44), .C2 (n_13_47) );
AOI211_X1 g_30_41 (.ZN (n_30_41), .A (n_31_38), .B (n_25_41), .C1 (n_21_43), .C2 (n_15_46) );
AOI211_X1 g_31_39 (.ZN (n_31_39), .A (n_32_40), .B (n_27_40), .C1 (n_23_42), .C2 (n_17_45) );
AOI211_X1 g_29_40 (.ZN (n_29_40), .A (n_30_41), .B (n_29_39), .C1 (n_25_41), .C2 (n_19_44) );
AOI211_X1 g_27_41 (.ZN (n_27_41), .A (n_31_39), .B (n_31_38), .C1 (n_27_40), .C2 (n_21_43) );
AOI211_X1 g_25_42 (.ZN (n_25_42), .A (n_29_40), .B (n_32_40), .C1 (n_29_39), .C2 (n_23_42) );
AOI211_X1 g_23_43 (.ZN (n_23_43), .A (n_27_41), .B (n_30_41), .C1 (n_31_38), .C2 (n_25_41) );
AOI211_X1 g_21_44 (.ZN (n_21_44), .A (n_25_42), .B (n_31_39), .C1 (n_32_40), .C2 (n_27_40) );
AOI211_X1 g_20_46 (.ZN (n_20_46), .A (n_23_43), .B (n_29_40), .C1 (n_30_41), .C2 (n_29_39) );
AOI211_X1 g_18_45 (.ZN (n_18_45), .A (n_21_44), .B (n_27_41), .C1 (n_31_39), .C2 (n_31_38) );
AOI211_X1 g_16_46 (.ZN (n_16_46), .A (n_20_46), .B (n_25_42), .C1 (n_29_40), .C2 (n_32_40) );
AOI211_X1 g_18_47 (.ZN (n_18_47), .A (n_18_45), .B (n_23_43), .C1 (n_27_41), .C2 (n_30_41) );
AOI211_X1 g_16_48 (.ZN (n_16_48), .A (n_16_46), .B (n_21_44), .C1 (n_25_42), .C2 (n_31_39) );
AOI211_X1 g_14_49 (.ZN (n_14_49), .A (n_18_47), .B (n_20_46), .C1 (n_23_43), .C2 (n_29_40) );
AOI211_X1 g_12_50 (.ZN (n_12_50), .A (n_16_48), .B (n_18_45), .C1 (n_21_44), .C2 (n_27_41) );
AOI211_X1 g_11_52 (.ZN (n_11_52), .A (n_14_49), .B (n_16_46), .C1 (n_20_46), .C2 (n_25_42) );
AOI211_X1 g_9_51 (.ZN (n_9_51), .A (n_12_50), .B (n_18_47), .C1 (n_18_45), .C2 (n_23_43) );
AOI211_X1 g_11_50 (.ZN (n_11_50), .A (n_11_52), .B (n_16_48), .C1 (n_16_46), .C2 (n_21_44) );
AOI211_X1 g_13_49 (.ZN (n_13_49), .A (n_9_51), .B (n_14_49), .C1 (n_18_47), .C2 (n_20_46) );
AOI211_X1 g_15_48 (.ZN (n_15_48), .A (n_11_50), .B (n_12_50), .C1 (n_16_48), .C2 (n_18_45) );
AOI211_X1 g_17_47 (.ZN (n_17_47), .A (n_13_49), .B (n_11_52), .C1 (n_14_49), .C2 (n_16_46) );
AOI211_X1 g_19_46 (.ZN (n_19_46), .A (n_15_48), .B (n_9_51), .C1 (n_12_50), .C2 (n_18_47) );
AOI211_X1 g_20_44 (.ZN (n_20_44), .A (n_17_47), .B (n_11_50), .C1 (n_11_52), .C2 (n_16_48) );
AOI211_X1 g_22_43 (.ZN (n_22_43), .A (n_19_46), .B (n_13_49), .C1 (n_9_51), .C2 (n_14_49) );
AOI211_X1 g_24_42 (.ZN (n_24_42), .A (n_20_44), .B (n_15_48), .C1 (n_11_50), .C2 (n_12_50) );
AOI211_X1 g_26_41 (.ZN (n_26_41), .A (n_22_43), .B (n_17_47), .C1 (n_13_49), .C2 (n_11_52) );
AOI211_X1 g_28_42 (.ZN (n_28_42), .A (n_24_42), .B (n_19_46), .C1 (n_15_48), .C2 (n_9_51) );
AOI211_X1 g_26_43 (.ZN (n_26_43), .A (n_26_41), .B (n_20_44), .C1 (n_17_47), .C2 (n_11_50) );
AOI211_X1 g_24_44 (.ZN (n_24_44), .A (n_28_42), .B (n_22_43), .C1 (n_19_46), .C2 (n_13_49) );
AOI211_X1 g_22_45 (.ZN (n_22_45), .A (n_26_43), .B (n_24_42), .C1 (n_20_44), .C2 (n_15_48) );
AOI211_X1 g_21_47 (.ZN (n_21_47), .A (n_24_44), .B (n_26_41), .C1 (n_22_43), .C2 (n_17_47) );
AOI211_X1 g_20_45 (.ZN (n_20_45), .A (n_22_45), .B (n_28_42), .C1 (n_24_42), .C2 (n_19_46) );
AOI211_X1 g_22_44 (.ZN (n_22_44), .A (n_21_47), .B (n_26_43), .C1 (n_26_41), .C2 (n_20_44) );
AOI211_X1 g_24_43 (.ZN (n_24_43), .A (n_20_45), .B (n_24_44), .C1 (n_28_42), .C2 (n_22_43) );
AOI211_X1 g_26_42 (.ZN (n_26_42), .A (n_22_44), .B (n_22_45), .C1 (n_26_43), .C2 (n_24_42) );
AOI211_X1 g_28_41 (.ZN (n_28_41), .A (n_24_43), .B (n_21_47), .C1 (n_24_44), .C2 (n_26_41) );
AOI211_X1 g_30_40 (.ZN (n_30_40), .A (n_26_42), .B (n_20_45), .C1 (n_22_45), .C2 (n_28_42) );
AOI211_X1 g_32_39 (.ZN (n_32_39), .A (n_28_41), .B (n_22_44), .C1 (n_21_47), .C2 (n_26_43) );
AOI211_X1 g_31_41 (.ZN (n_31_41), .A (n_30_40), .B (n_24_43), .C1 (n_20_45), .C2 (n_24_44) );
AOI211_X1 g_33_40 (.ZN (n_33_40), .A (n_32_39), .B (n_26_42), .C1 (n_22_44), .C2 (n_22_45) );
AOI211_X1 g_35_39 (.ZN (n_35_39), .A (n_31_41), .B (n_28_41), .C1 (n_24_43), .C2 (n_21_47) );
AOI211_X1 g_37_38 (.ZN (n_37_38), .A (n_33_40), .B (n_30_40), .C1 (n_26_42), .C2 (n_20_45) );
AOI211_X1 g_39_37 (.ZN (n_39_37), .A (n_35_39), .B (n_32_39), .C1 (n_28_41), .C2 (n_22_44) );
AOI211_X1 g_41_36 (.ZN (n_41_36), .A (n_37_38), .B (n_31_41), .C1 (n_30_40), .C2 (n_24_43) );
AOI211_X1 g_40_38 (.ZN (n_40_38), .A (n_39_37), .B (n_33_40), .C1 (n_32_39), .C2 (n_26_42) );
AOI211_X1 g_39_36 (.ZN (n_39_36), .A (n_41_36), .B (n_35_39), .C1 (n_31_41), .C2 (n_28_41) );
AOI211_X1 g_41_35 (.ZN (n_41_35), .A (n_40_38), .B (n_37_38), .C1 (n_33_40), .C2 (n_30_40) );
AOI211_X1 g_43_34 (.ZN (n_43_34), .A (n_39_36), .B (n_39_37), .C1 (n_35_39), .C2 (n_32_39) );
AOI211_X1 g_45_33 (.ZN (n_45_33), .A (n_41_35), .B (n_41_36), .C1 (n_37_38), .C2 (n_31_41) );
AOI211_X1 g_47_32 (.ZN (n_47_32), .A (n_43_34), .B (n_40_38), .C1 (n_39_37), .C2 (n_33_40) );
AOI211_X1 g_49_31 (.ZN (n_49_31), .A (n_45_33), .B (n_39_36), .C1 (n_41_36), .C2 (n_35_39) );
AOI211_X1 g_51_30 (.ZN (n_51_30), .A (n_47_32), .B (n_41_35), .C1 (n_40_38), .C2 (n_37_38) );
AOI211_X1 g_53_29 (.ZN (n_53_29), .A (n_49_31), .B (n_43_34), .C1 (n_39_36), .C2 (n_39_37) );
AOI211_X1 g_55_28 (.ZN (n_55_28), .A (n_51_30), .B (n_45_33), .C1 (n_41_35), .C2 (n_41_36) );
AOI211_X1 g_57_27 (.ZN (n_57_27), .A (n_53_29), .B (n_47_32), .C1 (n_43_34), .C2 (n_40_38) );
AOI211_X1 g_59_26 (.ZN (n_59_26), .A (n_55_28), .B (n_49_31), .C1 (n_45_33), .C2 (n_39_36) );
AOI211_X1 g_61_25 (.ZN (n_61_25), .A (n_57_27), .B (n_51_30), .C1 (n_47_32), .C2 (n_41_35) );
AOI211_X1 g_63_24 (.ZN (n_63_24), .A (n_59_26), .B (n_53_29), .C1 (n_49_31), .C2 (n_43_34) );
AOI211_X1 g_65_23 (.ZN (n_65_23), .A (n_61_25), .B (n_55_28), .C1 (n_51_30), .C2 (n_45_33) );
AOI211_X1 g_67_22 (.ZN (n_67_22), .A (n_63_24), .B (n_57_27), .C1 (n_53_29), .C2 (n_47_32) );
AOI211_X1 g_69_21 (.ZN (n_69_21), .A (n_65_23), .B (n_59_26), .C1 (n_55_28), .C2 (n_49_31) );
AOI211_X1 g_68_23 (.ZN (n_68_23), .A (n_67_22), .B (n_61_25), .C1 (n_57_27), .C2 (n_51_30) );
AOI211_X1 g_70_22 (.ZN (n_70_22), .A (n_69_21), .B (n_63_24), .C1 (n_59_26), .C2 (n_53_29) );
AOI211_X1 g_72_21 (.ZN (n_72_21), .A (n_68_23), .B (n_65_23), .C1 (n_61_25), .C2 (n_55_28) );
AOI211_X1 g_71_23 (.ZN (n_71_23), .A (n_70_22), .B (n_67_22), .C1 (n_63_24), .C2 (n_57_27) );
AOI211_X1 g_69_22 (.ZN (n_69_22), .A (n_72_21), .B (n_69_21), .C1 (n_65_23), .C2 (n_59_26) );
AOI211_X1 g_71_21 (.ZN (n_71_21), .A (n_71_23), .B (n_68_23), .C1 (n_67_22), .C2 (n_61_25) );
AOI211_X1 g_73_20 (.ZN (n_73_20), .A (n_69_22), .B (n_70_22), .C1 (n_69_21), .C2 (n_63_24) );
AOI211_X1 g_72_22 (.ZN (n_72_22), .A (n_71_21), .B (n_72_21), .C1 (n_68_23), .C2 (n_65_23) );
AOI211_X1 g_70_23 (.ZN (n_70_23), .A (n_73_20), .B (n_71_23), .C1 (n_70_22), .C2 (n_67_22) );
AOI211_X1 g_68_22 (.ZN (n_68_22), .A (n_72_22), .B (n_69_22), .C1 (n_72_21), .C2 (n_69_21) );
AOI211_X1 g_66_23 (.ZN (n_66_23), .A (n_70_23), .B (n_71_21), .C1 (n_71_23), .C2 (n_68_23) );
AOI211_X1 g_64_24 (.ZN (n_64_24), .A (n_68_22), .B (n_73_20), .C1 (n_69_22), .C2 (n_70_22) );
AOI211_X1 g_62_25 (.ZN (n_62_25), .A (n_66_23), .B (n_72_22), .C1 (n_71_21), .C2 (n_72_21) );
AOI211_X1 g_60_26 (.ZN (n_60_26), .A (n_64_24), .B (n_70_23), .C1 (n_73_20), .C2 (n_71_23) );
AOI211_X1 g_58_27 (.ZN (n_58_27), .A (n_62_25), .B (n_68_22), .C1 (n_72_22), .C2 (n_69_22) );
AOI211_X1 g_56_28 (.ZN (n_56_28), .A (n_60_26), .B (n_66_23), .C1 (n_70_23), .C2 (n_71_21) );
AOI211_X1 g_54_29 (.ZN (n_54_29), .A (n_58_27), .B (n_64_24), .C1 (n_68_22), .C2 (n_73_20) );
AOI211_X1 g_52_30 (.ZN (n_52_30), .A (n_56_28), .B (n_62_25), .C1 (n_66_23), .C2 (n_72_22) );
AOI211_X1 g_50_31 (.ZN (n_50_31), .A (n_54_29), .B (n_60_26), .C1 (n_64_24), .C2 (n_70_23) );
AOI211_X1 g_48_32 (.ZN (n_48_32), .A (n_52_30), .B (n_58_27), .C1 (n_62_25), .C2 (n_68_22) );
AOI211_X1 g_46_33 (.ZN (n_46_33), .A (n_50_31), .B (n_56_28), .C1 (n_60_26), .C2 (n_66_23) );
AOI211_X1 g_44_34 (.ZN (n_44_34), .A (n_48_32), .B (n_54_29), .C1 (n_58_27), .C2 (n_64_24) );
AOI211_X1 g_42_35 (.ZN (n_42_35), .A (n_46_33), .B (n_52_30), .C1 (n_56_28), .C2 (n_62_25) );
AOI211_X1 g_40_36 (.ZN (n_40_36), .A (n_44_34), .B (n_50_31), .C1 (n_54_29), .C2 (n_60_26) );
AOI211_X1 g_38_37 (.ZN (n_38_37), .A (n_42_35), .B (n_48_32), .C1 (n_52_30), .C2 (n_58_27) );
AOI211_X1 g_36_38 (.ZN (n_36_38), .A (n_40_36), .B (n_46_33), .C1 (n_50_31), .C2 (n_56_28) );
AOI211_X1 g_38_39 (.ZN (n_38_39), .A (n_38_37), .B (n_44_34), .C1 (n_48_32), .C2 (n_54_29) );
AOI211_X1 g_37_37 (.ZN (n_37_37), .A (n_36_38), .B (n_42_35), .C1 (n_46_33), .C2 (n_52_30) );
AOI211_X1 g_35_38 (.ZN (n_35_38), .A (n_38_39), .B (n_40_36), .C1 (n_44_34), .C2 (n_50_31) );
AOI211_X1 g_33_39 (.ZN (n_33_39), .A (n_37_37), .B (n_38_37), .C1 (n_42_35), .C2 (n_48_32) );
AOI211_X1 g_31_40 (.ZN (n_31_40), .A (n_35_38), .B (n_36_38), .C1 (n_40_36), .C2 (n_46_33) );
AOI211_X1 g_29_41 (.ZN (n_29_41), .A (n_33_39), .B (n_38_39), .C1 (n_38_37), .C2 (n_44_34) );
AOI211_X1 g_27_42 (.ZN (n_27_42), .A (n_31_40), .B (n_37_37), .C1 (n_36_38), .C2 (n_42_35) );
AOI211_X1 g_25_43 (.ZN (n_25_43), .A (n_29_41), .B (n_35_38), .C1 (n_38_39), .C2 (n_40_36) );
AOI211_X1 g_23_44 (.ZN (n_23_44), .A (n_27_42), .B (n_33_39), .C1 (n_37_37), .C2 (n_38_37) );
AOI211_X1 g_21_45 (.ZN (n_21_45), .A (n_25_43), .B (n_31_40), .C1 (n_35_38), .C2 (n_36_38) );
AOI211_X1 g_23_46 (.ZN (n_23_46), .A (n_23_44), .B (n_29_41), .C1 (n_33_39), .C2 (n_38_39) );
AOI211_X1 g_25_45 (.ZN (n_25_45), .A (n_21_45), .B (n_27_42), .C1 (n_31_40), .C2 (n_37_37) );
AOI211_X1 g_27_44 (.ZN (n_27_44), .A (n_23_46), .B (n_25_43), .C1 (n_29_41), .C2 (n_35_38) );
AOI211_X1 g_29_43 (.ZN (n_29_43), .A (n_25_45), .B (n_23_44), .C1 (n_27_42), .C2 (n_33_39) );
AOI211_X1 g_31_42 (.ZN (n_31_42), .A (n_27_44), .B (n_21_45), .C1 (n_25_43), .C2 (n_31_40) );
AOI211_X1 g_33_41 (.ZN (n_33_41), .A (n_29_43), .B (n_23_46), .C1 (n_23_44), .C2 (n_29_41) );
AOI211_X1 g_35_40 (.ZN (n_35_40), .A (n_31_42), .B (n_25_45), .C1 (n_21_45), .C2 (n_27_42) );
AOI211_X1 g_37_39 (.ZN (n_37_39), .A (n_33_41), .B (n_27_44), .C1 (n_23_46), .C2 (n_25_43) );
AOI211_X1 g_39_38 (.ZN (n_39_38), .A (n_35_40), .B (n_29_43), .C1 (n_25_45), .C2 (n_23_44) );
AOI211_X1 g_41_37 (.ZN (n_41_37), .A (n_37_39), .B (n_31_42), .C1 (n_27_44), .C2 (n_21_45) );
AOI211_X1 g_43_36 (.ZN (n_43_36), .A (n_39_38), .B (n_33_41), .C1 (n_29_43), .C2 (n_23_46) );
AOI211_X1 g_45_35 (.ZN (n_45_35), .A (n_41_37), .B (n_35_40), .C1 (n_31_42), .C2 (n_25_45) );
AOI211_X1 g_47_34 (.ZN (n_47_34), .A (n_43_36), .B (n_37_39), .C1 (n_33_41), .C2 (n_27_44) );
AOI211_X1 g_49_33 (.ZN (n_49_33), .A (n_45_35), .B (n_39_38), .C1 (n_35_40), .C2 (n_29_43) );
AOI211_X1 g_51_32 (.ZN (n_51_32), .A (n_47_34), .B (n_41_37), .C1 (n_37_39), .C2 (n_31_42) );
AOI211_X1 g_53_31 (.ZN (n_53_31), .A (n_49_33), .B (n_43_36), .C1 (n_39_38), .C2 (n_33_41) );
AOI211_X1 g_55_30 (.ZN (n_55_30), .A (n_51_32), .B (n_45_35), .C1 (n_41_37), .C2 (n_35_40) );
AOI211_X1 g_57_29 (.ZN (n_57_29), .A (n_53_31), .B (n_47_34), .C1 (n_43_36), .C2 (n_37_39) );
AOI211_X1 g_59_28 (.ZN (n_59_28), .A (n_55_30), .B (n_49_33), .C1 (n_45_35), .C2 (n_39_38) );
AOI211_X1 g_61_27 (.ZN (n_61_27), .A (n_57_29), .B (n_51_32), .C1 (n_47_34), .C2 (n_41_37) );
AOI211_X1 g_63_26 (.ZN (n_63_26), .A (n_59_28), .B (n_53_31), .C1 (n_49_33), .C2 (n_43_36) );
AOI211_X1 g_65_25 (.ZN (n_65_25), .A (n_61_27), .B (n_55_30), .C1 (n_51_32), .C2 (n_45_35) );
AOI211_X1 g_67_24 (.ZN (n_67_24), .A (n_63_26), .B (n_57_29), .C1 (n_53_31), .C2 (n_47_34) );
AOI211_X1 g_69_23 (.ZN (n_69_23), .A (n_65_25), .B (n_59_28), .C1 (n_55_30), .C2 (n_49_33) );
AOI211_X1 g_71_22 (.ZN (n_71_22), .A (n_67_24), .B (n_61_27), .C1 (n_57_29), .C2 (n_51_32) );
AOI211_X1 g_73_21 (.ZN (n_73_21), .A (n_69_23), .B (n_63_26), .C1 (n_59_28), .C2 (n_53_31) );
AOI211_X1 g_72_23 (.ZN (n_72_23), .A (n_71_22), .B (n_65_25), .C1 (n_61_27), .C2 (n_55_30) );
AOI211_X1 g_74_22 (.ZN (n_74_22), .A (n_73_21), .B (n_67_24), .C1 (n_63_26), .C2 (n_57_29) );
AOI211_X1 g_76_21 (.ZN (n_76_21), .A (n_72_23), .B (n_69_23), .C1 (n_65_25), .C2 (n_59_28) );
AOI211_X1 g_78_20 (.ZN (n_78_20), .A (n_74_22), .B (n_71_22), .C1 (n_67_24), .C2 (n_61_27) );
AOI211_X1 g_80_19 (.ZN (n_80_19), .A (n_76_21), .B (n_73_21), .C1 (n_69_23), .C2 (n_63_26) );
AOI211_X1 g_82_18 (.ZN (n_82_18), .A (n_78_20), .B (n_72_23), .C1 (n_71_22), .C2 (n_65_25) );
AOI211_X1 g_84_17 (.ZN (n_84_17), .A (n_80_19), .B (n_74_22), .C1 (n_73_21), .C2 (n_67_24) );
AOI211_X1 g_86_16 (.ZN (n_86_16), .A (n_82_18), .B (n_76_21), .C1 (n_72_23), .C2 (n_69_23) );
AOI211_X1 g_88_15 (.ZN (n_88_15), .A (n_84_17), .B (n_78_20), .C1 (n_74_22), .C2 (n_71_22) );
AOI211_X1 g_90_14 (.ZN (n_90_14), .A (n_86_16), .B (n_80_19), .C1 (n_76_21), .C2 (n_73_21) );
AOI211_X1 g_92_13 (.ZN (n_92_13), .A (n_88_15), .B (n_82_18), .C1 (n_78_20), .C2 (n_72_23) );
AOI211_X1 g_93_11 (.ZN (n_93_11), .A (n_90_14), .B (n_84_17), .C1 (n_80_19), .C2 (n_74_22) );
AOI211_X1 g_95_10 (.ZN (n_95_10), .A (n_92_13), .B (n_86_16), .C1 (n_82_18), .C2 (n_76_21) );
AOI211_X1 g_97_9 (.ZN (n_97_9), .A (n_93_11), .B (n_88_15), .C1 (n_84_17), .C2 (n_78_20) );
AOI211_X1 g_96_11 (.ZN (n_96_11), .A (n_95_10), .B (n_90_14), .C1 (n_86_16), .C2 (n_80_19) );
AOI211_X1 g_94_12 (.ZN (n_94_12), .A (n_97_9), .B (n_92_13), .C1 (n_88_15), .C2 (n_82_18) );
AOI211_X1 g_93_14 (.ZN (n_93_14), .A (n_96_11), .B (n_93_11), .C1 (n_90_14), .C2 (n_84_17) );
AOI211_X1 g_91_15 (.ZN (n_91_15), .A (n_94_12), .B (n_95_10), .C1 (n_92_13), .C2 (n_86_16) );
AOI211_X1 g_89_16 (.ZN (n_89_16), .A (n_93_14), .B (n_97_9), .C1 (n_93_11), .C2 (n_88_15) );
AOI211_X1 g_87_17 (.ZN (n_87_17), .A (n_91_15), .B (n_96_11), .C1 (n_95_10), .C2 (n_90_14) );
AOI211_X1 g_86_15 (.ZN (n_86_15), .A (n_89_16), .B (n_94_12), .C1 (n_97_9), .C2 (n_92_13) );
AOI211_X1 g_84_16 (.ZN (n_84_16), .A (n_87_17), .B (n_93_14), .C1 (n_96_11), .C2 (n_93_11) );
AOI211_X1 g_82_17 (.ZN (n_82_17), .A (n_86_15), .B (n_91_15), .C1 (n_94_12), .C2 (n_95_10) );
AOI211_X1 g_80_18 (.ZN (n_80_18), .A (n_84_16), .B (n_89_16), .C1 (n_93_14), .C2 (n_97_9) );
AOI211_X1 g_78_19 (.ZN (n_78_19), .A (n_82_17), .B (n_87_17), .C1 (n_91_15), .C2 (n_96_11) );
AOI211_X1 g_76_20 (.ZN (n_76_20), .A (n_80_18), .B (n_86_15), .C1 (n_89_16), .C2 (n_94_12) );
AOI211_X1 g_75_22 (.ZN (n_75_22), .A (n_78_19), .B (n_84_16), .C1 (n_87_17), .C2 (n_93_14) );
AOI211_X1 g_77_21 (.ZN (n_77_21), .A (n_76_20), .B (n_82_17), .C1 (n_86_15), .C2 (n_91_15) );
AOI211_X1 g_79_20 (.ZN (n_79_20), .A (n_75_22), .B (n_80_18), .C1 (n_84_16), .C2 (n_89_16) );
AOI211_X1 g_81_19 (.ZN (n_81_19), .A (n_77_21), .B (n_78_19), .C1 (n_82_17), .C2 (n_87_17) );
AOI211_X1 g_83_18 (.ZN (n_83_18), .A (n_79_20), .B (n_76_20), .C1 (n_80_18), .C2 (n_86_15) );
AOI211_X1 g_85_17 (.ZN (n_85_17), .A (n_81_19), .B (n_75_22), .C1 (n_78_19), .C2 (n_84_16) );
AOI211_X1 g_87_16 (.ZN (n_87_16), .A (n_83_18), .B (n_77_21), .C1 (n_76_20), .C2 (n_82_17) );
AOI211_X1 g_86_18 (.ZN (n_86_18), .A (n_85_17), .B (n_79_20), .C1 (n_75_22), .C2 (n_80_18) );
AOI211_X1 g_88_17 (.ZN (n_88_17), .A (n_87_16), .B (n_81_19), .C1 (n_77_21), .C2 (n_78_19) );
AOI211_X1 g_90_16 (.ZN (n_90_16), .A (n_86_18), .B (n_83_18), .C1 (n_79_20), .C2 (n_76_20) );
AOI211_X1 g_91_14 (.ZN (n_91_14), .A (n_88_17), .B (n_85_17), .C1 (n_81_19), .C2 (n_75_22) );
AOI211_X1 g_93_13 (.ZN (n_93_13), .A (n_90_16), .B (n_87_16), .C1 (n_83_18), .C2 (n_77_21) );
AOI211_X1 g_95_12 (.ZN (n_95_12), .A (n_91_14), .B (n_86_18), .C1 (n_85_17), .C2 (n_79_20) );
AOI211_X1 g_97_11 (.ZN (n_97_11), .A (n_93_13), .B (n_88_17), .C1 (n_87_16), .C2 (n_81_19) );
AOI211_X1 g_99_10 (.ZN (n_99_10), .A (n_95_12), .B (n_90_16), .C1 (n_86_18), .C2 (n_83_18) );
AOI211_X1 g_98_12 (.ZN (n_98_12), .A (n_97_11), .B (n_91_14), .C1 (n_88_17), .C2 (n_85_17) );
AOI211_X1 g_96_13 (.ZN (n_96_13), .A (n_99_10), .B (n_93_13), .C1 (n_90_16), .C2 (n_87_16) );
AOI211_X1 g_94_14 (.ZN (n_94_14), .A (n_98_12), .B (n_95_12), .C1 (n_91_14), .C2 (n_86_18) );
AOI211_X1 g_92_15 (.ZN (n_92_15), .A (n_96_13), .B (n_97_11), .C1 (n_93_13), .C2 (n_88_17) );
AOI211_X1 g_91_17 (.ZN (n_91_17), .A (n_94_14), .B (n_99_10), .C1 (n_95_12), .C2 (n_90_16) );
AOI211_X1 g_90_15 (.ZN (n_90_15), .A (n_92_15), .B (n_98_12), .C1 (n_97_11), .C2 (n_91_14) );
AOI211_X1 g_92_14 (.ZN (n_92_14), .A (n_91_17), .B (n_96_13), .C1 (n_99_10), .C2 (n_93_13) );
AOI211_X1 g_94_13 (.ZN (n_94_13), .A (n_90_15), .B (n_94_14), .C1 (n_98_12), .C2 (n_95_12) );
AOI211_X1 g_96_12 (.ZN (n_96_12), .A (n_92_14), .B (n_92_15), .C1 (n_96_13), .C2 (n_97_11) );
AOI211_X1 g_98_11 (.ZN (n_98_11), .A (n_94_13), .B (n_91_17), .C1 (n_94_14), .C2 (n_99_10) );
AOI211_X1 g_100_12 (.ZN (n_100_12), .A (n_96_12), .B (n_90_15), .C1 (n_92_15), .C2 (n_98_12) );
AOI211_X1 g_98_13 (.ZN (n_98_13), .A (n_98_11), .B (n_92_14), .C1 (n_91_17), .C2 (n_96_13) );
AOI211_X1 g_96_14 (.ZN (n_96_14), .A (n_100_12), .B (n_94_13), .C1 (n_90_15), .C2 (n_94_14) );
AOI211_X1 g_94_15 (.ZN (n_94_15), .A (n_98_13), .B (n_96_12), .C1 (n_92_14), .C2 (n_92_15) );
AOI211_X1 g_92_16 (.ZN (n_92_16), .A (n_96_14), .B (n_98_11), .C1 (n_94_13), .C2 (n_91_17) );
AOI211_X1 g_90_17 (.ZN (n_90_17), .A (n_94_15), .B (n_100_12), .C1 (n_96_12), .C2 (n_90_15) );
AOI211_X1 g_88_16 (.ZN (n_88_16), .A (n_92_16), .B (n_98_13), .C1 (n_98_11), .C2 (n_92_14) );
AOI211_X1 g_86_17 (.ZN (n_86_17), .A (n_90_17), .B (n_96_14), .C1 (n_100_12), .C2 (n_94_13) );
AOI211_X1 g_84_18 (.ZN (n_84_18), .A (n_88_16), .B (n_94_15), .C1 (n_98_13), .C2 (n_96_12) );
AOI211_X1 g_82_19 (.ZN (n_82_19), .A (n_86_17), .B (n_92_16), .C1 (n_96_14), .C2 (n_98_11) );
AOI211_X1 g_83_17 (.ZN (n_83_17), .A (n_84_18), .B (n_90_17), .C1 (n_94_15), .C2 (n_100_12) );
AOI211_X1 g_81_18 (.ZN (n_81_18), .A (n_82_19), .B (n_88_16), .C1 (n_92_16), .C2 (n_98_13) );
AOI211_X1 g_79_19 (.ZN (n_79_19), .A (n_83_17), .B (n_86_17), .C1 (n_90_17), .C2 (n_96_14) );
AOI211_X1 g_77_20 (.ZN (n_77_20), .A (n_81_18), .B (n_84_18), .C1 (n_88_16), .C2 (n_94_15) );
AOI211_X1 g_75_21 (.ZN (n_75_21), .A (n_79_19), .B (n_82_19), .C1 (n_86_17), .C2 (n_92_16) );
AOI211_X1 g_73_22 (.ZN (n_73_22), .A (n_77_20), .B (n_83_17), .C1 (n_84_18), .C2 (n_90_17) );
AOI211_X1 g_72_24 (.ZN (n_72_24), .A (n_75_21), .B (n_81_18), .C1 (n_82_19), .C2 (n_88_16) );
AOI211_X1 g_74_23 (.ZN (n_74_23), .A (n_73_22), .B (n_79_19), .C1 (n_83_17), .C2 (n_86_17) );
AOI211_X1 g_76_22 (.ZN (n_76_22), .A (n_72_24), .B (n_77_20), .C1 (n_81_18), .C2 (n_84_18) );
AOI211_X1 g_78_21 (.ZN (n_78_21), .A (n_74_23), .B (n_75_21), .C1 (n_79_19), .C2 (n_82_19) );
AOI211_X1 g_80_20 (.ZN (n_80_20), .A (n_76_22), .B (n_73_22), .C1 (n_77_20), .C2 (n_83_17) );
AOI211_X1 g_79_22 (.ZN (n_79_22), .A (n_78_21), .B (n_72_24), .C1 (n_75_21), .C2 (n_81_18) );
AOI211_X1 g_81_21 (.ZN (n_81_21), .A (n_80_20), .B (n_74_23), .C1 (n_73_22), .C2 (n_79_19) );
AOI211_X1 g_83_20 (.ZN (n_83_20), .A (n_79_22), .B (n_76_22), .C1 (n_72_24), .C2 (n_77_20) );
AOI211_X1 g_85_19 (.ZN (n_85_19), .A (n_81_21), .B (n_78_21), .C1 (n_74_23), .C2 (n_75_21) );
AOI211_X1 g_87_18 (.ZN (n_87_18), .A (n_83_20), .B (n_80_20), .C1 (n_76_22), .C2 (n_73_22) );
AOI211_X1 g_89_17 (.ZN (n_89_17), .A (n_85_19), .B (n_79_22), .C1 (n_78_21), .C2 (n_72_24) );
AOI211_X1 g_91_16 (.ZN (n_91_16), .A (n_87_18), .B (n_81_21), .C1 (n_80_20), .C2 (n_74_23) );
AOI211_X1 g_93_15 (.ZN (n_93_15), .A (n_89_17), .B (n_83_20), .C1 (n_79_22), .C2 (n_76_22) );
AOI211_X1 g_95_14 (.ZN (n_95_14), .A (n_91_16), .B (n_85_19), .C1 (n_81_21), .C2 (n_78_21) );
AOI211_X1 g_97_13 (.ZN (n_97_13), .A (n_93_15), .B (n_87_18), .C1 (n_83_20), .C2 (n_80_20) );
AOI211_X1 g_99_14 (.ZN (n_99_14), .A (n_95_14), .B (n_89_17), .C1 (n_85_19), .C2 (n_79_22) );
AOI211_X1 g_97_15 (.ZN (n_97_15), .A (n_97_13), .B (n_91_16), .C1 (n_87_18), .C2 (n_81_21) );
AOI211_X1 g_95_16 (.ZN (n_95_16), .A (n_99_14), .B (n_93_15), .C1 (n_89_17), .C2 (n_83_20) );
AOI211_X1 g_93_17 (.ZN (n_93_17), .A (n_97_15), .B (n_95_14), .C1 (n_91_16), .C2 (n_85_19) );
AOI211_X1 g_91_18 (.ZN (n_91_18), .A (n_95_16), .B (n_97_13), .C1 (n_93_15), .C2 (n_87_18) );
AOI211_X1 g_89_19 (.ZN (n_89_19), .A (n_93_17), .B (n_99_14), .C1 (n_95_14), .C2 (n_89_17) );
AOI211_X1 g_87_20 (.ZN (n_87_20), .A (n_91_18), .B (n_97_15), .C1 (n_97_13), .C2 (n_91_16) );
AOI211_X1 g_88_18 (.ZN (n_88_18), .A (n_89_19), .B (n_95_16), .C1 (n_99_14), .C2 (n_93_15) );
AOI211_X1 g_86_19 (.ZN (n_86_19), .A (n_87_20), .B (n_93_17), .C1 (n_97_15), .C2 (n_95_14) );
AOI211_X1 g_84_20 (.ZN (n_84_20), .A (n_88_18), .B (n_91_18), .C1 (n_95_16), .C2 (n_97_13) );
AOI211_X1 g_85_18 (.ZN (n_85_18), .A (n_86_19), .B (n_89_19), .C1 (n_93_17), .C2 (n_99_14) );
AOI211_X1 g_83_19 (.ZN (n_83_19), .A (n_84_20), .B (n_87_20), .C1 (n_91_18), .C2 (n_97_15) );
AOI211_X1 g_81_20 (.ZN (n_81_20), .A (n_85_18), .B (n_88_18), .C1 (n_89_19), .C2 (n_95_16) );
AOI211_X1 g_79_21 (.ZN (n_79_21), .A (n_83_19), .B (n_86_19), .C1 (n_87_20), .C2 (n_93_17) );
AOI211_X1 g_77_22 (.ZN (n_77_22), .A (n_81_20), .B (n_84_20), .C1 (n_88_18), .C2 (n_91_18) );
AOI211_X1 g_75_23 (.ZN (n_75_23), .A (n_79_21), .B (n_85_18), .C1 (n_86_19), .C2 (n_89_19) );
AOI211_X1 g_73_24 (.ZN (n_73_24), .A (n_77_22), .B (n_83_19), .C1 (n_84_20), .C2 (n_87_20) );
AOI211_X1 g_71_25 (.ZN (n_71_25), .A (n_75_23), .B (n_81_20), .C1 (n_85_18), .C2 (n_88_18) );
AOI211_X1 g_69_24 (.ZN (n_69_24), .A (n_73_24), .B (n_79_21), .C1 (n_83_19), .C2 (n_86_19) );
AOI211_X1 g_67_23 (.ZN (n_67_23), .A (n_71_25), .B (n_77_22), .C1 (n_81_20), .C2 (n_84_20) );
AOI211_X1 g_65_24 (.ZN (n_65_24), .A (n_69_24), .B (n_75_23), .C1 (n_79_21), .C2 (n_85_18) );
AOI211_X1 g_67_25 (.ZN (n_67_25), .A (n_67_23), .B (n_73_24), .C1 (n_77_22), .C2 (n_83_19) );
AOI211_X1 g_65_26 (.ZN (n_65_26), .A (n_65_24), .B (n_71_25), .C1 (n_75_23), .C2 (n_81_20) );
AOI211_X1 g_66_24 (.ZN (n_66_24), .A (n_67_25), .B (n_69_24), .C1 (n_73_24), .C2 (n_79_21) );
AOI211_X1 g_64_25 (.ZN (n_64_25), .A (n_65_26), .B (n_67_23), .C1 (n_71_25), .C2 (n_77_22) );
AOI211_X1 g_62_26 (.ZN (n_62_26), .A (n_66_24), .B (n_65_24), .C1 (n_69_24), .C2 (n_75_23) );
AOI211_X1 g_60_27 (.ZN (n_60_27), .A (n_64_25), .B (n_67_25), .C1 (n_67_23), .C2 (n_73_24) );
AOI211_X1 g_58_28 (.ZN (n_58_28), .A (n_62_26), .B (n_65_26), .C1 (n_65_24), .C2 (n_71_25) );
AOI211_X1 g_56_29 (.ZN (n_56_29), .A (n_60_27), .B (n_66_24), .C1 (n_67_25), .C2 (n_69_24) );
AOI211_X1 g_54_30 (.ZN (n_54_30), .A (n_58_28), .B (n_64_25), .C1 (n_65_26), .C2 (n_67_23) );
AOI211_X1 g_52_31 (.ZN (n_52_31), .A (n_56_29), .B (n_62_26), .C1 (n_66_24), .C2 (n_65_24) );
AOI211_X1 g_50_32 (.ZN (n_50_32), .A (n_54_30), .B (n_60_27), .C1 (n_64_25), .C2 (n_67_25) );
AOI211_X1 g_48_33 (.ZN (n_48_33), .A (n_52_31), .B (n_58_28), .C1 (n_62_26), .C2 (n_65_26) );
AOI211_X1 g_46_34 (.ZN (n_46_34), .A (n_50_32), .B (n_56_29), .C1 (n_60_27), .C2 (n_66_24) );
AOI211_X1 g_44_35 (.ZN (n_44_35), .A (n_48_33), .B (n_54_30), .C1 (n_58_28), .C2 (n_64_25) );
AOI211_X1 g_42_36 (.ZN (n_42_36), .A (n_46_34), .B (n_52_31), .C1 (n_56_29), .C2 (n_62_26) );
AOI211_X1 g_40_37 (.ZN (n_40_37), .A (n_44_35), .B (n_50_32), .C1 (n_54_30), .C2 (n_60_27) );
AOI211_X1 g_38_38 (.ZN (n_38_38), .A (n_42_36), .B (n_48_33), .C1 (n_52_31), .C2 (n_58_28) );
AOI211_X1 g_36_39 (.ZN (n_36_39), .A (n_40_37), .B (n_46_34), .C1 (n_50_32), .C2 (n_56_29) );
AOI211_X1 g_34_40 (.ZN (n_34_40), .A (n_38_38), .B (n_44_35), .C1 (n_48_33), .C2 (n_54_30) );
AOI211_X1 g_32_41 (.ZN (n_32_41), .A (n_36_39), .B (n_42_36), .C1 (n_46_34), .C2 (n_52_31) );
AOI211_X1 g_30_42 (.ZN (n_30_42), .A (n_34_40), .B (n_40_37), .C1 (n_44_35), .C2 (n_50_32) );
AOI211_X1 g_28_43 (.ZN (n_28_43), .A (n_32_41), .B (n_38_38), .C1 (n_42_36), .C2 (n_48_33) );
AOI211_X1 g_26_44 (.ZN (n_26_44), .A (n_30_42), .B (n_36_39), .C1 (n_40_37), .C2 (n_46_34) );
AOI211_X1 g_24_45 (.ZN (n_24_45), .A (n_28_43), .B (n_34_40), .C1 (n_38_38), .C2 (n_44_35) );
AOI211_X1 g_22_46 (.ZN (n_22_46), .A (n_26_44), .B (n_32_41), .C1 (n_36_39), .C2 (n_42_36) );
AOI211_X1 g_20_47 (.ZN (n_20_47), .A (n_24_45), .B (n_30_42), .C1 (n_34_40), .C2 (n_40_37) );
AOI211_X1 g_18_46 (.ZN (n_18_46), .A (n_22_46), .B (n_28_43), .C1 (n_32_41), .C2 (n_38_38) );
AOI211_X1 g_16_47 (.ZN (n_16_47), .A (n_20_47), .B (n_26_44), .C1 (n_30_42), .C2 (n_36_39) );
AOI211_X1 g_14_48 (.ZN (n_14_48), .A (n_18_46), .B (n_24_45), .C1 (n_28_43), .C2 (n_34_40) );
AOI211_X1 g_12_49 (.ZN (n_12_49), .A (n_16_47), .B (n_22_46), .C1 (n_26_44), .C2 (n_32_41) );
AOI211_X1 g_10_50 (.ZN (n_10_50), .A (n_14_48), .B (n_20_47), .C1 (n_24_45), .C2 (n_30_42) );
AOI211_X1 g_8_51 (.ZN (n_8_51), .A (n_12_49), .B (n_18_46), .C1 (n_22_46), .C2 (n_28_43) );
AOI211_X1 g_9_53 (.ZN (n_9_53), .A (n_10_50), .B (n_16_47), .C1 (n_20_47), .C2 (n_26_44) );
AOI211_X1 g_8_55 (.ZN (n_8_55), .A (n_8_51), .B (n_14_48), .C1 (n_18_46), .C2 (n_24_45) );
AOI211_X1 g_7_53 (.ZN (n_7_53), .A (n_9_53), .B (n_12_49), .C1 (n_16_47), .C2 (n_22_46) );
AOI211_X1 g_9_52 (.ZN (n_9_52), .A (n_8_55), .B (n_10_50), .C1 (n_14_48), .C2 (n_20_47) );
AOI211_X1 g_11_51 (.ZN (n_11_51), .A (n_7_53), .B (n_8_51), .C1 (n_12_49), .C2 (n_18_46) );
AOI211_X1 g_13_50 (.ZN (n_13_50), .A (n_9_52), .B (n_9_53), .C1 (n_10_50), .C2 (n_16_47) );
AOI211_X1 g_15_49 (.ZN (n_15_49), .A (n_11_51), .B (n_8_55), .C1 (n_8_51), .C2 (n_14_48) );
AOI211_X1 g_17_48 (.ZN (n_17_48), .A (n_13_50), .B (n_7_53), .C1 (n_9_53), .C2 (n_12_49) );
AOI211_X1 g_19_47 (.ZN (n_19_47), .A (n_15_49), .B (n_9_52), .C1 (n_8_55), .C2 (n_10_50) );
AOI211_X1 g_21_46 (.ZN (n_21_46), .A (n_17_48), .B (n_11_51), .C1 (n_7_53), .C2 (n_8_51) );
AOI211_X1 g_23_45 (.ZN (n_23_45), .A (n_19_47), .B (n_13_50), .C1 (n_9_52), .C2 (n_9_53) );
AOI211_X1 g_25_44 (.ZN (n_25_44), .A (n_21_46), .B (n_15_49), .C1 (n_11_51), .C2 (n_8_55) );
AOI211_X1 g_27_43 (.ZN (n_27_43), .A (n_23_45), .B (n_17_48), .C1 (n_13_50), .C2 (n_7_53) );
AOI211_X1 g_29_42 (.ZN (n_29_42), .A (n_25_44), .B (n_19_47), .C1 (n_15_49), .C2 (n_9_52) );
AOI211_X1 g_28_44 (.ZN (n_28_44), .A (n_27_43), .B (n_21_46), .C1 (n_17_48), .C2 (n_11_51) );
AOI211_X1 g_30_43 (.ZN (n_30_43), .A (n_29_42), .B (n_23_45), .C1 (n_19_47), .C2 (n_13_50) );
AOI211_X1 g_32_42 (.ZN (n_32_42), .A (n_28_44), .B (n_25_44), .C1 (n_21_46), .C2 (n_15_49) );
AOI211_X1 g_34_41 (.ZN (n_34_41), .A (n_30_43), .B (n_27_43), .C1 (n_23_45), .C2 (n_17_48) );
AOI211_X1 g_36_40 (.ZN (n_36_40), .A (n_32_42), .B (n_29_42), .C1 (n_25_44), .C2 (n_19_47) );
AOI211_X1 g_35_42 (.ZN (n_35_42), .A (n_34_41), .B (n_28_44), .C1 (n_27_43), .C2 (n_21_46) );
AOI211_X1 g_37_41 (.ZN (n_37_41), .A (n_36_40), .B (n_30_43), .C1 (n_29_42), .C2 (n_23_45) );
AOI211_X1 g_39_40 (.ZN (n_39_40), .A (n_35_42), .B (n_32_42), .C1 (n_28_44), .C2 (n_25_44) );
AOI211_X1 g_41_39 (.ZN (n_41_39), .A (n_37_41), .B (n_34_41), .C1 (n_30_43), .C2 (n_27_43) );
AOI211_X1 g_42_37 (.ZN (n_42_37), .A (n_39_40), .B (n_36_40), .C1 (n_32_42), .C2 (n_29_42) );
AOI211_X1 g_44_36 (.ZN (n_44_36), .A (n_41_39), .B (n_35_42), .C1 (n_34_41), .C2 (n_28_44) );
AOI211_X1 g_45_34 (.ZN (n_45_34), .A (n_42_37), .B (n_37_41), .C1 (n_36_40), .C2 (n_30_43) );
AOI211_X1 g_47_33 (.ZN (n_47_33), .A (n_44_36), .B (n_39_40), .C1 (n_35_42), .C2 (n_32_42) );
AOI211_X1 g_49_32 (.ZN (n_49_32), .A (n_45_34), .B (n_41_39), .C1 (n_37_41), .C2 (n_34_41) );
AOI211_X1 g_51_31 (.ZN (n_51_31), .A (n_47_33), .B (n_42_37), .C1 (n_39_40), .C2 (n_36_40) );
AOI211_X1 g_53_30 (.ZN (n_53_30), .A (n_49_32), .B (n_44_36), .C1 (n_41_39), .C2 (n_35_42) );
AOI211_X1 g_55_29 (.ZN (n_55_29), .A (n_51_31), .B (n_45_34), .C1 (n_42_37), .C2 (n_37_41) );
AOI211_X1 g_57_28 (.ZN (n_57_28), .A (n_53_30), .B (n_47_33), .C1 (n_44_36), .C2 (n_39_40) );
AOI211_X1 g_59_27 (.ZN (n_59_27), .A (n_55_29), .B (n_49_32), .C1 (n_45_34), .C2 (n_41_39) );
AOI211_X1 g_61_26 (.ZN (n_61_26), .A (n_57_28), .B (n_51_31), .C1 (n_47_33), .C2 (n_42_37) );
AOI211_X1 g_63_27 (.ZN (n_63_27), .A (n_59_27), .B (n_53_30), .C1 (n_49_32), .C2 (n_44_36) );
AOI211_X1 g_61_28 (.ZN (n_61_28), .A (n_61_26), .B (n_55_29), .C1 (n_51_31), .C2 (n_45_34) );
AOI211_X1 g_59_29 (.ZN (n_59_29), .A (n_63_27), .B (n_57_28), .C1 (n_53_30), .C2 (n_47_33) );
AOI211_X1 g_57_30 (.ZN (n_57_30), .A (n_61_28), .B (n_59_27), .C1 (n_55_29), .C2 (n_49_32) );
AOI211_X1 g_55_31 (.ZN (n_55_31), .A (n_59_29), .B (n_61_26), .C1 (n_57_28), .C2 (n_51_31) );
AOI211_X1 g_53_32 (.ZN (n_53_32), .A (n_57_30), .B (n_63_27), .C1 (n_59_27), .C2 (n_53_30) );
AOI211_X1 g_51_33 (.ZN (n_51_33), .A (n_55_31), .B (n_61_28), .C1 (n_61_26), .C2 (n_55_29) );
AOI211_X1 g_49_34 (.ZN (n_49_34), .A (n_53_32), .B (n_59_29), .C1 (n_63_27), .C2 (n_57_28) );
AOI211_X1 g_47_35 (.ZN (n_47_35), .A (n_51_33), .B (n_57_30), .C1 (n_61_28), .C2 (n_59_27) );
AOI211_X1 g_45_36 (.ZN (n_45_36), .A (n_49_34), .B (n_55_31), .C1 (n_59_29), .C2 (n_61_26) );
AOI211_X1 g_43_37 (.ZN (n_43_37), .A (n_47_35), .B (n_53_32), .C1 (n_57_30), .C2 (n_63_27) );
AOI211_X1 g_41_38 (.ZN (n_41_38), .A (n_45_36), .B (n_51_33), .C1 (n_55_31), .C2 (n_61_28) );
AOI211_X1 g_39_39 (.ZN (n_39_39), .A (n_43_37), .B (n_49_34), .C1 (n_53_32), .C2 (n_59_29) );
AOI211_X1 g_37_40 (.ZN (n_37_40), .A (n_41_38), .B (n_47_35), .C1 (n_51_33), .C2 (n_57_30) );
AOI211_X1 g_35_41 (.ZN (n_35_41), .A (n_39_39), .B (n_45_36), .C1 (n_49_34), .C2 (n_55_31) );
AOI211_X1 g_33_42 (.ZN (n_33_42), .A (n_37_40), .B (n_43_37), .C1 (n_47_35), .C2 (n_53_32) );
AOI211_X1 g_31_43 (.ZN (n_31_43), .A (n_35_41), .B (n_41_38), .C1 (n_45_36), .C2 (n_51_33) );
AOI211_X1 g_29_44 (.ZN (n_29_44), .A (n_33_42), .B (n_39_39), .C1 (n_43_37), .C2 (n_49_34) );
AOI211_X1 g_27_45 (.ZN (n_27_45), .A (n_31_43), .B (n_37_40), .C1 (n_41_38), .C2 (n_47_35) );
AOI211_X1 g_25_46 (.ZN (n_25_46), .A (n_29_44), .B (n_35_41), .C1 (n_39_39), .C2 (n_45_36) );
AOI211_X1 g_23_47 (.ZN (n_23_47), .A (n_27_45), .B (n_33_42), .C1 (n_37_40), .C2 (n_43_37) );
AOI211_X1 g_21_48 (.ZN (n_21_48), .A (n_25_46), .B (n_31_43), .C1 (n_35_41), .C2 (n_41_38) );
AOI211_X1 g_19_49 (.ZN (n_19_49), .A (n_23_47), .B (n_29_44), .C1 (n_33_42), .C2 (n_39_39) );
AOI211_X1 g_17_50 (.ZN (n_17_50), .A (n_21_48), .B (n_27_45), .C1 (n_31_43), .C2 (n_37_40) );
AOI211_X1 g_18_48 (.ZN (n_18_48), .A (n_19_49), .B (n_25_46), .C1 (n_29_44), .C2 (n_35_41) );
AOI211_X1 g_16_49 (.ZN (n_16_49), .A (n_17_50), .B (n_23_47), .C1 (n_27_45), .C2 (n_33_42) );
AOI211_X1 g_14_50 (.ZN (n_14_50), .A (n_18_48), .B (n_21_48), .C1 (n_25_46), .C2 (n_31_43) );
AOI211_X1 g_12_51 (.ZN (n_12_51), .A (n_16_49), .B (n_19_49), .C1 (n_23_47), .C2 (n_29_44) );
AOI211_X1 g_10_52 (.ZN (n_10_52), .A (n_14_50), .B (n_17_50), .C1 (n_21_48), .C2 (n_27_45) );
AOI211_X1 g_8_53 (.ZN (n_8_53), .A (n_12_51), .B (n_18_48), .C1 (n_19_49), .C2 (n_25_46) );
AOI211_X1 g_6_54 (.ZN (n_6_54), .A (n_10_52), .B (n_16_49), .C1 (n_17_50), .C2 (n_23_47) );
AOI211_X1 g_5_56 (.ZN (n_5_56), .A (n_8_53), .B (n_14_50), .C1 (n_18_48), .C2 (n_21_48) );
AOI211_X1 g_7_55 (.ZN (n_7_55), .A (n_6_54), .B (n_12_51), .C1 (n_16_49), .C2 (n_19_49) );
AOI211_X1 g_9_54 (.ZN (n_9_54), .A (n_5_56), .B (n_10_52), .C1 (n_14_50), .C2 (n_17_50) );
AOI211_X1 g_11_53 (.ZN (n_11_53), .A (n_7_55), .B (n_8_53), .C1 (n_12_51), .C2 (n_18_48) );
AOI211_X1 g_13_52 (.ZN (n_13_52), .A (n_9_54), .B (n_6_54), .C1 (n_10_52), .C2 (n_16_49) );
AOI211_X1 g_15_51 (.ZN (n_15_51), .A (n_11_53), .B (n_5_56), .C1 (n_8_53), .C2 (n_14_50) );
AOI211_X1 g_14_53 (.ZN (n_14_53), .A (n_13_52), .B (n_7_55), .C1 (n_6_54), .C2 (n_12_51) );
AOI211_X1 g_13_51 (.ZN (n_13_51), .A (n_15_51), .B (n_9_54), .C1 (n_5_56), .C2 (n_10_52) );
AOI211_X1 g_15_50 (.ZN (n_15_50), .A (n_14_53), .B (n_11_53), .C1 (n_7_55), .C2 (n_8_53) );
AOI211_X1 g_17_49 (.ZN (n_17_49), .A (n_13_51), .B (n_13_52), .C1 (n_9_54), .C2 (n_6_54) );
AOI211_X1 g_19_48 (.ZN (n_19_48), .A (n_15_50), .B (n_15_51), .C1 (n_11_53), .C2 (n_5_56) );
AOI211_X1 g_18_50 (.ZN (n_18_50), .A (n_17_49), .B (n_14_53), .C1 (n_13_52), .C2 (n_7_55) );
AOI211_X1 g_20_49 (.ZN (n_20_49), .A (n_19_48), .B (n_13_51), .C1 (n_15_51), .C2 (n_9_54) );
AOI211_X1 g_22_48 (.ZN (n_22_48), .A (n_18_50), .B (n_15_50), .C1 (n_14_53), .C2 (n_11_53) );
AOI211_X1 g_24_47 (.ZN (n_24_47), .A (n_20_49), .B (n_17_49), .C1 (n_13_51), .C2 (n_13_52) );
AOI211_X1 g_26_46 (.ZN (n_26_46), .A (n_22_48), .B (n_19_48), .C1 (n_15_50), .C2 (n_15_51) );
AOI211_X1 g_28_45 (.ZN (n_28_45), .A (n_24_47), .B (n_18_50), .C1 (n_17_49), .C2 (n_14_53) );
AOI211_X1 g_30_44 (.ZN (n_30_44), .A (n_26_46), .B (n_20_49), .C1 (n_19_48), .C2 (n_13_51) );
AOI211_X1 g_32_43 (.ZN (n_32_43), .A (n_28_45), .B (n_22_48), .C1 (n_18_50), .C2 (n_15_50) );
AOI211_X1 g_34_42 (.ZN (n_34_42), .A (n_30_44), .B (n_24_47), .C1 (n_20_49), .C2 (n_17_49) );
AOI211_X1 g_36_41 (.ZN (n_36_41), .A (n_32_43), .B (n_26_46), .C1 (n_22_48), .C2 (n_19_48) );
AOI211_X1 g_38_40 (.ZN (n_38_40), .A (n_34_42), .B (n_28_45), .C1 (n_24_47), .C2 (n_18_50) );
AOI211_X1 g_40_39 (.ZN (n_40_39), .A (n_36_41), .B (n_30_44), .C1 (n_26_46), .C2 (n_20_49) );
AOI211_X1 g_42_38 (.ZN (n_42_38), .A (n_38_40), .B (n_32_43), .C1 (n_28_45), .C2 (n_22_48) );
AOI211_X1 g_44_37 (.ZN (n_44_37), .A (n_40_39), .B (n_34_42), .C1 (n_30_44), .C2 (n_24_47) );
AOI211_X1 g_46_36 (.ZN (n_46_36), .A (n_42_38), .B (n_36_41), .C1 (n_32_43), .C2 (n_26_46) );
AOI211_X1 g_48_35 (.ZN (n_48_35), .A (n_44_37), .B (n_38_40), .C1 (n_34_42), .C2 (n_28_45) );
AOI211_X1 g_50_34 (.ZN (n_50_34), .A (n_46_36), .B (n_40_39), .C1 (n_36_41), .C2 (n_30_44) );
AOI211_X1 g_52_33 (.ZN (n_52_33), .A (n_48_35), .B (n_42_38), .C1 (n_38_40), .C2 (n_32_43) );
AOI211_X1 g_54_32 (.ZN (n_54_32), .A (n_50_34), .B (n_44_37), .C1 (n_40_39), .C2 (n_34_42) );
AOI211_X1 g_56_31 (.ZN (n_56_31), .A (n_52_33), .B (n_46_36), .C1 (n_42_38), .C2 (n_36_41) );
AOI211_X1 g_58_30 (.ZN (n_58_30), .A (n_54_32), .B (n_48_35), .C1 (n_44_37), .C2 (n_38_40) );
AOI211_X1 g_60_29 (.ZN (n_60_29), .A (n_56_31), .B (n_50_34), .C1 (n_46_36), .C2 (n_40_39) );
AOI211_X1 g_62_28 (.ZN (n_62_28), .A (n_58_30), .B (n_52_33), .C1 (n_48_35), .C2 (n_42_38) );
AOI211_X1 g_64_27 (.ZN (n_64_27), .A (n_60_29), .B (n_54_32), .C1 (n_50_34), .C2 (n_44_37) );
AOI211_X1 g_66_26 (.ZN (n_66_26), .A (n_62_28), .B (n_56_31), .C1 (n_52_33), .C2 (n_46_36) );
AOI211_X1 g_68_25 (.ZN (n_68_25), .A (n_64_27), .B (n_58_30), .C1 (n_54_32), .C2 (n_48_35) );
AOI211_X1 g_70_24 (.ZN (n_70_24), .A (n_66_26), .B (n_60_29), .C1 (n_56_31), .C2 (n_50_34) );
AOI211_X1 g_69_26 (.ZN (n_69_26), .A (n_68_25), .B (n_62_28), .C1 (n_58_30), .C2 (n_52_33) );
AOI211_X1 g_68_24 (.ZN (n_68_24), .A (n_70_24), .B (n_64_27), .C1 (n_60_29), .C2 (n_54_32) );
AOI211_X1 g_66_25 (.ZN (n_66_25), .A (n_69_26), .B (n_66_26), .C1 (n_62_28), .C2 (n_56_31) );
AOI211_X1 g_64_26 (.ZN (n_64_26), .A (n_68_24), .B (n_68_25), .C1 (n_64_27), .C2 (n_58_30) );
AOI211_X1 g_62_27 (.ZN (n_62_27), .A (n_66_25), .B (n_70_24), .C1 (n_66_26), .C2 (n_60_29) );
AOI211_X1 g_60_28 (.ZN (n_60_28), .A (n_64_26), .B (n_69_26), .C1 (n_68_25), .C2 (n_62_28) );
AOI211_X1 g_58_29 (.ZN (n_58_29), .A (n_62_27), .B (n_68_24), .C1 (n_70_24), .C2 (n_64_27) );
AOI211_X1 g_56_30 (.ZN (n_56_30), .A (n_60_28), .B (n_66_25), .C1 (n_69_26), .C2 (n_66_26) );
AOI211_X1 g_54_31 (.ZN (n_54_31), .A (n_58_29), .B (n_64_26), .C1 (n_68_24), .C2 (n_68_25) );
AOI211_X1 g_52_32 (.ZN (n_52_32), .A (n_56_30), .B (n_62_27), .C1 (n_66_25), .C2 (n_70_24) );
AOI211_X1 g_50_33 (.ZN (n_50_33), .A (n_54_31), .B (n_60_28), .C1 (n_64_26), .C2 (n_69_26) );
AOI211_X1 g_48_34 (.ZN (n_48_34), .A (n_52_32), .B (n_58_29), .C1 (n_62_27), .C2 (n_68_24) );
AOI211_X1 g_46_35 (.ZN (n_46_35), .A (n_50_33), .B (n_56_30), .C1 (n_60_28), .C2 (n_66_25) );
AOI211_X1 g_45_37 (.ZN (n_45_37), .A (n_48_34), .B (n_54_31), .C1 (n_58_29), .C2 (n_64_26) );
AOI211_X1 g_43_38 (.ZN (n_43_38), .A (n_46_35), .B (n_52_32), .C1 (n_56_30), .C2 (n_62_27) );
AOI211_X1 g_42_40 (.ZN (n_42_40), .A (n_45_37), .B (n_50_33), .C1 (n_54_31), .C2 (n_60_28) );
AOI211_X1 g_44_39 (.ZN (n_44_39), .A (n_43_38), .B (n_48_34), .C1 (n_52_32), .C2 (n_58_29) );
AOI211_X1 g_46_38 (.ZN (n_46_38), .A (n_42_40), .B (n_46_35), .C1 (n_50_33), .C2 (n_56_30) );
AOI211_X1 g_47_36 (.ZN (n_47_36), .A (n_44_39), .B (n_45_37), .C1 (n_48_34), .C2 (n_54_31) );
AOI211_X1 g_49_35 (.ZN (n_49_35), .A (n_46_38), .B (n_43_38), .C1 (n_46_35), .C2 (n_52_32) );
AOI211_X1 g_51_34 (.ZN (n_51_34), .A (n_47_36), .B (n_42_40), .C1 (n_45_37), .C2 (n_50_33) );
AOI211_X1 g_53_33 (.ZN (n_53_33), .A (n_49_35), .B (n_44_39), .C1 (n_43_38), .C2 (n_48_34) );
AOI211_X1 g_55_32 (.ZN (n_55_32), .A (n_51_34), .B (n_46_38), .C1 (n_42_40), .C2 (n_46_35) );
AOI211_X1 g_57_31 (.ZN (n_57_31), .A (n_53_33), .B (n_47_36), .C1 (n_44_39), .C2 (n_45_37) );
AOI211_X1 g_59_30 (.ZN (n_59_30), .A (n_55_32), .B (n_49_35), .C1 (n_46_38), .C2 (n_43_38) );
AOI211_X1 g_61_29 (.ZN (n_61_29), .A (n_57_31), .B (n_51_34), .C1 (n_47_36), .C2 (n_42_40) );
AOI211_X1 g_63_28 (.ZN (n_63_28), .A (n_59_30), .B (n_53_33), .C1 (n_49_35), .C2 (n_44_39) );
AOI211_X1 g_65_27 (.ZN (n_65_27), .A (n_61_29), .B (n_55_32), .C1 (n_51_34), .C2 (n_46_38) );
AOI211_X1 g_67_26 (.ZN (n_67_26), .A (n_63_28), .B (n_57_31), .C1 (n_53_33), .C2 (n_47_36) );
AOI211_X1 g_69_25 (.ZN (n_69_25), .A (n_65_27), .B (n_59_30), .C1 (n_55_32), .C2 (n_49_35) );
AOI211_X1 g_71_24 (.ZN (n_71_24), .A (n_67_26), .B (n_61_29), .C1 (n_57_31), .C2 (n_51_34) );
AOI211_X1 g_73_23 (.ZN (n_73_23), .A (n_69_25), .B (n_63_28), .C1 (n_59_30), .C2 (n_53_33) );
AOI211_X1 g_72_25 (.ZN (n_72_25), .A (n_71_24), .B (n_65_27), .C1 (n_61_29), .C2 (n_55_32) );
AOI211_X1 g_74_24 (.ZN (n_74_24), .A (n_73_23), .B (n_67_26), .C1 (n_63_28), .C2 (n_57_31) );
AOI211_X1 g_76_23 (.ZN (n_76_23), .A (n_72_25), .B (n_69_25), .C1 (n_65_27), .C2 (n_59_30) );
AOI211_X1 g_78_22 (.ZN (n_78_22), .A (n_74_24), .B (n_71_24), .C1 (n_67_26), .C2 (n_61_29) );
AOI211_X1 g_80_21 (.ZN (n_80_21), .A (n_76_23), .B (n_73_23), .C1 (n_69_25), .C2 (n_63_28) );
AOI211_X1 g_82_20 (.ZN (n_82_20), .A (n_78_22), .B (n_72_25), .C1 (n_71_24), .C2 (n_65_27) );
AOI211_X1 g_84_19 (.ZN (n_84_19), .A (n_80_21), .B (n_74_24), .C1 (n_73_23), .C2 (n_67_26) );
AOI211_X1 g_85_21 (.ZN (n_85_21), .A (n_82_20), .B (n_76_23), .C1 (n_72_25), .C2 (n_69_25) );
AOI211_X1 g_83_22 (.ZN (n_83_22), .A (n_84_19), .B (n_78_22), .C1 (n_74_24), .C2 (n_71_24) );
AOI211_X1 g_81_23 (.ZN (n_81_23), .A (n_85_21), .B (n_80_21), .C1 (n_76_23), .C2 (n_73_23) );
AOI211_X1 g_82_21 (.ZN (n_82_21), .A (n_83_22), .B (n_82_20), .C1 (n_78_22), .C2 (n_72_25) );
AOI211_X1 g_80_22 (.ZN (n_80_22), .A (n_81_23), .B (n_84_19), .C1 (n_80_21), .C2 (n_74_24) );
AOI211_X1 g_78_23 (.ZN (n_78_23), .A (n_82_21), .B (n_85_21), .C1 (n_82_20), .C2 (n_76_23) );
AOI211_X1 g_76_24 (.ZN (n_76_24), .A (n_80_22), .B (n_83_22), .C1 (n_84_19), .C2 (n_78_22) );
AOI211_X1 g_74_25 (.ZN (n_74_25), .A (n_78_23), .B (n_81_23), .C1 (n_85_21), .C2 (n_80_21) );
AOI211_X1 g_72_26 (.ZN (n_72_26), .A (n_76_24), .B (n_82_21), .C1 (n_83_22), .C2 (n_82_20) );
AOI211_X1 g_70_25 (.ZN (n_70_25), .A (n_74_25), .B (n_80_22), .C1 (n_81_23), .C2 (n_84_19) );
AOI211_X1 g_68_26 (.ZN (n_68_26), .A (n_72_26), .B (n_78_23), .C1 (n_82_21), .C2 (n_85_21) );
AOI211_X1 g_66_27 (.ZN (n_66_27), .A (n_70_25), .B (n_76_24), .C1 (n_80_22), .C2 (n_83_22) );
AOI211_X1 g_64_28 (.ZN (n_64_28), .A (n_68_26), .B (n_74_25), .C1 (n_78_23), .C2 (n_81_23) );
AOI211_X1 g_62_29 (.ZN (n_62_29), .A (n_66_27), .B (n_72_26), .C1 (n_76_24), .C2 (n_82_21) );
AOI211_X1 g_60_30 (.ZN (n_60_30), .A (n_64_28), .B (n_70_25), .C1 (n_74_25), .C2 (n_80_22) );
AOI211_X1 g_58_31 (.ZN (n_58_31), .A (n_62_29), .B (n_68_26), .C1 (n_72_26), .C2 (n_78_23) );
AOI211_X1 g_56_32 (.ZN (n_56_32), .A (n_60_30), .B (n_66_27), .C1 (n_70_25), .C2 (n_76_24) );
AOI211_X1 g_54_33 (.ZN (n_54_33), .A (n_58_31), .B (n_64_28), .C1 (n_68_26), .C2 (n_74_25) );
AOI211_X1 g_52_34 (.ZN (n_52_34), .A (n_56_32), .B (n_62_29), .C1 (n_66_27), .C2 (n_72_26) );
AOI211_X1 g_50_35 (.ZN (n_50_35), .A (n_54_33), .B (n_60_30), .C1 (n_64_28), .C2 (n_70_25) );
AOI211_X1 g_48_36 (.ZN (n_48_36), .A (n_52_34), .B (n_58_31), .C1 (n_62_29), .C2 (n_68_26) );
AOI211_X1 g_46_37 (.ZN (n_46_37), .A (n_50_35), .B (n_56_32), .C1 (n_60_30), .C2 (n_66_27) );
AOI211_X1 g_44_38 (.ZN (n_44_38), .A (n_48_36), .B (n_54_33), .C1 (n_58_31), .C2 (n_64_28) );
AOI211_X1 g_42_39 (.ZN (n_42_39), .A (n_46_37), .B (n_52_34), .C1 (n_56_32), .C2 (n_62_29) );
AOI211_X1 g_40_40 (.ZN (n_40_40), .A (n_44_38), .B (n_50_35), .C1 (n_54_33), .C2 (n_60_30) );
AOI211_X1 g_38_41 (.ZN (n_38_41), .A (n_42_39), .B (n_48_36), .C1 (n_52_34), .C2 (n_58_31) );
AOI211_X1 g_36_42 (.ZN (n_36_42), .A (n_40_40), .B (n_46_37), .C1 (n_50_35), .C2 (n_56_32) );
AOI211_X1 g_34_43 (.ZN (n_34_43), .A (n_38_41), .B (n_44_38), .C1 (n_48_36), .C2 (n_54_33) );
AOI211_X1 g_32_44 (.ZN (n_32_44), .A (n_36_42), .B (n_42_39), .C1 (n_46_37), .C2 (n_52_34) );
AOI211_X1 g_30_45 (.ZN (n_30_45), .A (n_34_43), .B (n_40_40), .C1 (n_44_38), .C2 (n_50_35) );
AOI211_X1 g_28_46 (.ZN (n_28_46), .A (n_32_44), .B (n_38_41), .C1 (n_42_39), .C2 (n_48_36) );
AOI211_X1 g_26_45 (.ZN (n_26_45), .A (n_30_45), .B (n_36_42), .C1 (n_40_40), .C2 (n_46_37) );
AOI211_X1 g_24_46 (.ZN (n_24_46), .A (n_28_46), .B (n_34_43), .C1 (n_38_41), .C2 (n_44_38) );
AOI211_X1 g_22_47 (.ZN (n_22_47), .A (n_26_45), .B (n_32_44), .C1 (n_36_42), .C2 (n_42_39) );
AOI211_X1 g_20_48 (.ZN (n_20_48), .A (n_24_46), .B (n_30_45), .C1 (n_34_43), .C2 (n_40_40) );
AOI211_X1 g_18_49 (.ZN (n_18_49), .A (n_22_47), .B (n_28_46), .C1 (n_32_44), .C2 (n_38_41) );
AOI211_X1 g_16_50 (.ZN (n_16_50), .A (n_20_48), .B (n_26_45), .C1 (n_30_45), .C2 (n_36_42) );
AOI211_X1 g_14_51 (.ZN (n_14_51), .A (n_18_49), .B (n_24_46), .C1 (n_28_46), .C2 (n_34_43) );
AOI211_X1 g_12_52 (.ZN (n_12_52), .A (n_16_50), .B (n_22_47), .C1 (n_26_45), .C2 (n_32_44) );
AOI211_X1 g_10_53 (.ZN (n_10_53), .A (n_14_51), .B (n_20_48), .C1 (n_24_46), .C2 (n_30_45) );
AOI211_X1 g_8_54 (.ZN (n_8_54), .A (n_12_52), .B (n_18_49), .C1 (n_22_47), .C2 (n_28_46) );
AOI211_X1 g_6_55 (.ZN (n_6_55), .A (n_10_53), .B (n_16_50), .C1 (n_20_48), .C2 (n_26_45) );
AOI211_X1 g_5_57 (.ZN (n_5_57), .A (n_8_54), .B (n_14_51), .C1 (n_18_49), .C2 (n_24_46) );
AOI211_X1 g_4_59 (.ZN (n_4_59), .A (n_6_55), .B (n_12_52), .C1 (n_16_50), .C2 (n_22_47) );
AOI211_X1 g_6_58 (.ZN (n_6_58), .A (n_5_57), .B (n_10_53), .C1 (n_14_51), .C2 (n_20_48) );
AOI211_X1 g_7_56 (.ZN (n_7_56), .A (n_4_59), .B (n_8_54), .C1 (n_12_52), .C2 (n_18_49) );
AOI211_X1 g_9_55 (.ZN (n_9_55), .A (n_6_58), .B (n_6_55), .C1 (n_10_53), .C2 (n_16_50) );
AOI211_X1 g_11_54 (.ZN (n_11_54), .A (n_7_56), .B (n_5_57), .C1 (n_8_54), .C2 (n_14_51) );
AOI211_X1 g_13_53 (.ZN (n_13_53), .A (n_9_55), .B (n_4_59), .C1 (n_6_55), .C2 (n_12_52) );
AOI211_X1 g_15_52 (.ZN (n_15_52), .A (n_11_54), .B (n_6_58), .C1 (n_5_57), .C2 (n_10_53) );
AOI211_X1 g_17_51 (.ZN (n_17_51), .A (n_13_53), .B (n_7_56), .C1 (n_4_59), .C2 (n_8_54) );
AOI211_X1 g_19_50 (.ZN (n_19_50), .A (n_15_52), .B (n_9_55), .C1 (n_6_58), .C2 (n_6_55) );
AOI211_X1 g_21_49 (.ZN (n_21_49), .A (n_17_51), .B (n_11_54), .C1 (n_7_56), .C2 (n_5_57) );
AOI211_X1 g_23_48 (.ZN (n_23_48), .A (n_19_50), .B (n_13_53), .C1 (n_9_55), .C2 (n_4_59) );
AOI211_X1 g_25_47 (.ZN (n_25_47), .A (n_21_49), .B (n_15_52), .C1 (n_11_54), .C2 (n_6_58) );
AOI211_X1 g_27_46 (.ZN (n_27_46), .A (n_23_48), .B (n_17_51), .C1 (n_13_53), .C2 (n_7_56) );
AOI211_X1 g_29_45 (.ZN (n_29_45), .A (n_25_47), .B (n_19_50), .C1 (n_15_52), .C2 (n_9_55) );
AOI211_X1 g_31_44 (.ZN (n_31_44), .A (n_27_46), .B (n_21_49), .C1 (n_17_51), .C2 (n_11_54) );
AOI211_X1 g_33_43 (.ZN (n_33_43), .A (n_29_45), .B (n_23_48), .C1 (n_19_50), .C2 (n_13_53) );
AOI211_X1 g_32_45 (.ZN (n_32_45), .A (n_31_44), .B (n_25_47), .C1 (n_21_49), .C2 (n_15_52) );
AOI211_X1 g_34_44 (.ZN (n_34_44), .A (n_33_43), .B (n_27_46), .C1 (n_23_48), .C2 (n_17_51) );
AOI211_X1 g_36_43 (.ZN (n_36_43), .A (n_32_45), .B (n_29_45), .C1 (n_25_47), .C2 (n_19_50) );
AOI211_X1 g_38_42 (.ZN (n_38_42), .A (n_34_44), .B (n_31_44), .C1 (n_27_46), .C2 (n_21_49) );
AOI211_X1 g_40_41 (.ZN (n_40_41), .A (n_36_43), .B (n_33_43), .C1 (n_29_45), .C2 (n_23_48) );
AOI211_X1 g_39_43 (.ZN (n_39_43), .A (n_38_42), .B (n_32_45), .C1 (n_31_44), .C2 (n_25_47) );
AOI211_X1 g_37_42 (.ZN (n_37_42), .A (n_40_41), .B (n_34_44), .C1 (n_33_43), .C2 (n_27_46) );
AOI211_X1 g_39_41 (.ZN (n_39_41), .A (n_39_43), .B (n_36_43), .C1 (n_32_45), .C2 (n_29_45) );
AOI211_X1 g_41_40 (.ZN (n_41_40), .A (n_37_42), .B (n_38_42), .C1 (n_34_44), .C2 (n_31_44) );
AOI211_X1 g_43_39 (.ZN (n_43_39), .A (n_39_41), .B (n_40_41), .C1 (n_36_43), .C2 (n_33_43) );
AOI211_X1 g_45_38 (.ZN (n_45_38), .A (n_41_40), .B (n_39_43), .C1 (n_38_42), .C2 (n_32_45) );
AOI211_X1 g_47_37 (.ZN (n_47_37), .A (n_43_39), .B (n_37_42), .C1 (n_40_41), .C2 (n_34_44) );
AOI211_X1 g_49_36 (.ZN (n_49_36), .A (n_45_38), .B (n_39_41), .C1 (n_39_43), .C2 (n_36_43) );
AOI211_X1 g_51_35 (.ZN (n_51_35), .A (n_47_37), .B (n_41_40), .C1 (n_37_42), .C2 (n_38_42) );
AOI211_X1 g_53_34 (.ZN (n_53_34), .A (n_49_36), .B (n_43_39), .C1 (n_39_41), .C2 (n_40_41) );
AOI211_X1 g_55_33 (.ZN (n_55_33), .A (n_51_35), .B (n_45_38), .C1 (n_41_40), .C2 (n_39_43) );
AOI211_X1 g_57_32 (.ZN (n_57_32), .A (n_53_34), .B (n_47_37), .C1 (n_43_39), .C2 (n_37_42) );
AOI211_X1 g_59_31 (.ZN (n_59_31), .A (n_55_33), .B (n_49_36), .C1 (n_45_38), .C2 (n_39_41) );
AOI211_X1 g_61_30 (.ZN (n_61_30), .A (n_57_32), .B (n_51_35), .C1 (n_47_37), .C2 (n_41_40) );
AOI211_X1 g_63_29 (.ZN (n_63_29), .A (n_59_31), .B (n_53_34), .C1 (n_49_36), .C2 (n_43_39) );
AOI211_X1 g_65_28 (.ZN (n_65_28), .A (n_61_30), .B (n_55_33), .C1 (n_51_35), .C2 (n_45_38) );
AOI211_X1 g_67_27 (.ZN (n_67_27), .A (n_63_29), .B (n_57_32), .C1 (n_53_34), .C2 (n_47_37) );
AOI211_X1 g_66_29 (.ZN (n_66_29), .A (n_65_28), .B (n_59_31), .C1 (n_55_33), .C2 (n_49_36) );
AOI211_X1 g_68_28 (.ZN (n_68_28), .A (n_67_27), .B (n_61_30), .C1 (n_57_32), .C2 (n_51_35) );
AOI211_X1 g_70_27 (.ZN (n_70_27), .A (n_66_29), .B (n_63_29), .C1 (n_59_31), .C2 (n_53_34) );
AOI211_X1 g_69_29 (.ZN (n_69_29), .A (n_68_28), .B (n_65_28), .C1 (n_61_30), .C2 (n_55_33) );
AOI211_X1 g_68_27 (.ZN (n_68_27), .A (n_70_27), .B (n_67_27), .C1 (n_63_29), .C2 (n_57_32) );
AOI211_X1 g_70_26 (.ZN (n_70_26), .A (n_69_29), .B (n_66_29), .C1 (n_65_28), .C2 (n_59_31) );
AOI211_X1 g_69_28 (.ZN (n_69_28), .A (n_68_27), .B (n_68_28), .C1 (n_67_27), .C2 (n_61_30) );
AOI211_X1 g_71_27 (.ZN (n_71_27), .A (n_70_26), .B (n_70_27), .C1 (n_66_29), .C2 (n_63_29) );
AOI211_X1 g_73_26 (.ZN (n_73_26), .A (n_69_28), .B (n_69_29), .C1 (n_68_28), .C2 (n_65_28) );
AOI211_X1 g_75_25 (.ZN (n_75_25), .A (n_71_27), .B (n_68_27), .C1 (n_70_27), .C2 (n_67_27) );
AOI211_X1 g_77_24 (.ZN (n_77_24), .A (n_73_26), .B (n_70_26), .C1 (n_69_29), .C2 (n_66_29) );
AOI211_X1 g_79_23 (.ZN (n_79_23), .A (n_75_25), .B (n_69_28), .C1 (n_68_27), .C2 (n_68_28) );
AOI211_X1 g_81_22 (.ZN (n_81_22), .A (n_77_24), .B (n_71_27), .C1 (n_70_26), .C2 (n_70_27) );
AOI211_X1 g_83_21 (.ZN (n_83_21), .A (n_79_23), .B (n_73_26), .C1 (n_69_28), .C2 (n_69_29) );
AOI211_X1 g_85_20 (.ZN (n_85_20), .A (n_81_22), .B (n_75_25), .C1 (n_71_27), .C2 (n_68_27) );
AOI211_X1 g_87_19 (.ZN (n_87_19), .A (n_83_21), .B (n_77_24), .C1 (n_73_26), .C2 (n_70_26) );
AOI211_X1 g_89_18 (.ZN (n_89_18), .A (n_85_20), .B (n_79_23), .C1 (n_75_25), .C2 (n_69_28) );
AOI211_X1 g_88_20 (.ZN (n_88_20), .A (n_87_19), .B (n_81_22), .C1 (n_77_24), .C2 (n_71_27) );
AOI211_X1 g_90_19 (.ZN (n_90_19), .A (n_89_18), .B (n_83_21), .C1 (n_79_23), .C2 (n_73_26) );
AOI211_X1 g_92_18 (.ZN (n_92_18), .A (n_88_20), .B (n_85_20), .C1 (n_81_22), .C2 (n_75_25) );
AOI211_X1 g_93_16 (.ZN (n_93_16), .A (n_90_19), .B (n_87_19), .C1 (n_83_21), .C2 (n_77_24) );
AOI211_X1 g_95_15 (.ZN (n_95_15), .A (n_92_18), .B (n_89_18), .C1 (n_85_20), .C2 (n_79_23) );
AOI211_X1 g_97_14 (.ZN (n_97_14), .A (n_93_16), .B (n_88_20), .C1 (n_87_19), .C2 (n_81_22) );
AOI211_X1 g_99_15 (.ZN (n_99_15), .A (n_95_15), .B (n_90_19), .C1 (n_89_18), .C2 (n_83_21) );
AOI211_X1 g_100_17 (.ZN (n_100_17), .A (n_97_14), .B (n_92_18), .C1 (n_88_20), .C2 (n_85_20) );
AOI211_X1 g_98_16 (.ZN (n_98_16), .A (n_99_15), .B (n_93_16), .C1 (n_90_19), .C2 (n_87_19) );
AOI211_X1 g_96_15 (.ZN (n_96_15), .A (n_100_17), .B (n_95_15), .C1 (n_92_18), .C2 (n_89_18) );
AOI211_X1 g_94_16 (.ZN (n_94_16), .A (n_98_16), .B (n_97_14), .C1 (n_93_16), .C2 (n_88_20) );
AOI211_X1 g_92_17 (.ZN (n_92_17), .A (n_96_15), .B (n_99_15), .C1 (n_95_15), .C2 (n_90_19) );
AOI211_X1 g_90_18 (.ZN (n_90_18), .A (n_94_16), .B (n_100_17), .C1 (n_97_14), .C2 (n_92_18) );
AOI211_X1 g_88_19 (.ZN (n_88_19), .A (n_92_17), .B (n_98_16), .C1 (n_99_15), .C2 (n_93_16) );
AOI211_X1 g_86_20 (.ZN (n_86_20), .A (n_90_18), .B (n_96_15), .C1 (n_100_17), .C2 (n_95_15) );
AOI211_X1 g_84_21 (.ZN (n_84_21), .A (n_88_19), .B (n_94_16), .C1 (n_98_16), .C2 (n_97_14) );
AOI211_X1 g_82_22 (.ZN (n_82_22), .A (n_86_20), .B (n_92_17), .C1 (n_96_15), .C2 (n_99_15) );
AOI211_X1 g_80_23 (.ZN (n_80_23), .A (n_84_21), .B (n_90_18), .C1 (n_94_16), .C2 (n_100_17) );
AOI211_X1 g_78_24 (.ZN (n_78_24), .A (n_82_22), .B (n_88_19), .C1 (n_92_17), .C2 (n_98_16) );
AOI211_X1 g_76_25 (.ZN (n_76_25), .A (n_80_23), .B (n_86_20), .C1 (n_90_18), .C2 (n_96_15) );
AOI211_X1 g_77_23 (.ZN (n_77_23), .A (n_78_24), .B (n_84_21), .C1 (n_88_19), .C2 (n_94_16) );
AOI211_X1 g_75_24 (.ZN (n_75_24), .A (n_76_25), .B (n_82_22), .C1 (n_86_20), .C2 (n_92_17) );
AOI211_X1 g_73_25 (.ZN (n_73_25), .A (n_77_23), .B (n_80_23), .C1 (n_84_21), .C2 (n_90_18) );
AOI211_X1 g_71_26 (.ZN (n_71_26), .A (n_75_24), .B (n_78_24), .C1 (n_82_22), .C2 (n_88_19) );
AOI211_X1 g_69_27 (.ZN (n_69_27), .A (n_73_25), .B (n_76_25), .C1 (n_80_23), .C2 (n_86_20) );
AOI211_X1 g_67_28 (.ZN (n_67_28), .A (n_71_26), .B (n_77_23), .C1 (n_78_24), .C2 (n_84_21) );
AOI211_X1 g_65_29 (.ZN (n_65_29), .A (n_69_27), .B (n_75_24), .C1 (n_76_25), .C2 (n_82_22) );
AOI211_X1 g_63_30 (.ZN (n_63_30), .A (n_67_28), .B (n_73_25), .C1 (n_77_23), .C2 (n_80_23) );
AOI211_X1 g_61_31 (.ZN (n_61_31), .A (n_65_29), .B (n_71_26), .C1 (n_75_24), .C2 (n_78_24) );
AOI211_X1 g_59_32 (.ZN (n_59_32), .A (n_63_30), .B (n_69_27), .C1 (n_73_25), .C2 (n_76_25) );
AOI211_X1 g_57_33 (.ZN (n_57_33), .A (n_61_31), .B (n_67_28), .C1 (n_71_26), .C2 (n_77_23) );
AOI211_X1 g_55_34 (.ZN (n_55_34), .A (n_59_32), .B (n_65_29), .C1 (n_69_27), .C2 (n_75_24) );
AOI211_X1 g_53_35 (.ZN (n_53_35), .A (n_57_33), .B (n_63_30), .C1 (n_67_28), .C2 (n_73_25) );
AOI211_X1 g_51_36 (.ZN (n_51_36), .A (n_55_34), .B (n_61_31), .C1 (n_65_29), .C2 (n_71_26) );
AOI211_X1 g_49_37 (.ZN (n_49_37), .A (n_53_35), .B (n_59_32), .C1 (n_63_30), .C2 (n_69_27) );
AOI211_X1 g_47_38 (.ZN (n_47_38), .A (n_51_36), .B (n_57_33), .C1 (n_61_31), .C2 (n_67_28) );
AOI211_X1 g_45_39 (.ZN (n_45_39), .A (n_49_37), .B (n_55_34), .C1 (n_59_32), .C2 (n_65_29) );
AOI211_X1 g_43_40 (.ZN (n_43_40), .A (n_47_38), .B (n_53_35), .C1 (n_57_33), .C2 (n_63_30) );
AOI211_X1 g_41_41 (.ZN (n_41_41), .A (n_45_39), .B (n_51_36), .C1 (n_55_34), .C2 (n_61_31) );
AOI211_X1 g_39_42 (.ZN (n_39_42), .A (n_43_40), .B (n_49_37), .C1 (n_53_35), .C2 (n_59_32) );
AOI211_X1 g_37_43 (.ZN (n_37_43), .A (n_41_41), .B (n_47_38), .C1 (n_51_36), .C2 (n_57_33) );
AOI211_X1 g_35_44 (.ZN (n_35_44), .A (n_39_42), .B (n_45_39), .C1 (n_49_37), .C2 (n_55_34) );
AOI211_X1 g_33_45 (.ZN (n_33_45), .A (n_37_43), .B (n_43_40), .C1 (n_47_38), .C2 (n_53_35) );
AOI211_X1 g_31_46 (.ZN (n_31_46), .A (n_35_44), .B (n_41_41), .C1 (n_45_39), .C2 (n_51_36) );
AOI211_X1 g_29_47 (.ZN (n_29_47), .A (n_33_45), .B (n_39_42), .C1 (n_43_40), .C2 (n_49_37) );
AOI211_X1 g_27_48 (.ZN (n_27_48), .A (n_31_46), .B (n_37_43), .C1 (n_41_41), .C2 (n_47_38) );
AOI211_X1 g_25_49 (.ZN (n_25_49), .A (n_29_47), .B (n_35_44), .C1 (n_39_42), .C2 (n_45_39) );
AOI211_X1 g_26_47 (.ZN (n_26_47), .A (n_27_48), .B (n_33_45), .C1 (n_37_43), .C2 (n_43_40) );
AOI211_X1 g_24_48 (.ZN (n_24_48), .A (n_25_49), .B (n_31_46), .C1 (n_35_44), .C2 (n_41_41) );
AOI211_X1 g_22_49 (.ZN (n_22_49), .A (n_26_47), .B (n_29_47), .C1 (n_33_45), .C2 (n_39_42) );
AOI211_X1 g_20_50 (.ZN (n_20_50), .A (n_24_48), .B (n_27_48), .C1 (n_31_46), .C2 (n_37_43) );
AOI211_X1 g_18_51 (.ZN (n_18_51), .A (n_22_49), .B (n_25_49), .C1 (n_29_47), .C2 (n_35_44) );
AOI211_X1 g_16_52 (.ZN (n_16_52), .A (n_20_50), .B (n_26_47), .C1 (n_27_48), .C2 (n_33_45) );
AOI211_X1 g_15_54 (.ZN (n_15_54), .A (n_18_51), .B (n_24_48), .C1 (n_25_49), .C2 (n_31_46) );
AOI211_X1 g_14_52 (.ZN (n_14_52), .A (n_16_52), .B (n_22_49), .C1 (n_26_47), .C2 (n_29_47) );
AOI211_X1 g_16_51 (.ZN (n_16_51), .A (n_15_54), .B (n_20_50), .C1 (n_24_48), .C2 (n_27_48) );
AOI211_X1 g_17_53 (.ZN (n_17_53), .A (n_14_52), .B (n_18_51), .C1 (n_22_49), .C2 (n_25_49) );
AOI211_X1 g_19_52 (.ZN (n_19_52), .A (n_16_51), .B (n_16_52), .C1 (n_20_50), .C2 (n_26_47) );
AOI211_X1 g_21_51 (.ZN (n_21_51), .A (n_17_53), .B (n_15_54), .C1 (n_18_51), .C2 (n_24_48) );
AOI211_X1 g_23_50 (.ZN (n_23_50), .A (n_19_52), .B (n_14_52), .C1 (n_16_52), .C2 (n_22_49) );
AOI211_X1 g_22_52 (.ZN (n_22_52), .A (n_21_51), .B (n_16_51), .C1 (n_15_54), .C2 (n_20_50) );
AOI211_X1 g_21_50 (.ZN (n_21_50), .A (n_23_50), .B (n_17_53), .C1 (n_14_52), .C2 (n_18_51) );
AOI211_X1 g_23_49 (.ZN (n_23_49), .A (n_22_52), .B (n_19_52), .C1 (n_16_51), .C2 (n_16_52) );
AOI211_X1 g_25_48 (.ZN (n_25_48), .A (n_21_50), .B (n_21_51), .C1 (n_17_53), .C2 (n_15_54) );
AOI211_X1 g_27_47 (.ZN (n_27_47), .A (n_23_49), .B (n_23_50), .C1 (n_19_52), .C2 (n_14_52) );
AOI211_X1 g_29_46 (.ZN (n_29_46), .A (n_25_48), .B (n_22_52), .C1 (n_21_51), .C2 (n_16_51) );
AOI211_X1 g_31_45 (.ZN (n_31_45), .A (n_27_47), .B (n_21_50), .C1 (n_23_50), .C2 (n_17_53) );
AOI211_X1 g_33_44 (.ZN (n_33_44), .A (n_29_46), .B (n_23_49), .C1 (n_22_52), .C2 (n_19_52) );
AOI211_X1 g_35_43 (.ZN (n_35_43), .A (n_31_45), .B (n_25_48), .C1 (n_21_50), .C2 (n_21_51) );
AOI211_X1 g_37_44 (.ZN (n_37_44), .A (n_33_44), .B (n_27_47), .C1 (n_23_49), .C2 (n_23_50) );
AOI211_X1 g_35_45 (.ZN (n_35_45), .A (n_35_43), .B (n_29_46), .C1 (n_25_48), .C2 (n_22_52) );
AOI211_X1 g_33_46 (.ZN (n_33_46), .A (n_37_44), .B (n_31_45), .C1 (n_27_47), .C2 (n_21_50) );
AOI211_X1 g_31_47 (.ZN (n_31_47), .A (n_35_45), .B (n_33_44), .C1 (n_29_46), .C2 (n_23_49) );
AOI211_X1 g_29_48 (.ZN (n_29_48), .A (n_33_46), .B (n_35_43), .C1 (n_31_45), .C2 (n_25_48) );
AOI211_X1 g_30_46 (.ZN (n_30_46), .A (n_31_47), .B (n_37_44), .C1 (n_33_44), .C2 (n_27_47) );
AOI211_X1 g_28_47 (.ZN (n_28_47), .A (n_29_48), .B (n_35_45), .C1 (n_35_43), .C2 (n_29_46) );
AOI211_X1 g_26_48 (.ZN (n_26_48), .A (n_30_46), .B (n_33_46), .C1 (n_37_44), .C2 (n_31_45) );
AOI211_X1 g_24_49 (.ZN (n_24_49), .A (n_28_47), .B (n_31_47), .C1 (n_35_45), .C2 (n_33_44) );
AOI211_X1 g_22_50 (.ZN (n_22_50), .A (n_26_48), .B (n_29_48), .C1 (n_33_46), .C2 (n_35_43) );
AOI211_X1 g_20_51 (.ZN (n_20_51), .A (n_24_49), .B (n_30_46), .C1 (n_31_47), .C2 (n_37_44) );
AOI211_X1 g_18_52 (.ZN (n_18_52), .A (n_22_50), .B (n_28_47), .C1 (n_29_48), .C2 (n_35_45) );
AOI211_X1 g_16_53 (.ZN (n_16_53), .A (n_20_51), .B (n_26_48), .C1 (n_30_46), .C2 (n_33_46) );
AOI211_X1 g_14_54 (.ZN (n_14_54), .A (n_18_52), .B (n_24_49), .C1 (n_28_47), .C2 (n_31_47) );
AOI211_X1 g_12_53 (.ZN (n_12_53), .A (n_16_53), .B (n_22_50), .C1 (n_26_48), .C2 (n_29_48) );
AOI211_X1 g_10_54 (.ZN (n_10_54), .A (n_14_54), .B (n_20_51), .C1 (n_24_49), .C2 (n_30_46) );
AOI211_X1 g_12_55 (.ZN (n_12_55), .A (n_12_53), .B (n_18_52), .C1 (n_22_50), .C2 (n_28_47) );
AOI211_X1 g_10_56 (.ZN (n_10_56), .A (n_10_54), .B (n_16_53), .C1 (n_20_51), .C2 (n_26_48) );
AOI211_X1 g_8_57 (.ZN (n_8_57), .A (n_12_55), .B (n_14_54), .C1 (n_18_52), .C2 (n_24_49) );
AOI211_X1 g_7_59 (.ZN (n_7_59), .A (n_10_56), .B (n_12_53), .C1 (n_16_53), .C2 (n_22_50) );
AOI211_X1 g_6_57 (.ZN (n_6_57), .A (n_8_57), .B (n_10_54), .C1 (n_14_54), .C2 (n_20_51) );
AOI211_X1 g_4_58 (.ZN (n_4_58), .A (n_7_59), .B (n_12_55), .C1 (n_12_53), .C2 (n_18_52) );
AOI211_X1 g_5_60 (.ZN (n_5_60), .A (n_6_57), .B (n_10_56), .C1 (n_10_54), .C2 (n_16_53) );
AOI211_X1 g_4_62 (.ZN (n_4_62), .A (n_4_58), .B (n_8_57), .C1 (n_12_55), .C2 (n_14_54) );
AOI211_X1 g_3_60 (.ZN (n_3_60), .A (n_5_60), .B (n_7_59), .C1 (n_10_56), .C2 (n_12_53) );
AOI211_X1 g_2_62 (.ZN (n_2_62), .A (n_4_62), .B (n_6_57), .C1 (n_8_57), .C2 (n_10_54) );
AOI211_X1 g_4_61 (.ZN (n_4_61), .A (n_3_60), .B (n_4_58), .C1 (n_7_59), .C2 (n_12_55) );
AOI211_X1 g_5_59 (.ZN (n_5_59), .A (n_2_62), .B (n_5_60), .C1 (n_6_57), .C2 (n_10_56) );
AOI211_X1 g_6_61 (.ZN (n_6_61), .A (n_4_61), .B (n_4_62), .C1 (n_4_58), .C2 (n_8_57) );
AOI211_X1 g_5_63 (.ZN (n_5_63), .A (n_5_59), .B (n_3_60), .C1 (n_5_60), .C2 (n_7_59) );
AOI211_X1 g_3_64 (.ZN (n_3_64), .A (n_6_61), .B (n_2_62), .C1 (n_4_62), .C2 (n_6_57) );
AOI211_X1 g_2_66 (.ZN (n_2_66), .A (n_5_63), .B (n_4_61), .C1 (n_3_60), .C2 (n_4_58) );
AOI211_X1 g_4_65 (.ZN (n_4_65), .A (n_3_64), .B (n_5_59), .C1 (n_2_62), .C2 (n_5_60) );
AOI211_X1 g_6_64 (.ZN (n_6_64), .A (n_2_66), .B (n_6_61), .C1 (n_4_61), .C2 (n_4_62) );
AOI211_X1 g_4_63 (.ZN (n_4_63), .A (n_4_65), .B (n_5_63), .C1 (n_5_59), .C2 (n_3_60) );
AOI211_X1 g_5_61 (.ZN (n_5_61), .A (n_6_64), .B (n_3_64), .C1 (n_6_61), .C2 (n_2_62) );
AOI211_X1 g_6_59 (.ZN (n_6_59), .A (n_4_63), .B (n_2_66), .C1 (n_5_63), .C2 (n_4_61) );
AOI211_X1 g_7_57 (.ZN (n_7_57), .A (n_5_61), .B (n_4_65), .C1 (n_3_64), .C2 (n_5_59) );
AOI211_X1 g_9_56 (.ZN (n_9_56), .A (n_6_59), .B (n_6_64), .C1 (n_2_66), .C2 (n_6_61) );
AOI211_X1 g_11_55 (.ZN (n_11_55), .A (n_7_57), .B (n_4_63), .C1 (n_4_65), .C2 (n_5_63) );
AOI211_X1 g_13_54 (.ZN (n_13_54), .A (n_9_56), .B (n_5_61), .C1 (n_6_64), .C2 (n_3_64) );
AOI211_X1 g_15_53 (.ZN (n_15_53), .A (n_11_55), .B (n_6_59), .C1 (n_4_63), .C2 (n_2_66) );
AOI211_X1 g_17_52 (.ZN (n_17_52), .A (n_13_54), .B (n_7_57), .C1 (n_5_61), .C2 (n_4_65) );
AOI211_X1 g_19_51 (.ZN (n_19_51), .A (n_15_53), .B (n_9_56), .C1 (n_6_59), .C2 (n_6_64) );
AOI211_X1 g_20_53 (.ZN (n_20_53), .A (n_17_52), .B (n_11_55), .C1 (n_7_57), .C2 (n_4_63) );
AOI211_X1 g_18_54 (.ZN (n_18_54), .A (n_19_51), .B (n_13_54), .C1 (n_9_56), .C2 (n_5_61) );
AOI211_X1 g_16_55 (.ZN (n_16_55), .A (n_20_53), .B (n_15_53), .C1 (n_11_55), .C2 (n_6_59) );
AOI211_X1 g_14_56 (.ZN (n_14_56), .A (n_18_54), .B (n_17_52), .C1 (n_13_54), .C2 (n_7_57) );
AOI211_X1 g_12_57 (.ZN (n_12_57), .A (n_16_55), .B (n_19_51), .C1 (n_15_53), .C2 (n_9_56) );
AOI211_X1 g_13_55 (.ZN (n_13_55), .A (n_14_56), .B (n_20_53), .C1 (n_17_52), .C2 (n_11_55) );
AOI211_X1 g_11_56 (.ZN (n_11_56), .A (n_12_57), .B (n_18_54), .C1 (n_19_51), .C2 (n_13_54) );
AOI211_X1 g_12_54 (.ZN (n_12_54), .A (n_13_55), .B (n_16_55), .C1 (n_20_53), .C2 (n_15_53) );
AOI211_X1 g_10_55 (.ZN (n_10_55), .A (n_11_56), .B (n_14_56), .C1 (n_18_54), .C2 (n_17_52) );
AOI211_X1 g_8_56 (.ZN (n_8_56), .A (n_12_54), .B (n_12_57), .C1 (n_16_55), .C2 (n_19_51) );
AOI211_X1 g_7_58 (.ZN (n_7_58), .A (n_10_55), .B (n_13_55), .C1 (n_14_56), .C2 (n_20_53) );
AOI211_X1 g_9_57 (.ZN (n_9_57), .A (n_8_56), .B (n_11_56), .C1 (n_12_57), .C2 (n_18_54) );
AOI211_X1 g_8_59 (.ZN (n_8_59), .A (n_7_58), .B (n_12_54), .C1 (n_13_55), .C2 (n_16_55) );
AOI211_X1 g_6_60 (.ZN (n_6_60), .A (n_9_57), .B (n_10_55), .C1 (n_11_56), .C2 (n_14_56) );
AOI211_X1 g_7_62 (.ZN (n_7_62), .A (n_8_59), .B (n_8_56), .C1 (n_12_54), .C2 (n_12_57) );
AOI211_X1 g_8_60 (.ZN (n_8_60), .A (n_6_60), .B (n_7_58), .C1 (n_10_55), .C2 (n_13_55) );
AOI211_X1 g_9_58 (.ZN (n_9_58), .A (n_7_62), .B (n_9_57), .C1 (n_8_56), .C2 (n_11_56) );
AOI211_X1 g_11_57 (.ZN (n_11_57), .A (n_8_60), .B (n_8_59), .C1 (n_7_58), .C2 (n_12_54) );
AOI211_X1 g_13_56 (.ZN (n_13_56), .A (n_9_58), .B (n_6_60), .C1 (n_9_57), .C2 (n_10_55) );
AOI211_X1 g_15_55 (.ZN (n_15_55), .A (n_11_57), .B (n_7_62), .C1 (n_8_59), .C2 (n_8_56) );
AOI211_X1 g_17_54 (.ZN (n_17_54), .A (n_13_56), .B (n_8_60), .C1 (n_6_60), .C2 (n_7_58) );
AOI211_X1 g_19_53 (.ZN (n_19_53), .A (n_15_55), .B (n_9_58), .C1 (n_7_62), .C2 (n_9_57) );
AOI211_X1 g_21_52 (.ZN (n_21_52), .A (n_17_54), .B (n_11_57), .C1 (n_8_60), .C2 (n_8_59) );
AOI211_X1 g_23_51 (.ZN (n_23_51), .A (n_19_53), .B (n_13_56), .C1 (n_9_58), .C2 (n_6_60) );
AOI211_X1 g_25_50 (.ZN (n_25_50), .A (n_21_52), .B (n_15_55), .C1 (n_11_57), .C2 (n_7_62) );
AOI211_X1 g_27_49 (.ZN (n_27_49), .A (n_23_51), .B (n_17_54), .C1 (n_13_56), .C2 (n_8_60) );
AOI211_X1 g_26_51 (.ZN (n_26_51), .A (n_25_50), .B (n_19_53), .C1 (n_15_55), .C2 (n_9_58) );
AOI211_X1 g_24_50 (.ZN (n_24_50), .A (n_27_49), .B (n_21_52), .C1 (n_17_54), .C2 (n_11_57) );
AOI211_X1 g_26_49 (.ZN (n_26_49), .A (n_26_51), .B (n_23_51), .C1 (n_19_53), .C2 (n_13_56) );
AOI211_X1 g_28_48 (.ZN (n_28_48), .A (n_24_50), .B (n_25_50), .C1 (n_21_52), .C2 (n_15_55) );
AOI211_X1 g_30_47 (.ZN (n_30_47), .A (n_26_49), .B (n_27_49), .C1 (n_23_51), .C2 (n_17_54) );
AOI211_X1 g_32_46 (.ZN (n_32_46), .A (n_28_48), .B (n_26_51), .C1 (n_25_50), .C2 (n_19_53) );
AOI211_X1 g_34_45 (.ZN (n_34_45), .A (n_30_47), .B (n_24_50), .C1 (n_27_49), .C2 (n_21_52) );
AOI211_X1 g_36_44 (.ZN (n_36_44), .A (n_32_46), .B (n_26_49), .C1 (n_26_51), .C2 (n_23_51) );
AOI211_X1 g_38_43 (.ZN (n_38_43), .A (n_34_45), .B (n_28_48), .C1 (n_24_50), .C2 (n_25_50) );
AOI211_X1 g_40_42 (.ZN (n_40_42), .A (n_36_44), .B (n_30_47), .C1 (n_26_49), .C2 (n_27_49) );
AOI211_X1 g_42_41 (.ZN (n_42_41), .A (n_38_43), .B (n_32_46), .C1 (n_28_48), .C2 (n_26_51) );
AOI211_X1 g_44_40 (.ZN (n_44_40), .A (n_40_42), .B (n_34_45), .C1 (n_30_47), .C2 (n_24_50) );
AOI211_X1 g_46_39 (.ZN (n_46_39), .A (n_42_41), .B (n_36_44), .C1 (n_32_46), .C2 (n_26_49) );
AOI211_X1 g_48_38 (.ZN (n_48_38), .A (n_44_40), .B (n_38_43), .C1 (n_34_45), .C2 (n_28_48) );
AOI211_X1 g_50_37 (.ZN (n_50_37), .A (n_46_39), .B (n_40_42), .C1 (n_36_44), .C2 (n_30_47) );
AOI211_X1 g_52_36 (.ZN (n_52_36), .A (n_48_38), .B (n_42_41), .C1 (n_38_43), .C2 (n_32_46) );
AOI211_X1 g_54_35 (.ZN (n_54_35), .A (n_50_37), .B (n_44_40), .C1 (n_40_42), .C2 (n_34_45) );
AOI211_X1 g_56_34 (.ZN (n_56_34), .A (n_52_36), .B (n_46_39), .C1 (n_42_41), .C2 (n_36_44) );
AOI211_X1 g_58_33 (.ZN (n_58_33), .A (n_54_35), .B (n_48_38), .C1 (n_44_40), .C2 (n_38_43) );
AOI211_X1 g_60_32 (.ZN (n_60_32), .A (n_56_34), .B (n_50_37), .C1 (n_46_39), .C2 (n_40_42) );
AOI211_X1 g_62_31 (.ZN (n_62_31), .A (n_58_33), .B (n_52_36), .C1 (n_48_38), .C2 (n_42_41) );
AOI211_X1 g_64_30 (.ZN (n_64_30), .A (n_60_32), .B (n_54_35), .C1 (n_50_37), .C2 (n_44_40) );
AOI211_X1 g_63_32 (.ZN (n_63_32), .A (n_62_31), .B (n_56_34), .C1 (n_52_36), .C2 (n_46_39) );
AOI211_X1 g_62_30 (.ZN (n_62_30), .A (n_64_30), .B (n_58_33), .C1 (n_54_35), .C2 (n_48_38) );
AOI211_X1 g_64_29 (.ZN (n_64_29), .A (n_63_32), .B (n_60_32), .C1 (n_56_34), .C2 (n_50_37) );
AOI211_X1 g_66_28 (.ZN (n_66_28), .A (n_62_30), .B (n_62_31), .C1 (n_58_33), .C2 (n_52_36) );
AOI211_X1 g_67_30 (.ZN (n_67_30), .A (n_64_29), .B (n_64_30), .C1 (n_60_32), .C2 (n_54_35) );
AOI211_X1 g_65_31 (.ZN (n_65_31), .A (n_66_28), .B (n_63_32), .C1 (n_62_31), .C2 (n_56_34) );
AOI211_X1 g_64_33 (.ZN (n_64_33), .A (n_67_30), .B (n_62_30), .C1 (n_64_30), .C2 (n_58_33) );
AOI211_X1 g_63_31 (.ZN (n_63_31), .A (n_65_31), .B (n_64_29), .C1 (n_63_32), .C2 (n_60_32) );
AOI211_X1 g_65_30 (.ZN (n_65_30), .A (n_64_33), .B (n_66_28), .C1 (n_62_30), .C2 (n_62_31) );
AOI211_X1 g_67_29 (.ZN (n_67_29), .A (n_63_31), .B (n_67_30), .C1 (n_64_29), .C2 (n_64_30) );
AOI211_X1 g_66_31 (.ZN (n_66_31), .A (n_65_30), .B (n_65_31), .C1 (n_66_28), .C2 (n_63_32) );
AOI211_X1 g_68_30 (.ZN (n_68_30), .A (n_67_29), .B (n_64_33), .C1 (n_67_30), .C2 (n_62_30) );
AOI211_X1 g_70_29 (.ZN (n_70_29), .A (n_66_31), .B (n_63_31), .C1 (n_65_31), .C2 (n_64_29) );
AOI211_X1 g_72_28 (.ZN (n_72_28), .A (n_68_30), .B (n_65_30), .C1 (n_64_33), .C2 (n_66_28) );
AOI211_X1 g_74_27 (.ZN (n_74_27), .A (n_70_29), .B (n_67_29), .C1 (n_63_31), .C2 (n_67_30) );
AOI211_X1 g_76_26 (.ZN (n_76_26), .A (n_72_28), .B (n_66_31), .C1 (n_65_30), .C2 (n_65_31) );
AOI211_X1 g_78_25 (.ZN (n_78_25), .A (n_74_27), .B (n_68_30), .C1 (n_67_29), .C2 (n_64_33) );
AOI211_X1 g_80_24 (.ZN (n_80_24), .A (n_76_26), .B (n_70_29), .C1 (n_66_31), .C2 (n_63_31) );
AOI211_X1 g_82_23 (.ZN (n_82_23), .A (n_78_25), .B (n_72_28), .C1 (n_68_30), .C2 (n_65_30) );
AOI211_X1 g_84_22 (.ZN (n_84_22), .A (n_80_24), .B (n_74_27), .C1 (n_70_29), .C2 (n_67_29) );
AOI211_X1 g_86_21 (.ZN (n_86_21), .A (n_82_23), .B (n_76_26), .C1 (n_72_28), .C2 (n_66_31) );
AOI211_X1 g_85_23 (.ZN (n_85_23), .A (n_84_22), .B (n_78_25), .C1 (n_74_27), .C2 (n_68_30) );
AOI211_X1 g_87_22 (.ZN (n_87_22), .A (n_86_21), .B (n_80_24), .C1 (n_76_26), .C2 (n_70_29) );
AOI211_X1 g_89_21 (.ZN (n_89_21), .A (n_85_23), .B (n_82_23), .C1 (n_78_25), .C2 (n_72_28) );
AOI211_X1 g_91_20 (.ZN (n_91_20), .A (n_87_22), .B (n_84_22), .C1 (n_80_24), .C2 (n_74_27) );
AOI211_X1 g_93_19 (.ZN (n_93_19), .A (n_89_21), .B (n_86_21), .C1 (n_82_23), .C2 (n_76_26) );
AOI211_X1 g_94_17 (.ZN (n_94_17), .A (n_91_20), .B (n_85_23), .C1 (n_84_22), .C2 (n_78_25) );
AOI211_X1 g_96_16 (.ZN (n_96_16), .A (n_93_19), .B (n_87_22), .C1 (n_86_21), .C2 (n_80_24) );
AOI211_X1 g_98_15 (.ZN (n_98_15), .A (n_94_17), .B (n_89_21), .C1 (n_85_23), .C2 (n_82_23) );
AOI211_X1 g_100_16 (.ZN (n_100_16), .A (n_96_16), .B (n_91_20), .C1 (n_87_22), .C2 (n_84_22) );
AOI211_X1 g_98_17 (.ZN (n_98_17), .A (n_98_15), .B (n_93_19), .C1 (n_89_21), .C2 (n_86_21) );
AOI211_X1 g_99_19 (.ZN (n_99_19), .A (n_100_16), .B (n_94_17), .C1 (n_91_20), .C2 (n_85_23) );
AOI211_X1 g_100_21 (.ZN (n_100_21), .A (n_98_17), .B (n_96_16), .C1 (n_93_19), .C2 (n_87_22) );
AOI211_X1 g_98_22 (.ZN (n_98_22), .A (n_99_19), .B (n_98_15), .C1 (n_94_17), .C2 (n_89_21) );
AOI211_X1 g_100_23 (.ZN (n_100_23), .A (n_100_21), .B (n_100_16), .C1 (n_96_16), .C2 (n_91_20) );
AOI211_X1 g_99_21 (.ZN (n_99_21), .A (n_98_22), .B (n_98_17), .C1 (n_98_15), .C2 (n_93_19) );
AOI211_X1 g_100_19 (.ZN (n_100_19), .A (n_100_23), .B (n_99_19), .C1 (n_100_16), .C2 (n_94_17) );
AOI211_X1 g_99_17 (.ZN (n_99_17), .A (n_99_21), .B (n_100_21), .C1 (n_98_17), .C2 (n_96_16) );
AOI211_X1 g_97_16 (.ZN (n_97_16), .A (n_100_19), .B (n_98_22), .C1 (n_99_19), .C2 (n_98_15) );
AOI211_X1 g_98_18 (.ZN (n_98_18), .A (n_99_17), .B (n_100_23), .C1 (n_100_21), .C2 (n_100_16) );
AOI211_X1 g_96_17 (.ZN (n_96_17), .A (n_97_16), .B (n_99_21), .C1 (n_98_22), .C2 (n_98_17) );
AOI211_X1 g_94_18 (.ZN (n_94_18), .A (n_98_18), .B (n_100_19), .C1 (n_100_23), .C2 (n_99_19) );
AOI211_X1 g_92_19 (.ZN (n_92_19), .A (n_96_17), .B (n_99_17), .C1 (n_99_21), .C2 (n_100_21) );
AOI211_X1 g_90_20 (.ZN (n_90_20), .A (n_94_18), .B (n_97_16), .C1 (n_100_19), .C2 (n_98_22) );
AOI211_X1 g_88_21 (.ZN (n_88_21), .A (n_92_19), .B (n_98_18), .C1 (n_99_17), .C2 (n_100_23) );
AOI211_X1 g_86_22 (.ZN (n_86_22), .A (n_90_20), .B (n_96_17), .C1 (n_97_16), .C2 (n_99_21) );
AOI211_X1 g_84_23 (.ZN (n_84_23), .A (n_88_21), .B (n_94_18), .C1 (n_98_18), .C2 (n_100_19) );
AOI211_X1 g_82_24 (.ZN (n_82_24), .A (n_86_22), .B (n_92_19), .C1 (n_96_17), .C2 (n_99_17) );
AOI211_X1 g_80_25 (.ZN (n_80_25), .A (n_84_23), .B (n_90_20), .C1 (n_94_18), .C2 (n_97_16) );
AOI211_X1 g_78_26 (.ZN (n_78_26), .A (n_82_24), .B (n_88_21), .C1 (n_92_19), .C2 (n_98_18) );
AOI211_X1 g_79_24 (.ZN (n_79_24), .A (n_80_25), .B (n_86_22), .C1 (n_90_20), .C2 (n_96_17) );
AOI211_X1 g_77_25 (.ZN (n_77_25), .A (n_78_26), .B (n_84_23), .C1 (n_88_21), .C2 (n_94_18) );
AOI211_X1 g_75_26 (.ZN (n_75_26), .A (n_79_24), .B (n_82_24), .C1 (n_86_22), .C2 (n_92_19) );
AOI211_X1 g_73_27 (.ZN (n_73_27), .A (n_77_25), .B (n_80_25), .C1 (n_84_23), .C2 (n_90_20) );
AOI211_X1 g_71_28 (.ZN (n_71_28), .A (n_75_26), .B (n_78_26), .C1 (n_82_24), .C2 (n_88_21) );
AOI211_X1 g_70_30 (.ZN (n_70_30), .A (n_73_27), .B (n_79_24), .C1 (n_80_25), .C2 (n_86_22) );
AOI211_X1 g_68_29 (.ZN (n_68_29), .A (n_71_28), .B (n_77_25), .C1 (n_78_26), .C2 (n_84_23) );
AOI211_X1 g_70_28 (.ZN (n_70_28), .A (n_70_30), .B (n_75_26), .C1 (n_79_24), .C2 (n_82_24) );
AOI211_X1 g_72_27 (.ZN (n_72_27), .A (n_68_29), .B (n_73_27), .C1 (n_77_25), .C2 (n_80_25) );
AOI211_X1 g_74_26 (.ZN (n_74_26), .A (n_70_28), .B (n_71_28), .C1 (n_75_26), .C2 (n_78_26) );
AOI211_X1 g_76_27 (.ZN (n_76_27), .A (n_72_27), .B (n_70_30), .C1 (n_73_27), .C2 (n_79_24) );
AOI211_X1 g_74_28 (.ZN (n_74_28), .A (n_74_26), .B (n_68_29), .C1 (n_71_28), .C2 (n_77_25) );
AOI211_X1 g_72_29 (.ZN (n_72_29), .A (n_76_27), .B (n_70_28), .C1 (n_70_30), .C2 (n_75_26) );
AOI211_X1 g_71_31 (.ZN (n_71_31), .A (n_74_28), .B (n_72_27), .C1 (n_68_29), .C2 (n_73_27) );
AOI211_X1 g_69_30 (.ZN (n_69_30), .A (n_72_29), .B (n_74_26), .C1 (n_70_28), .C2 (n_71_28) );
AOI211_X1 g_71_29 (.ZN (n_71_29), .A (n_71_31), .B (n_76_27), .C1 (n_72_27), .C2 (n_70_30) );
AOI211_X1 g_73_28 (.ZN (n_73_28), .A (n_69_30), .B (n_74_28), .C1 (n_74_26), .C2 (n_68_29) );
AOI211_X1 g_75_27 (.ZN (n_75_27), .A (n_71_29), .B (n_72_29), .C1 (n_76_27), .C2 (n_70_28) );
AOI211_X1 g_77_26 (.ZN (n_77_26), .A (n_73_28), .B (n_71_31), .C1 (n_74_28), .C2 (n_72_27) );
AOI211_X1 g_79_25 (.ZN (n_79_25), .A (n_75_27), .B (n_69_30), .C1 (n_72_29), .C2 (n_74_26) );
AOI211_X1 g_81_24 (.ZN (n_81_24), .A (n_77_26), .B (n_71_29), .C1 (n_71_31), .C2 (n_76_27) );
AOI211_X1 g_83_23 (.ZN (n_83_23), .A (n_79_25), .B (n_73_28), .C1 (n_69_30), .C2 (n_74_28) );
AOI211_X1 g_85_22 (.ZN (n_85_22), .A (n_81_24), .B (n_75_27), .C1 (n_71_29), .C2 (n_72_29) );
AOI211_X1 g_87_21 (.ZN (n_87_21), .A (n_83_23), .B (n_77_26), .C1 (n_73_28), .C2 (n_71_31) );
AOI211_X1 g_89_20 (.ZN (n_89_20), .A (n_85_22), .B (n_79_25), .C1 (n_75_27), .C2 (n_69_30) );
AOI211_X1 g_91_19 (.ZN (n_91_19), .A (n_87_21), .B (n_81_24), .C1 (n_77_26), .C2 (n_71_29) );
AOI211_X1 g_93_18 (.ZN (n_93_18), .A (n_89_20), .B (n_83_23), .C1 (n_79_25), .C2 (n_73_28) );
AOI211_X1 g_95_17 (.ZN (n_95_17), .A (n_91_19), .B (n_85_22), .C1 (n_81_24), .C2 (n_75_27) );
AOI211_X1 g_97_18 (.ZN (n_97_18), .A (n_93_18), .B (n_87_21), .C1 (n_83_23), .C2 (n_77_26) );
AOI211_X1 g_95_19 (.ZN (n_95_19), .A (n_95_17), .B (n_89_20), .C1 (n_85_22), .C2 (n_79_25) );
AOI211_X1 g_97_20 (.ZN (n_97_20), .A (n_97_18), .B (n_91_19), .C1 (n_87_21), .C2 (n_81_24) );
AOI211_X1 g_96_18 (.ZN (n_96_18), .A (n_95_19), .B (n_93_18), .C1 (n_89_20), .C2 (n_83_23) );
AOI211_X1 g_94_19 (.ZN (n_94_19), .A (n_97_20), .B (n_95_17), .C1 (n_91_19), .C2 (n_85_22) );
AOI211_X1 g_92_20 (.ZN (n_92_20), .A (n_96_18), .B (n_97_18), .C1 (n_93_18), .C2 (n_87_21) );
AOI211_X1 g_90_21 (.ZN (n_90_21), .A (n_94_19), .B (n_95_19), .C1 (n_95_17), .C2 (n_89_20) );
AOI211_X1 g_88_22 (.ZN (n_88_22), .A (n_92_20), .B (n_97_20), .C1 (n_97_18), .C2 (n_91_19) );
AOI211_X1 g_86_23 (.ZN (n_86_23), .A (n_90_21), .B (n_96_18), .C1 (n_95_19), .C2 (n_93_18) );
AOI211_X1 g_84_24 (.ZN (n_84_24), .A (n_88_22), .B (n_94_19), .C1 (n_97_20), .C2 (n_95_17) );
AOI211_X1 g_82_25 (.ZN (n_82_25), .A (n_86_23), .B (n_92_20), .C1 (n_96_18), .C2 (n_97_18) );
AOI211_X1 g_80_26 (.ZN (n_80_26), .A (n_84_24), .B (n_90_21), .C1 (n_94_19), .C2 (n_95_19) );
AOI211_X1 g_78_27 (.ZN (n_78_27), .A (n_82_25), .B (n_88_22), .C1 (n_92_20), .C2 (n_97_20) );
AOI211_X1 g_76_28 (.ZN (n_76_28), .A (n_80_26), .B (n_86_23), .C1 (n_90_21), .C2 (n_96_18) );
AOI211_X1 g_74_29 (.ZN (n_74_29), .A (n_78_27), .B (n_84_24), .C1 (n_88_22), .C2 (n_94_19) );
AOI211_X1 g_72_30 (.ZN (n_72_30), .A (n_76_28), .B (n_82_25), .C1 (n_86_23), .C2 (n_92_20) );
AOI211_X1 g_70_31 (.ZN (n_70_31), .A (n_74_29), .B (n_80_26), .C1 (n_84_24), .C2 (n_90_21) );
AOI211_X1 g_68_32 (.ZN (n_68_32), .A (n_72_30), .B (n_78_27), .C1 (n_82_25), .C2 (n_88_22) );
AOI211_X1 g_66_33 (.ZN (n_66_33), .A (n_70_31), .B (n_76_28), .C1 (n_80_26), .C2 (n_86_23) );
AOI211_X1 g_67_31 (.ZN (n_67_31), .A (n_68_32), .B (n_74_29), .C1 (n_78_27), .C2 (n_84_24) );
AOI211_X1 g_69_32 (.ZN (n_69_32), .A (n_66_33), .B (n_72_30), .C1 (n_76_28), .C2 (n_82_25) );
AOI211_X1 g_67_33 (.ZN (n_67_33), .A (n_67_31), .B (n_70_31), .C1 (n_74_29), .C2 (n_80_26) );
AOI211_X1 g_68_31 (.ZN (n_68_31), .A (n_69_32), .B (n_68_32), .C1 (n_72_30), .C2 (n_78_27) );
AOI211_X1 g_66_30 (.ZN (n_66_30), .A (n_67_33), .B (n_66_33), .C1 (n_70_31), .C2 (n_76_28) );
AOI211_X1 g_65_32 (.ZN (n_65_32), .A (n_68_31), .B (n_67_31), .C1 (n_68_32), .C2 (n_74_29) );
AOI211_X1 g_64_34 (.ZN (n_64_34), .A (n_66_30), .B (n_69_32), .C1 (n_66_33), .C2 (n_72_30) );
AOI211_X1 g_62_33 (.ZN (n_62_33), .A (n_65_32), .B (n_67_33), .C1 (n_67_31), .C2 (n_70_31) );
AOI211_X1 g_64_32 (.ZN (n_64_32), .A (n_64_34), .B (n_68_31), .C1 (n_69_32), .C2 (n_68_32) );
AOI211_X1 g_65_34 (.ZN (n_65_34), .A (n_62_33), .B (n_66_30), .C1 (n_67_33), .C2 (n_66_33) );
AOI211_X1 g_66_32 (.ZN (n_66_32), .A (n_64_32), .B (n_65_32), .C1 (n_68_31), .C2 (n_67_31) );
AOI211_X1 g_64_31 (.ZN (n_64_31), .A (n_65_34), .B (n_64_34), .C1 (n_66_30), .C2 (n_69_32) );
AOI211_X1 g_62_32 (.ZN (n_62_32), .A (n_66_32), .B (n_62_33), .C1 (n_65_32), .C2 (n_67_33) );
AOI211_X1 g_60_31 (.ZN (n_60_31), .A (n_64_31), .B (n_64_32), .C1 (n_64_34), .C2 (n_68_31) );
AOI211_X1 g_58_32 (.ZN (n_58_32), .A (n_62_32), .B (n_65_34), .C1 (n_62_33), .C2 (n_66_30) );
AOI211_X1 g_56_33 (.ZN (n_56_33), .A (n_60_31), .B (n_66_32), .C1 (n_64_32), .C2 (n_65_32) );
AOI211_X1 g_54_34 (.ZN (n_54_34), .A (n_58_32), .B (n_64_31), .C1 (n_65_34), .C2 (n_64_34) );
AOI211_X1 g_52_35 (.ZN (n_52_35), .A (n_56_33), .B (n_62_32), .C1 (n_66_32), .C2 (n_62_33) );
AOI211_X1 g_50_36 (.ZN (n_50_36), .A (n_54_34), .B (n_60_31), .C1 (n_64_31), .C2 (n_64_32) );
AOI211_X1 g_48_37 (.ZN (n_48_37), .A (n_52_35), .B (n_58_32), .C1 (n_62_32), .C2 (n_65_34) );
AOI211_X1 g_47_39 (.ZN (n_47_39), .A (n_50_36), .B (n_56_33), .C1 (n_60_31), .C2 (n_66_32) );
AOI211_X1 g_49_38 (.ZN (n_49_38), .A (n_48_37), .B (n_54_34), .C1 (n_58_32), .C2 (n_64_31) );
AOI211_X1 g_51_37 (.ZN (n_51_37), .A (n_47_39), .B (n_52_35), .C1 (n_56_33), .C2 (n_62_32) );
AOI211_X1 g_53_36 (.ZN (n_53_36), .A (n_49_38), .B (n_50_36), .C1 (n_54_34), .C2 (n_60_31) );
AOI211_X1 g_55_35 (.ZN (n_55_35), .A (n_51_37), .B (n_48_37), .C1 (n_52_35), .C2 (n_58_32) );
AOI211_X1 g_57_34 (.ZN (n_57_34), .A (n_53_36), .B (n_47_39), .C1 (n_50_36), .C2 (n_56_33) );
AOI211_X1 g_59_33 (.ZN (n_59_33), .A (n_55_35), .B (n_49_38), .C1 (n_48_37), .C2 (n_54_34) );
AOI211_X1 g_61_32 (.ZN (n_61_32), .A (n_57_34), .B (n_51_37), .C1 (n_47_39), .C2 (n_52_35) );
AOI211_X1 g_63_33 (.ZN (n_63_33), .A (n_59_33), .B (n_53_36), .C1 (n_49_38), .C2 (n_50_36) );
AOI211_X1 g_61_34 (.ZN (n_61_34), .A (n_61_32), .B (n_55_35), .C1 (n_51_37), .C2 (n_48_37) );
AOI211_X1 g_63_35 (.ZN (n_63_35), .A (n_63_33), .B (n_57_34), .C1 (n_53_36), .C2 (n_47_39) );
AOI211_X1 g_65_36 (.ZN (n_65_36), .A (n_61_34), .B (n_59_33), .C1 (n_55_35), .C2 (n_49_38) );
AOI211_X1 g_67_35 (.ZN (n_67_35), .A (n_63_35), .B (n_61_32), .C1 (n_57_34), .C2 (n_51_37) );
AOI211_X1 g_69_34 (.ZN (n_69_34), .A (n_65_36), .B (n_63_33), .C1 (n_59_33), .C2 (n_53_36) );
AOI211_X1 g_71_33 (.ZN (n_71_33), .A (n_67_35), .B (n_61_34), .C1 (n_61_32), .C2 (n_55_35) );
AOI211_X1 g_73_32 (.ZN (n_73_32), .A (n_69_34), .B (n_63_35), .C1 (n_63_33), .C2 (n_57_34) );
AOI211_X1 g_74_30 (.ZN (n_74_30), .A (n_71_33), .B (n_65_36), .C1 (n_61_34), .C2 (n_59_33) );
AOI211_X1 g_75_28 (.ZN (n_75_28), .A (n_73_32), .B (n_67_35), .C1 (n_63_35), .C2 (n_61_32) );
AOI211_X1 g_77_27 (.ZN (n_77_27), .A (n_74_30), .B (n_69_34), .C1 (n_65_36), .C2 (n_63_33) );
AOI211_X1 g_79_26 (.ZN (n_79_26), .A (n_75_28), .B (n_71_33), .C1 (n_67_35), .C2 (n_61_34) );
AOI211_X1 g_81_25 (.ZN (n_81_25), .A (n_77_27), .B (n_73_32), .C1 (n_69_34), .C2 (n_63_35) );
AOI211_X1 g_83_24 (.ZN (n_83_24), .A (n_79_26), .B (n_74_30), .C1 (n_71_33), .C2 (n_65_36) );
AOI211_X1 g_82_26 (.ZN (n_82_26), .A (n_81_25), .B (n_75_28), .C1 (n_73_32), .C2 (n_67_35) );
AOI211_X1 g_84_25 (.ZN (n_84_25), .A (n_83_24), .B (n_77_27), .C1 (n_74_30), .C2 (n_69_34) );
AOI211_X1 g_86_24 (.ZN (n_86_24), .A (n_82_26), .B (n_79_26), .C1 (n_75_28), .C2 (n_71_33) );
AOI211_X1 g_88_23 (.ZN (n_88_23), .A (n_84_25), .B (n_81_25), .C1 (n_77_27), .C2 (n_73_32) );
AOI211_X1 g_90_22 (.ZN (n_90_22), .A (n_86_24), .B (n_83_24), .C1 (n_79_26), .C2 (n_74_30) );
AOI211_X1 g_92_21 (.ZN (n_92_21), .A (n_88_23), .B (n_82_26), .C1 (n_81_25), .C2 (n_75_28) );
AOI211_X1 g_94_20 (.ZN (n_94_20), .A (n_90_22), .B (n_84_25), .C1 (n_83_24), .C2 (n_77_27) );
AOI211_X1 g_95_18 (.ZN (n_95_18), .A (n_92_21), .B (n_86_24), .C1 (n_82_26), .C2 (n_79_26) );
AOI211_X1 g_97_17 (.ZN (n_97_17), .A (n_94_20), .B (n_88_23), .C1 (n_84_25), .C2 (n_81_25) );
AOI211_X1 g_96_19 (.ZN (n_96_19), .A (n_95_18), .B (n_90_22), .C1 (n_86_24), .C2 (n_83_24) );
AOI211_X1 g_98_20 (.ZN (n_98_20), .A (n_97_17), .B (n_92_21), .C1 (n_88_23), .C2 (n_82_26) );
AOI211_X1 g_99_18 (.ZN (n_99_18), .A (n_96_19), .B (n_94_20), .C1 (n_90_22), .C2 (n_84_25) );
AOI211_X1 g_97_19 (.ZN (n_97_19), .A (n_98_20), .B (n_95_18), .C1 (n_92_21), .C2 (n_86_24) );
AOI211_X1 g_96_21 (.ZN (n_96_21), .A (n_99_18), .B (n_97_17), .C1 (n_94_20), .C2 (n_88_23) );
AOI211_X1 g_94_22 (.ZN (n_94_22), .A (n_97_19), .B (n_96_19), .C1 (n_95_18), .C2 (n_90_22) );
AOI211_X1 g_95_20 (.ZN (n_95_20), .A (n_96_21), .B (n_98_20), .C1 (n_97_17), .C2 (n_92_21) );
AOI211_X1 g_93_21 (.ZN (n_93_21), .A (n_94_22), .B (n_99_18), .C1 (n_96_19), .C2 (n_94_20) );
AOI211_X1 g_91_22 (.ZN (n_91_22), .A (n_95_20), .B (n_97_19), .C1 (n_98_20), .C2 (n_95_18) );
AOI211_X1 g_89_23 (.ZN (n_89_23), .A (n_93_21), .B (n_96_21), .C1 (n_99_18), .C2 (n_97_17) );
AOI211_X1 g_87_24 (.ZN (n_87_24), .A (n_91_22), .B (n_94_22), .C1 (n_97_19), .C2 (n_96_19) );
AOI211_X1 g_85_25 (.ZN (n_85_25), .A (n_89_23), .B (n_95_20), .C1 (n_96_21), .C2 (n_98_20) );
AOI211_X1 g_83_26 (.ZN (n_83_26), .A (n_87_24), .B (n_93_21), .C1 (n_94_22), .C2 (n_99_18) );
AOI211_X1 g_81_27 (.ZN (n_81_27), .A (n_85_25), .B (n_91_22), .C1 (n_95_20), .C2 (n_97_19) );
AOI211_X1 g_79_28 (.ZN (n_79_28), .A (n_83_26), .B (n_89_23), .C1 (n_93_21), .C2 (n_96_21) );
AOI211_X1 g_77_29 (.ZN (n_77_29), .A (n_81_27), .B (n_87_24), .C1 (n_91_22), .C2 (n_94_22) );
AOI211_X1 g_75_30 (.ZN (n_75_30), .A (n_79_28), .B (n_85_25), .C1 (n_89_23), .C2 (n_95_20) );
AOI211_X1 g_73_29 (.ZN (n_73_29), .A (n_77_29), .B (n_83_26), .C1 (n_87_24), .C2 (n_93_21) );
AOI211_X1 g_72_31 (.ZN (n_72_31), .A (n_75_30), .B (n_81_27), .C1 (n_85_25), .C2 (n_91_22) );
AOI211_X1 g_70_32 (.ZN (n_70_32), .A (n_73_29), .B (n_79_28), .C1 (n_83_26), .C2 (n_89_23) );
AOI211_X1 g_71_30 (.ZN (n_71_30), .A (n_72_31), .B (n_77_29), .C1 (n_81_27), .C2 (n_87_24) );
AOI211_X1 g_69_31 (.ZN (n_69_31), .A (n_70_32), .B (n_75_30), .C1 (n_79_28), .C2 (n_85_25) );
AOI211_X1 g_68_33 (.ZN (n_68_33), .A (n_71_30), .B (n_73_29), .C1 (n_77_29), .C2 (n_83_26) );
AOI211_X1 g_66_34 (.ZN (n_66_34), .A (n_69_31), .B (n_72_31), .C1 (n_75_30), .C2 (n_81_27) );
AOI211_X1 g_67_32 (.ZN (n_67_32), .A (n_68_33), .B (n_70_32), .C1 (n_73_29), .C2 (n_79_28) );
AOI211_X1 g_65_33 (.ZN (n_65_33), .A (n_66_34), .B (n_71_30), .C1 (n_72_31), .C2 (n_77_29) );
AOI211_X1 g_63_34 (.ZN (n_63_34), .A (n_67_32), .B (n_69_31), .C1 (n_70_32), .C2 (n_75_30) );
AOI211_X1 g_61_33 (.ZN (n_61_33), .A (n_65_33), .B (n_68_33), .C1 (n_71_30), .C2 (n_73_29) );
AOI211_X1 g_59_34 (.ZN (n_59_34), .A (n_63_34), .B (n_66_34), .C1 (n_69_31), .C2 (n_72_31) );
AOI211_X1 g_57_35 (.ZN (n_57_35), .A (n_61_33), .B (n_67_32), .C1 (n_68_33), .C2 (n_70_32) );
AOI211_X1 g_55_36 (.ZN (n_55_36), .A (n_59_34), .B (n_65_33), .C1 (n_66_34), .C2 (n_71_30) );
AOI211_X1 g_53_37 (.ZN (n_53_37), .A (n_57_35), .B (n_63_34), .C1 (n_67_32), .C2 (n_69_31) );
AOI211_X1 g_51_38 (.ZN (n_51_38), .A (n_55_36), .B (n_61_33), .C1 (n_65_33), .C2 (n_68_33) );
AOI211_X1 g_49_39 (.ZN (n_49_39), .A (n_53_37), .B (n_59_34), .C1 (n_63_34), .C2 (n_66_34) );
AOI211_X1 g_47_40 (.ZN (n_47_40), .A (n_51_38), .B (n_57_35), .C1 (n_61_33), .C2 (n_67_32) );
AOI211_X1 g_45_41 (.ZN (n_45_41), .A (n_49_39), .B (n_55_36), .C1 (n_59_34), .C2 (n_65_33) );
AOI211_X1 g_43_42 (.ZN (n_43_42), .A (n_47_40), .B (n_53_37), .C1 (n_57_35), .C2 (n_63_34) );
AOI211_X1 g_41_43 (.ZN (n_41_43), .A (n_45_41), .B (n_51_38), .C1 (n_55_36), .C2 (n_61_33) );
AOI211_X1 g_39_44 (.ZN (n_39_44), .A (n_43_42), .B (n_49_39), .C1 (n_53_37), .C2 (n_59_34) );
AOI211_X1 g_37_45 (.ZN (n_37_45), .A (n_41_43), .B (n_47_40), .C1 (n_51_38), .C2 (n_57_35) );
AOI211_X1 g_35_46 (.ZN (n_35_46), .A (n_39_44), .B (n_45_41), .C1 (n_49_39), .C2 (n_55_36) );
AOI211_X1 g_33_47 (.ZN (n_33_47), .A (n_37_45), .B (n_43_42), .C1 (n_47_40), .C2 (n_53_37) );
AOI211_X1 g_31_48 (.ZN (n_31_48), .A (n_35_46), .B (n_41_43), .C1 (n_45_41), .C2 (n_51_38) );
AOI211_X1 g_29_49 (.ZN (n_29_49), .A (n_33_47), .B (n_39_44), .C1 (n_43_42), .C2 (n_49_39) );
AOI211_X1 g_27_50 (.ZN (n_27_50), .A (n_31_48), .B (n_37_45), .C1 (n_41_43), .C2 (n_47_40) );
AOI211_X1 g_25_51 (.ZN (n_25_51), .A (n_29_49), .B (n_35_46), .C1 (n_39_44), .C2 (n_45_41) );
AOI211_X1 g_23_52 (.ZN (n_23_52), .A (n_27_50), .B (n_33_47), .C1 (n_37_45), .C2 (n_43_42) );
AOI211_X1 g_21_53 (.ZN (n_21_53), .A (n_25_51), .B (n_31_48), .C1 (n_35_46), .C2 (n_41_43) );
AOI211_X1 g_22_51 (.ZN (n_22_51), .A (n_23_52), .B (n_29_49), .C1 (n_33_47), .C2 (n_39_44) );
AOI211_X1 g_20_52 (.ZN (n_20_52), .A (n_21_53), .B (n_27_50), .C1 (n_31_48), .C2 (n_37_45) );
AOI211_X1 g_18_53 (.ZN (n_18_53), .A (n_22_51), .B (n_25_51), .C1 (n_29_49), .C2 (n_35_46) );
AOI211_X1 g_16_54 (.ZN (n_16_54), .A (n_20_52), .B (n_23_52), .C1 (n_27_50), .C2 (n_33_47) );
AOI211_X1 g_14_55 (.ZN (n_14_55), .A (n_18_53), .B (n_21_53), .C1 (n_25_51), .C2 (n_31_48) );
AOI211_X1 g_12_56 (.ZN (n_12_56), .A (n_16_54), .B (n_22_51), .C1 (n_23_52), .C2 (n_29_49) );
AOI211_X1 g_10_57 (.ZN (n_10_57), .A (n_14_55), .B (n_20_52), .C1 (n_21_53), .C2 (n_27_50) );
AOI211_X1 g_8_58 (.ZN (n_8_58), .A (n_12_56), .B (n_18_53), .C1 (n_22_51), .C2 (n_25_51) );
AOI211_X1 g_7_60 (.ZN (n_7_60), .A (n_10_57), .B (n_16_54), .C1 (n_20_52), .C2 (n_23_52) );
AOI211_X1 g_9_59 (.ZN (n_9_59), .A (n_8_58), .B (n_14_55), .C1 (n_18_53), .C2 (n_21_53) );
AOI211_X1 g_11_58 (.ZN (n_11_58), .A (n_7_60), .B (n_12_56), .C1 (n_16_54), .C2 (n_22_51) );
AOI211_X1 g_13_57 (.ZN (n_13_57), .A (n_9_59), .B (n_10_57), .C1 (n_14_55), .C2 (n_20_52) );
AOI211_X1 g_15_56 (.ZN (n_15_56), .A (n_11_58), .B (n_8_58), .C1 (n_12_56), .C2 (n_18_53) );
AOI211_X1 g_17_55 (.ZN (n_17_55), .A (n_13_57), .B (n_7_60), .C1 (n_10_57), .C2 (n_16_54) );
AOI211_X1 g_19_54 (.ZN (n_19_54), .A (n_15_56), .B (n_9_59), .C1 (n_8_58), .C2 (n_14_55) );
AOI211_X1 g_18_56 (.ZN (n_18_56), .A (n_17_55), .B (n_11_58), .C1 (n_7_60), .C2 (n_12_56) );
AOI211_X1 g_20_55 (.ZN (n_20_55), .A (n_19_54), .B (n_13_57), .C1 (n_9_59), .C2 (n_10_57) );
AOI211_X1 g_22_54 (.ZN (n_22_54), .A (n_18_56), .B (n_15_56), .C1 (n_11_58), .C2 (n_8_58) );
AOI211_X1 g_24_53 (.ZN (n_24_53), .A (n_20_55), .B (n_17_55), .C1 (n_13_57), .C2 (n_7_60) );
AOI211_X1 g_26_52 (.ZN (n_26_52), .A (n_22_54), .B (n_19_54), .C1 (n_15_56), .C2 (n_9_59) );
AOI211_X1 g_24_51 (.ZN (n_24_51), .A (n_24_53), .B (n_18_56), .C1 (n_17_55), .C2 (n_11_58) );
AOI211_X1 g_26_50 (.ZN (n_26_50), .A (n_26_52), .B (n_20_55), .C1 (n_19_54), .C2 (n_13_57) );
AOI211_X1 g_28_49 (.ZN (n_28_49), .A (n_24_51), .B (n_22_54), .C1 (n_18_56), .C2 (n_15_56) );
AOI211_X1 g_30_48 (.ZN (n_30_48), .A (n_26_50), .B (n_24_53), .C1 (n_20_55), .C2 (n_17_55) );
AOI211_X1 g_32_47 (.ZN (n_32_47), .A (n_28_49), .B (n_26_52), .C1 (n_22_54), .C2 (n_19_54) );
AOI211_X1 g_34_46 (.ZN (n_34_46), .A (n_30_48), .B (n_24_51), .C1 (n_24_53), .C2 (n_18_56) );
AOI211_X1 g_36_45 (.ZN (n_36_45), .A (n_32_47), .B (n_26_50), .C1 (n_26_52), .C2 (n_20_55) );
AOI211_X1 g_38_44 (.ZN (n_38_44), .A (n_34_46), .B (n_28_49), .C1 (n_24_51), .C2 (n_22_54) );
AOI211_X1 g_40_43 (.ZN (n_40_43), .A (n_36_45), .B (n_30_48), .C1 (n_26_50), .C2 (n_24_53) );
AOI211_X1 g_42_42 (.ZN (n_42_42), .A (n_38_44), .B (n_32_47), .C1 (n_28_49), .C2 (n_26_52) );
AOI211_X1 g_44_41 (.ZN (n_44_41), .A (n_40_43), .B (n_34_46), .C1 (n_30_48), .C2 (n_24_51) );
AOI211_X1 g_46_40 (.ZN (n_46_40), .A (n_42_42), .B (n_36_45), .C1 (n_32_47), .C2 (n_26_50) );
AOI211_X1 g_48_39 (.ZN (n_48_39), .A (n_44_41), .B (n_38_44), .C1 (n_34_46), .C2 (n_28_49) );
AOI211_X1 g_50_38 (.ZN (n_50_38), .A (n_46_40), .B (n_40_43), .C1 (n_36_45), .C2 (n_30_48) );
AOI211_X1 g_52_37 (.ZN (n_52_37), .A (n_48_39), .B (n_42_42), .C1 (n_38_44), .C2 (n_32_47) );
AOI211_X1 g_54_36 (.ZN (n_54_36), .A (n_50_38), .B (n_44_41), .C1 (n_40_43), .C2 (n_34_46) );
AOI211_X1 g_56_35 (.ZN (n_56_35), .A (n_52_37), .B (n_46_40), .C1 (n_42_42), .C2 (n_36_45) );
AOI211_X1 g_58_34 (.ZN (n_58_34), .A (n_54_36), .B (n_48_39), .C1 (n_44_41), .C2 (n_38_44) );
AOI211_X1 g_60_33 (.ZN (n_60_33), .A (n_56_35), .B (n_50_38), .C1 (n_46_40), .C2 (n_40_43) );
AOI211_X1 g_59_35 (.ZN (n_59_35), .A (n_58_34), .B (n_52_37), .C1 (n_48_39), .C2 (n_42_42) );
AOI211_X1 g_57_36 (.ZN (n_57_36), .A (n_60_33), .B (n_54_36), .C1 (n_50_38), .C2 (n_44_41) );
AOI211_X1 g_55_37 (.ZN (n_55_37), .A (n_59_35), .B (n_56_35), .C1 (n_52_37), .C2 (n_46_40) );
AOI211_X1 g_53_38 (.ZN (n_53_38), .A (n_57_36), .B (n_58_34), .C1 (n_54_36), .C2 (n_48_39) );
AOI211_X1 g_51_39 (.ZN (n_51_39), .A (n_55_37), .B (n_60_33), .C1 (n_56_35), .C2 (n_50_38) );
AOI211_X1 g_49_40 (.ZN (n_49_40), .A (n_53_38), .B (n_59_35), .C1 (n_58_34), .C2 (n_52_37) );
AOI211_X1 g_47_41 (.ZN (n_47_41), .A (n_51_39), .B (n_57_36), .C1 (n_60_33), .C2 (n_54_36) );
AOI211_X1 g_45_40 (.ZN (n_45_40), .A (n_49_40), .B (n_55_37), .C1 (n_59_35), .C2 (n_56_35) );
AOI211_X1 g_43_41 (.ZN (n_43_41), .A (n_47_41), .B (n_53_38), .C1 (n_57_36), .C2 (n_58_34) );
AOI211_X1 g_41_42 (.ZN (n_41_42), .A (n_45_40), .B (n_51_39), .C1 (n_55_37), .C2 (n_60_33) );
AOI211_X1 g_40_44 (.ZN (n_40_44), .A (n_43_41), .B (n_49_40), .C1 (n_53_38), .C2 (n_59_35) );
AOI211_X1 g_42_43 (.ZN (n_42_43), .A (n_41_42), .B (n_47_41), .C1 (n_51_39), .C2 (n_57_36) );
AOI211_X1 g_44_42 (.ZN (n_44_42), .A (n_40_44), .B (n_45_40), .C1 (n_49_40), .C2 (n_55_37) );
AOI211_X1 g_46_41 (.ZN (n_46_41), .A (n_42_43), .B (n_43_41), .C1 (n_47_41), .C2 (n_53_38) );
AOI211_X1 g_48_40 (.ZN (n_48_40), .A (n_44_42), .B (n_41_42), .C1 (n_45_40), .C2 (n_51_39) );
AOI211_X1 g_50_39 (.ZN (n_50_39), .A (n_46_41), .B (n_40_44), .C1 (n_43_41), .C2 (n_49_40) );
AOI211_X1 g_52_38 (.ZN (n_52_38), .A (n_48_40), .B (n_42_43), .C1 (n_41_42), .C2 (n_47_41) );
AOI211_X1 g_54_37 (.ZN (n_54_37), .A (n_50_39), .B (n_44_42), .C1 (n_40_44), .C2 (n_45_40) );
AOI211_X1 g_56_36 (.ZN (n_56_36), .A (n_52_38), .B (n_46_41), .C1 (n_42_43), .C2 (n_43_41) );
AOI211_X1 g_58_35 (.ZN (n_58_35), .A (n_54_37), .B (n_48_40), .C1 (n_44_42), .C2 (n_41_42) );
AOI211_X1 g_60_34 (.ZN (n_60_34), .A (n_56_36), .B (n_50_39), .C1 (n_46_41), .C2 (n_40_44) );
AOI211_X1 g_62_35 (.ZN (n_62_35), .A (n_58_35), .B (n_52_38), .C1 (n_48_40), .C2 (n_42_43) );
AOI211_X1 g_60_36 (.ZN (n_60_36), .A (n_60_34), .B (n_54_37), .C1 (n_50_39), .C2 (n_44_42) );
AOI211_X1 g_58_37 (.ZN (n_58_37), .A (n_62_35), .B (n_56_36), .C1 (n_52_38), .C2 (n_46_41) );
AOI211_X1 g_56_38 (.ZN (n_56_38), .A (n_60_36), .B (n_58_35), .C1 (n_54_37), .C2 (n_48_40) );
AOI211_X1 g_54_39 (.ZN (n_54_39), .A (n_58_37), .B (n_60_34), .C1 (n_56_36), .C2 (n_50_39) );
AOI211_X1 g_52_40 (.ZN (n_52_40), .A (n_56_38), .B (n_62_35), .C1 (n_58_35), .C2 (n_52_38) );
AOI211_X1 g_50_41 (.ZN (n_50_41), .A (n_54_39), .B (n_60_36), .C1 (n_60_34), .C2 (n_54_37) );
AOI211_X1 g_48_42 (.ZN (n_48_42), .A (n_52_40), .B (n_58_37), .C1 (n_62_35), .C2 (n_56_36) );
AOI211_X1 g_46_43 (.ZN (n_46_43), .A (n_50_41), .B (n_56_38), .C1 (n_60_36), .C2 (n_58_35) );
AOI211_X1 g_44_44 (.ZN (n_44_44), .A (n_48_42), .B (n_54_39), .C1 (n_58_37), .C2 (n_60_34) );
AOI211_X1 g_45_42 (.ZN (n_45_42), .A (n_46_43), .B (n_52_40), .C1 (n_56_38), .C2 (n_62_35) );
AOI211_X1 g_43_43 (.ZN (n_43_43), .A (n_44_44), .B (n_50_41), .C1 (n_54_39), .C2 (n_60_36) );
AOI211_X1 g_41_44 (.ZN (n_41_44), .A (n_45_42), .B (n_48_42), .C1 (n_52_40), .C2 (n_58_37) );
AOI211_X1 g_39_45 (.ZN (n_39_45), .A (n_43_43), .B (n_46_43), .C1 (n_50_41), .C2 (n_56_38) );
AOI211_X1 g_37_46 (.ZN (n_37_46), .A (n_41_44), .B (n_44_44), .C1 (n_48_42), .C2 (n_54_39) );
AOI211_X1 g_35_47 (.ZN (n_35_47), .A (n_39_45), .B (n_45_42), .C1 (n_46_43), .C2 (n_52_40) );
AOI211_X1 g_33_48 (.ZN (n_33_48), .A (n_37_46), .B (n_43_43), .C1 (n_44_44), .C2 (n_50_41) );
AOI211_X1 g_31_49 (.ZN (n_31_49), .A (n_35_47), .B (n_41_44), .C1 (n_45_42), .C2 (n_48_42) );
AOI211_X1 g_29_50 (.ZN (n_29_50), .A (n_33_48), .B (n_39_45), .C1 (n_43_43), .C2 (n_46_43) );
AOI211_X1 g_27_51 (.ZN (n_27_51), .A (n_31_49), .B (n_37_46), .C1 (n_41_44), .C2 (n_44_44) );
AOI211_X1 g_25_52 (.ZN (n_25_52), .A (n_29_50), .B (n_35_47), .C1 (n_39_45), .C2 (n_45_42) );
AOI211_X1 g_23_53 (.ZN (n_23_53), .A (n_27_51), .B (n_33_48), .C1 (n_37_46), .C2 (n_43_43) );
AOI211_X1 g_21_54 (.ZN (n_21_54), .A (n_25_52), .B (n_31_49), .C1 (n_35_47), .C2 (n_41_44) );
AOI211_X1 g_19_55 (.ZN (n_19_55), .A (n_23_53), .B (n_29_50), .C1 (n_33_48), .C2 (n_39_45) );
AOI211_X1 g_17_56 (.ZN (n_17_56), .A (n_21_54), .B (n_27_51), .C1 (n_31_49), .C2 (n_37_46) );
AOI211_X1 g_15_57 (.ZN (n_15_57), .A (n_19_55), .B (n_25_52), .C1 (n_29_50), .C2 (n_35_47) );
AOI211_X1 g_13_58 (.ZN (n_13_58), .A (n_17_56), .B (n_23_53), .C1 (n_27_51), .C2 (n_33_48) );
AOI211_X1 g_11_59 (.ZN (n_11_59), .A (n_15_57), .B (n_21_54), .C1 (n_25_52), .C2 (n_31_49) );
AOI211_X1 g_9_60 (.ZN (n_9_60), .A (n_13_58), .B (n_19_55), .C1 (n_23_53), .C2 (n_29_50) );
AOI211_X1 g_10_58 (.ZN (n_10_58), .A (n_11_59), .B (n_17_56), .C1 (n_21_54), .C2 (n_27_51) );
AOI211_X1 g_12_59 (.ZN (n_12_59), .A (n_9_60), .B (n_15_57), .C1 (n_19_55), .C2 (n_25_52) );
AOI211_X1 g_14_58 (.ZN (n_14_58), .A (n_10_58), .B (n_13_58), .C1 (n_17_56), .C2 (n_23_53) );
AOI211_X1 g_16_57 (.ZN (n_16_57), .A (n_12_59), .B (n_11_59), .C1 (n_15_57), .C2 (n_21_54) );
AOI211_X1 g_15_59 (.ZN (n_15_59), .A (n_14_58), .B (n_9_60), .C1 (n_13_58), .C2 (n_19_55) );
AOI211_X1 g_14_57 (.ZN (n_14_57), .A (n_16_57), .B (n_10_58), .C1 (n_11_59), .C2 (n_17_56) );
AOI211_X1 g_16_56 (.ZN (n_16_56), .A (n_15_59), .B (n_12_59), .C1 (n_9_60), .C2 (n_15_57) );
AOI211_X1 g_18_55 (.ZN (n_18_55), .A (n_14_57), .B (n_14_58), .C1 (n_10_58), .C2 (n_13_58) );
AOI211_X1 g_20_54 (.ZN (n_20_54), .A (n_16_56), .B (n_16_57), .C1 (n_12_59), .C2 (n_11_59) );
AOI211_X1 g_22_53 (.ZN (n_22_53), .A (n_18_55), .B (n_15_59), .C1 (n_14_58), .C2 (n_9_60) );
AOI211_X1 g_24_52 (.ZN (n_24_52), .A (n_20_54), .B (n_14_57), .C1 (n_16_57), .C2 (n_10_58) );
AOI211_X1 g_23_54 (.ZN (n_23_54), .A (n_22_53), .B (n_16_56), .C1 (n_15_59), .C2 (n_12_59) );
AOI211_X1 g_25_53 (.ZN (n_25_53), .A (n_24_52), .B (n_18_55), .C1 (n_14_57), .C2 (n_14_58) );
AOI211_X1 g_27_52 (.ZN (n_27_52), .A (n_23_54), .B (n_20_54), .C1 (n_16_56), .C2 (n_16_57) );
AOI211_X1 g_28_50 (.ZN (n_28_50), .A (n_25_53), .B (n_22_53), .C1 (n_18_55), .C2 (n_15_59) );
AOI211_X1 g_30_49 (.ZN (n_30_49), .A (n_27_52), .B (n_24_52), .C1 (n_20_54), .C2 (n_14_57) );
AOI211_X1 g_32_48 (.ZN (n_32_48), .A (n_28_50), .B (n_23_54), .C1 (n_22_53), .C2 (n_16_56) );
AOI211_X1 g_34_47 (.ZN (n_34_47), .A (n_30_49), .B (n_25_53), .C1 (n_24_52), .C2 (n_18_55) );
AOI211_X1 g_36_46 (.ZN (n_36_46), .A (n_32_48), .B (n_27_52), .C1 (n_23_54), .C2 (n_20_54) );
AOI211_X1 g_38_45 (.ZN (n_38_45), .A (n_34_47), .B (n_28_50), .C1 (n_25_53), .C2 (n_22_53) );
AOI211_X1 g_37_47 (.ZN (n_37_47), .A (n_36_46), .B (n_30_49), .C1 (n_27_52), .C2 (n_24_52) );
AOI211_X1 g_39_46 (.ZN (n_39_46), .A (n_38_45), .B (n_32_48), .C1 (n_28_50), .C2 (n_23_54) );
AOI211_X1 g_41_45 (.ZN (n_41_45), .A (n_37_47), .B (n_34_47), .C1 (n_30_49), .C2 (n_25_53) );
AOI211_X1 g_43_44 (.ZN (n_43_44), .A (n_39_46), .B (n_36_46), .C1 (n_32_48), .C2 (n_27_52) );
AOI211_X1 g_45_43 (.ZN (n_45_43), .A (n_41_45), .B (n_38_45), .C1 (n_34_47), .C2 (n_28_50) );
AOI211_X1 g_47_42 (.ZN (n_47_42), .A (n_43_44), .B (n_37_47), .C1 (n_36_46), .C2 (n_30_49) );
AOI211_X1 g_49_41 (.ZN (n_49_41), .A (n_45_43), .B (n_39_46), .C1 (n_38_45), .C2 (n_32_48) );
AOI211_X1 g_51_40 (.ZN (n_51_40), .A (n_47_42), .B (n_41_45), .C1 (n_37_47), .C2 (n_34_47) );
AOI211_X1 g_53_39 (.ZN (n_53_39), .A (n_49_41), .B (n_43_44), .C1 (n_39_46), .C2 (n_36_46) );
AOI211_X1 g_55_38 (.ZN (n_55_38), .A (n_51_40), .B (n_45_43), .C1 (n_41_45), .C2 (n_38_45) );
AOI211_X1 g_57_37 (.ZN (n_57_37), .A (n_53_39), .B (n_47_42), .C1 (n_43_44), .C2 (n_37_47) );
AOI211_X1 g_59_36 (.ZN (n_59_36), .A (n_55_38), .B (n_49_41), .C1 (n_45_43), .C2 (n_39_46) );
AOI211_X1 g_61_35 (.ZN (n_61_35), .A (n_57_37), .B (n_51_40), .C1 (n_47_42), .C2 (n_41_45) );
AOI211_X1 g_62_37 (.ZN (n_62_37), .A (n_59_36), .B (n_53_39), .C1 (n_49_41), .C2 (n_43_44) );
AOI211_X1 g_64_36 (.ZN (n_64_36), .A (n_61_35), .B (n_55_38), .C1 (n_51_40), .C2 (n_45_43) );
AOI211_X1 g_66_35 (.ZN (n_66_35), .A (n_62_37), .B (n_57_37), .C1 (n_53_39), .C2 (n_47_42) );
AOI211_X1 g_68_34 (.ZN (n_68_34), .A (n_64_36), .B (n_59_36), .C1 (n_55_38), .C2 (n_49_41) );
AOI211_X1 g_70_33 (.ZN (n_70_33), .A (n_66_35), .B (n_61_35), .C1 (n_57_37), .C2 (n_51_40) );
AOI211_X1 g_72_32 (.ZN (n_72_32), .A (n_68_34), .B (n_62_37), .C1 (n_59_36), .C2 (n_53_39) );
AOI211_X1 g_73_30 (.ZN (n_73_30), .A (n_70_33), .B (n_64_36), .C1 (n_61_35), .C2 (n_55_38) );
AOI211_X1 g_75_29 (.ZN (n_75_29), .A (n_72_32), .B (n_66_35), .C1 (n_62_37), .C2 (n_57_37) );
AOI211_X1 g_77_28 (.ZN (n_77_28), .A (n_73_30), .B (n_68_34), .C1 (n_64_36), .C2 (n_59_36) );
AOI211_X1 g_79_27 (.ZN (n_79_27), .A (n_75_29), .B (n_70_33), .C1 (n_66_35), .C2 (n_61_35) );
AOI211_X1 g_81_26 (.ZN (n_81_26), .A (n_77_28), .B (n_72_32), .C1 (n_68_34), .C2 (n_62_37) );
AOI211_X1 g_83_25 (.ZN (n_83_25), .A (n_79_27), .B (n_73_30), .C1 (n_70_33), .C2 (n_64_36) );
AOI211_X1 g_85_24 (.ZN (n_85_24), .A (n_81_26), .B (n_75_29), .C1 (n_72_32), .C2 (n_66_35) );
AOI211_X1 g_87_23 (.ZN (n_87_23), .A (n_83_25), .B (n_77_28), .C1 (n_73_30), .C2 (n_68_34) );
AOI211_X1 g_89_22 (.ZN (n_89_22), .A (n_85_24), .B (n_79_27), .C1 (n_75_29), .C2 (n_70_33) );
AOI211_X1 g_91_21 (.ZN (n_91_21), .A (n_87_23), .B (n_81_26), .C1 (n_77_28), .C2 (n_72_32) );
AOI211_X1 g_93_20 (.ZN (n_93_20), .A (n_89_22), .B (n_83_25), .C1 (n_79_27), .C2 (n_73_30) );
AOI211_X1 g_95_21 (.ZN (n_95_21), .A (n_91_21), .B (n_85_24), .C1 (n_81_26), .C2 (n_75_29) );
AOI211_X1 g_93_22 (.ZN (n_93_22), .A (n_93_20), .B (n_87_23), .C1 (n_83_25), .C2 (n_77_28) );
AOI211_X1 g_91_23 (.ZN (n_91_23), .A (n_95_21), .B (n_89_22), .C1 (n_85_24), .C2 (n_79_27) );
AOI211_X1 g_89_24 (.ZN (n_89_24), .A (n_93_22), .B (n_91_21), .C1 (n_87_23), .C2 (n_81_26) );
AOI211_X1 g_87_25 (.ZN (n_87_25), .A (n_91_23), .B (n_93_20), .C1 (n_89_22), .C2 (n_83_25) );
AOI211_X1 g_85_26 (.ZN (n_85_26), .A (n_89_24), .B (n_95_21), .C1 (n_91_21), .C2 (n_85_24) );
AOI211_X1 g_83_27 (.ZN (n_83_27), .A (n_87_25), .B (n_93_22), .C1 (n_93_20), .C2 (n_87_23) );
AOI211_X1 g_81_28 (.ZN (n_81_28), .A (n_85_26), .B (n_91_23), .C1 (n_95_21), .C2 (n_89_22) );
AOI211_X1 g_79_29 (.ZN (n_79_29), .A (n_83_27), .B (n_89_24), .C1 (n_93_22), .C2 (n_91_21) );
AOI211_X1 g_80_27 (.ZN (n_80_27), .A (n_81_28), .B (n_87_25), .C1 (n_91_23), .C2 (n_93_20) );
AOI211_X1 g_78_28 (.ZN (n_78_28), .A (n_79_29), .B (n_85_26), .C1 (n_89_24), .C2 (n_95_21) );
AOI211_X1 g_76_29 (.ZN (n_76_29), .A (n_80_27), .B (n_83_27), .C1 (n_87_25), .C2 (n_93_22) );
AOI211_X1 g_75_31 (.ZN (n_75_31), .A (n_78_28), .B (n_81_28), .C1 (n_85_26), .C2 (n_91_23) );
AOI211_X1 g_77_30 (.ZN (n_77_30), .A (n_76_29), .B (n_79_29), .C1 (n_83_27), .C2 (n_89_24) );
AOI211_X1 g_76_32 (.ZN (n_76_32), .A (n_75_31), .B (n_80_27), .C1 (n_81_28), .C2 (n_87_25) );
AOI211_X1 g_74_31 (.ZN (n_74_31), .A (n_77_30), .B (n_78_28), .C1 (n_79_29), .C2 (n_85_26) );
AOI211_X1 g_76_30 (.ZN (n_76_30), .A (n_76_32), .B (n_76_29), .C1 (n_80_27), .C2 (n_83_27) );
AOI211_X1 g_78_29 (.ZN (n_78_29), .A (n_74_31), .B (n_75_31), .C1 (n_78_28), .C2 (n_81_28) );
AOI211_X1 g_80_28 (.ZN (n_80_28), .A (n_76_30), .B (n_77_30), .C1 (n_76_29), .C2 (n_79_29) );
AOI211_X1 g_82_27 (.ZN (n_82_27), .A (n_78_29), .B (n_76_32), .C1 (n_75_31), .C2 (n_80_27) );
AOI211_X1 g_84_26 (.ZN (n_84_26), .A (n_80_28), .B (n_74_31), .C1 (n_77_30), .C2 (n_78_28) );
AOI211_X1 g_86_25 (.ZN (n_86_25), .A (n_82_27), .B (n_76_30), .C1 (n_76_32), .C2 (n_76_29) );
AOI211_X1 g_88_24 (.ZN (n_88_24), .A (n_84_26), .B (n_78_29), .C1 (n_74_31), .C2 (n_75_31) );
AOI211_X1 g_90_23 (.ZN (n_90_23), .A (n_86_25), .B (n_80_28), .C1 (n_76_30), .C2 (n_77_30) );
AOI211_X1 g_92_22 (.ZN (n_92_22), .A (n_88_24), .B (n_82_27), .C1 (n_78_29), .C2 (n_76_32) );
AOI211_X1 g_94_21 (.ZN (n_94_21), .A (n_90_23), .B (n_84_26), .C1 (n_80_28), .C2 (n_74_31) );
AOI211_X1 g_96_20 (.ZN (n_96_20), .A (n_92_22), .B (n_86_25), .C1 (n_82_27), .C2 (n_76_30) );
AOI211_X1 g_98_19 (.ZN (n_98_19), .A (n_94_21), .B (n_88_24), .C1 (n_84_26), .C2 (n_78_29) );
AOI211_X1 g_100_20 (.ZN (n_100_20), .A (n_96_20), .B (n_90_23), .C1 (n_86_25), .C2 (n_80_28) );
AOI211_X1 g_98_21 (.ZN (n_98_21), .A (n_98_19), .B (n_92_22), .C1 (n_88_24), .C2 (n_82_27) );
AOI211_X1 g_96_22 (.ZN (n_96_22), .A (n_100_20), .B (n_94_21), .C1 (n_90_23), .C2 (n_84_26) );
AOI211_X1 g_94_23 (.ZN (n_94_23), .A (n_98_21), .B (n_96_20), .C1 (n_92_22), .C2 (n_86_25) );
AOI211_X1 g_92_24 (.ZN (n_92_24), .A (n_96_22), .B (n_98_19), .C1 (n_94_21), .C2 (n_88_24) );
AOI211_X1 g_90_25 (.ZN (n_90_25), .A (n_94_23), .B (n_100_20), .C1 (n_96_20), .C2 (n_90_23) );
AOI211_X1 g_88_26 (.ZN (n_88_26), .A (n_92_24), .B (n_98_21), .C1 (n_98_19), .C2 (n_92_22) );
AOI211_X1 g_86_27 (.ZN (n_86_27), .A (n_90_25), .B (n_96_22), .C1 (n_100_20), .C2 (n_94_21) );
AOI211_X1 g_84_28 (.ZN (n_84_28), .A (n_88_26), .B (n_94_23), .C1 (n_98_21), .C2 (n_96_20) );
AOI211_X1 g_82_29 (.ZN (n_82_29), .A (n_86_27), .B (n_92_24), .C1 (n_96_22), .C2 (n_98_19) );
AOI211_X1 g_80_30 (.ZN (n_80_30), .A (n_84_28), .B (n_90_25), .C1 (n_94_23), .C2 (n_100_20) );
AOI211_X1 g_78_31 (.ZN (n_78_31), .A (n_82_29), .B (n_88_26), .C1 (n_92_24), .C2 (n_98_21) );
AOI211_X1 g_77_33 (.ZN (n_77_33), .A (n_80_30), .B (n_86_27), .C1 (n_90_25), .C2 (n_96_22) );
AOI211_X1 g_76_31 (.ZN (n_76_31), .A (n_78_31), .B (n_84_28), .C1 (n_88_26), .C2 (n_94_23) );
AOI211_X1 g_78_30 (.ZN (n_78_30), .A (n_77_33), .B (n_82_29), .C1 (n_86_27), .C2 (n_92_24) );
AOI211_X1 g_80_29 (.ZN (n_80_29), .A (n_76_31), .B (n_80_30), .C1 (n_84_28), .C2 (n_90_25) );
AOI211_X1 g_82_28 (.ZN (n_82_28), .A (n_78_30), .B (n_78_31), .C1 (n_82_29), .C2 (n_88_26) );
AOI211_X1 g_84_27 (.ZN (n_84_27), .A (n_80_29), .B (n_77_33), .C1 (n_80_30), .C2 (n_86_27) );
AOI211_X1 g_86_26 (.ZN (n_86_26), .A (n_82_28), .B (n_76_31), .C1 (n_78_31), .C2 (n_84_28) );
AOI211_X1 g_88_25 (.ZN (n_88_25), .A (n_84_27), .B (n_78_30), .C1 (n_77_33), .C2 (n_82_29) );
AOI211_X1 g_90_24 (.ZN (n_90_24), .A (n_86_26), .B (n_80_29), .C1 (n_76_31), .C2 (n_80_30) );
AOI211_X1 g_92_23 (.ZN (n_92_23), .A (n_88_25), .B (n_82_28), .C1 (n_78_30), .C2 (n_78_31) );
AOI211_X1 g_91_25 (.ZN (n_91_25), .A (n_90_24), .B (n_84_27), .C1 (n_80_29), .C2 (n_77_33) );
AOI211_X1 g_93_24 (.ZN (n_93_24), .A (n_92_23), .B (n_86_26), .C1 (n_82_28), .C2 (n_76_31) );
AOI211_X1 g_95_23 (.ZN (n_95_23), .A (n_91_25), .B (n_88_25), .C1 (n_84_27), .C2 (n_78_30) );
AOI211_X1 g_97_22 (.ZN (n_97_22), .A (n_93_24), .B (n_90_24), .C1 (n_86_26), .C2 (n_80_29) );
AOI211_X1 g_99_23 (.ZN (n_99_23), .A (n_95_23), .B (n_92_23), .C1 (n_88_25), .C2 (n_82_28) );
AOI211_X1 g_100_25 (.ZN (n_100_25), .A (n_97_22), .B (n_91_25), .C1 (n_90_24), .C2 (n_84_27) );
AOI211_X1 g_98_24 (.ZN (n_98_24), .A (n_99_23), .B (n_93_24), .C1 (n_92_23), .C2 (n_86_26) );
AOI211_X1 g_99_22 (.ZN (n_99_22), .A (n_100_25), .B (n_95_23), .C1 (n_91_25), .C2 (n_88_25) );
AOI211_X1 g_97_21 (.ZN (n_97_21), .A (n_98_24), .B (n_97_22), .C1 (n_93_24), .C2 (n_90_24) );
AOI211_X1 g_96_23 (.ZN (n_96_23), .A (n_99_22), .B (n_99_23), .C1 (n_95_23), .C2 (n_92_23) );
AOI211_X1 g_94_24 (.ZN (n_94_24), .A (n_97_21), .B (n_100_25), .C1 (n_97_22), .C2 (n_91_25) );
AOI211_X1 g_95_22 (.ZN (n_95_22), .A (n_96_23), .B (n_98_24), .C1 (n_99_23), .C2 (n_93_24) );
AOI211_X1 g_97_23 (.ZN (n_97_23), .A (n_94_24), .B (n_99_22), .C1 (n_100_25), .C2 (n_95_23) );
AOI211_X1 g_96_25 (.ZN (n_96_25), .A (n_95_22), .B (n_97_21), .C1 (n_98_24), .C2 (n_97_22) );
AOI211_X1 g_98_26 (.ZN (n_98_26), .A (n_97_23), .B (n_96_23), .C1 (n_99_22), .C2 (n_99_23) );
AOI211_X1 g_97_24 (.ZN (n_97_24), .A (n_96_25), .B (n_94_24), .C1 (n_97_21), .C2 (n_100_25) );
AOI211_X1 g_95_25 (.ZN (n_95_25), .A (n_98_26), .B (n_95_22), .C1 (n_96_23), .C2 (n_98_24) );
AOI211_X1 g_93_26 (.ZN (n_93_26), .A (n_97_24), .B (n_97_23), .C1 (n_94_24), .C2 (n_99_22) );
AOI211_X1 g_91_27 (.ZN (n_91_27), .A (n_95_25), .B (n_96_25), .C1 (n_95_22), .C2 (n_97_21) );
AOI211_X1 g_89_26 (.ZN (n_89_26), .A (n_93_26), .B (n_98_26), .C1 (n_97_23), .C2 (n_96_23) );
AOI211_X1 g_87_27 (.ZN (n_87_27), .A (n_91_27), .B (n_97_24), .C1 (n_96_25), .C2 (n_94_24) );
AOI211_X1 g_85_28 (.ZN (n_85_28), .A (n_89_26), .B (n_95_25), .C1 (n_98_26), .C2 (n_95_22) );
AOI211_X1 g_83_29 (.ZN (n_83_29), .A (n_87_27), .B (n_93_26), .C1 (n_97_24), .C2 (n_97_23) );
AOI211_X1 g_81_30 (.ZN (n_81_30), .A (n_85_28), .B (n_91_27), .C1 (n_95_25), .C2 (n_96_25) );
AOI211_X1 g_79_31 (.ZN (n_79_31), .A (n_83_29), .B (n_89_26), .C1 (n_93_26), .C2 (n_98_26) );
AOI211_X1 g_77_32 (.ZN (n_77_32), .A (n_81_30), .B (n_87_27), .C1 (n_91_27), .C2 (n_97_24) );
AOI211_X1 g_75_33 (.ZN (n_75_33), .A (n_79_31), .B (n_85_28), .C1 (n_89_26), .C2 (n_95_25) );
AOI211_X1 g_73_34 (.ZN (n_73_34), .A (n_77_32), .B (n_83_29), .C1 (n_87_27), .C2 (n_93_26) );
AOI211_X1 g_74_32 (.ZN (n_74_32), .A (n_75_33), .B (n_81_30), .C1 (n_85_28), .C2 (n_91_27) );
AOI211_X1 g_72_33 (.ZN (n_72_33), .A (n_73_34), .B (n_79_31), .C1 (n_83_29), .C2 (n_89_26) );
AOI211_X1 g_73_31 (.ZN (n_73_31), .A (n_74_32), .B (n_77_32), .C1 (n_81_30), .C2 (n_87_27) );
AOI211_X1 g_71_32 (.ZN (n_71_32), .A (n_72_33), .B (n_75_33), .C1 (n_79_31), .C2 (n_85_28) );
AOI211_X1 g_69_33 (.ZN (n_69_33), .A (n_73_31), .B (n_73_34), .C1 (n_77_32), .C2 (n_83_29) );
AOI211_X1 g_67_34 (.ZN (n_67_34), .A (n_71_32), .B (n_74_32), .C1 (n_75_33), .C2 (n_81_30) );
AOI211_X1 g_65_35 (.ZN (n_65_35), .A (n_69_33), .B (n_72_33), .C1 (n_73_34), .C2 (n_79_31) );
AOI211_X1 g_63_36 (.ZN (n_63_36), .A (n_67_34), .B (n_73_31), .C1 (n_74_32), .C2 (n_77_32) );
AOI211_X1 g_62_34 (.ZN (n_62_34), .A (n_65_35), .B (n_71_32), .C1 (n_72_33), .C2 (n_75_33) );
AOI211_X1 g_60_35 (.ZN (n_60_35), .A (n_63_36), .B (n_69_33), .C1 (n_73_31), .C2 (n_73_34) );
AOI211_X1 g_58_36 (.ZN (n_58_36), .A (n_62_34), .B (n_67_34), .C1 (n_71_32), .C2 (n_74_32) );
AOI211_X1 g_56_37 (.ZN (n_56_37), .A (n_60_35), .B (n_65_35), .C1 (n_69_33), .C2 (n_72_33) );
AOI211_X1 g_54_38 (.ZN (n_54_38), .A (n_58_36), .B (n_63_36), .C1 (n_67_34), .C2 (n_73_31) );
AOI211_X1 g_52_39 (.ZN (n_52_39), .A (n_56_37), .B (n_62_34), .C1 (n_65_35), .C2 (n_71_32) );
AOI211_X1 g_50_40 (.ZN (n_50_40), .A (n_54_38), .B (n_60_35), .C1 (n_63_36), .C2 (n_69_33) );
AOI211_X1 g_48_41 (.ZN (n_48_41), .A (n_52_39), .B (n_58_36), .C1 (n_62_34), .C2 (n_67_34) );
AOI211_X1 g_46_42 (.ZN (n_46_42), .A (n_50_40), .B (n_56_37), .C1 (n_60_35), .C2 (n_65_35) );
AOI211_X1 g_44_43 (.ZN (n_44_43), .A (n_48_41), .B (n_54_38), .C1 (n_58_36), .C2 (n_63_36) );
AOI211_X1 g_42_44 (.ZN (n_42_44), .A (n_46_42), .B (n_52_39), .C1 (n_56_37), .C2 (n_62_34) );
AOI211_X1 g_40_45 (.ZN (n_40_45), .A (n_44_43), .B (n_50_40), .C1 (n_54_38), .C2 (n_60_35) );
AOI211_X1 g_38_46 (.ZN (n_38_46), .A (n_42_44), .B (n_48_41), .C1 (n_52_39), .C2 (n_58_36) );
AOI211_X1 g_36_47 (.ZN (n_36_47), .A (n_40_45), .B (n_46_42), .C1 (n_50_40), .C2 (n_56_37) );
AOI211_X1 g_34_48 (.ZN (n_34_48), .A (n_38_46), .B (n_44_43), .C1 (n_48_41), .C2 (n_54_38) );
AOI211_X1 g_32_49 (.ZN (n_32_49), .A (n_36_47), .B (n_42_44), .C1 (n_46_42), .C2 (n_52_39) );
AOI211_X1 g_30_50 (.ZN (n_30_50), .A (n_34_48), .B (n_40_45), .C1 (n_44_43), .C2 (n_50_40) );
AOI211_X1 g_28_51 (.ZN (n_28_51), .A (n_32_49), .B (n_38_46), .C1 (n_42_44), .C2 (n_48_41) );
AOI211_X1 g_27_53 (.ZN (n_27_53), .A (n_30_50), .B (n_36_47), .C1 (n_40_45), .C2 (n_46_42) );
AOI211_X1 g_29_52 (.ZN (n_29_52), .A (n_28_51), .B (n_34_48), .C1 (n_38_46), .C2 (n_44_43) );
AOI211_X1 g_31_51 (.ZN (n_31_51), .A (n_27_53), .B (n_32_49), .C1 (n_36_47), .C2 (n_42_44) );
AOI211_X1 g_33_50 (.ZN (n_33_50), .A (n_29_52), .B (n_30_50), .C1 (n_34_48), .C2 (n_40_45) );
AOI211_X1 g_35_49 (.ZN (n_35_49), .A (n_31_51), .B (n_28_51), .C1 (n_32_49), .C2 (n_38_46) );
AOI211_X1 g_37_48 (.ZN (n_37_48), .A (n_33_50), .B (n_27_53), .C1 (n_30_50), .C2 (n_36_47) );
AOI211_X1 g_39_47 (.ZN (n_39_47), .A (n_35_49), .B (n_29_52), .C1 (n_28_51), .C2 (n_34_48) );
AOI211_X1 g_41_46 (.ZN (n_41_46), .A (n_37_48), .B (n_31_51), .C1 (n_27_53), .C2 (n_32_49) );
AOI211_X1 g_43_45 (.ZN (n_43_45), .A (n_39_47), .B (n_33_50), .C1 (n_29_52), .C2 (n_30_50) );
AOI211_X1 g_45_44 (.ZN (n_45_44), .A (n_41_46), .B (n_35_49), .C1 (n_31_51), .C2 (n_28_51) );
AOI211_X1 g_47_43 (.ZN (n_47_43), .A (n_43_45), .B (n_37_48), .C1 (n_33_50), .C2 (n_27_53) );
AOI211_X1 g_49_42 (.ZN (n_49_42), .A (n_45_44), .B (n_39_47), .C1 (n_35_49), .C2 (n_29_52) );
AOI211_X1 g_51_41 (.ZN (n_51_41), .A (n_47_43), .B (n_41_46), .C1 (n_37_48), .C2 (n_31_51) );
AOI211_X1 g_53_40 (.ZN (n_53_40), .A (n_49_42), .B (n_43_45), .C1 (n_39_47), .C2 (n_33_50) );
AOI211_X1 g_55_39 (.ZN (n_55_39), .A (n_51_41), .B (n_45_44), .C1 (n_41_46), .C2 (n_35_49) );
AOI211_X1 g_57_38 (.ZN (n_57_38), .A (n_53_40), .B (n_47_43), .C1 (n_43_45), .C2 (n_37_48) );
AOI211_X1 g_59_37 (.ZN (n_59_37), .A (n_55_39), .B (n_49_42), .C1 (n_45_44), .C2 (n_39_47) );
AOI211_X1 g_61_36 (.ZN (n_61_36), .A (n_57_38), .B (n_51_41), .C1 (n_47_43), .C2 (n_41_46) );
AOI211_X1 g_60_38 (.ZN (n_60_38), .A (n_59_37), .B (n_53_40), .C1 (n_49_42), .C2 (n_43_45) );
AOI211_X1 g_58_39 (.ZN (n_58_39), .A (n_61_36), .B (n_55_39), .C1 (n_51_41), .C2 (n_45_44) );
AOI211_X1 g_56_40 (.ZN (n_56_40), .A (n_60_38), .B (n_57_38), .C1 (n_53_40), .C2 (n_47_43) );
AOI211_X1 g_54_41 (.ZN (n_54_41), .A (n_58_39), .B (n_59_37), .C1 (n_55_39), .C2 (n_49_42) );
AOI211_X1 g_52_42 (.ZN (n_52_42), .A (n_56_40), .B (n_61_36), .C1 (n_57_38), .C2 (n_51_41) );
AOI211_X1 g_50_43 (.ZN (n_50_43), .A (n_54_41), .B (n_60_38), .C1 (n_59_37), .C2 (n_53_40) );
AOI211_X1 g_48_44 (.ZN (n_48_44), .A (n_52_42), .B (n_58_39), .C1 (n_61_36), .C2 (n_55_39) );
AOI211_X1 g_46_45 (.ZN (n_46_45), .A (n_50_43), .B (n_56_40), .C1 (n_60_38), .C2 (n_57_38) );
AOI211_X1 g_44_46 (.ZN (n_44_46), .A (n_48_44), .B (n_54_41), .C1 (n_58_39), .C2 (n_59_37) );
AOI211_X1 g_42_45 (.ZN (n_42_45), .A (n_46_45), .B (n_52_42), .C1 (n_56_40), .C2 (n_61_36) );
AOI211_X1 g_40_46 (.ZN (n_40_46), .A (n_44_46), .B (n_50_43), .C1 (n_54_41), .C2 (n_60_38) );
AOI211_X1 g_38_47 (.ZN (n_38_47), .A (n_42_45), .B (n_48_44), .C1 (n_52_42), .C2 (n_58_39) );
AOI211_X1 g_36_48 (.ZN (n_36_48), .A (n_40_46), .B (n_46_45), .C1 (n_50_43), .C2 (n_56_40) );
AOI211_X1 g_34_49 (.ZN (n_34_49), .A (n_38_47), .B (n_44_46), .C1 (n_48_44), .C2 (n_54_41) );
AOI211_X1 g_32_50 (.ZN (n_32_50), .A (n_36_48), .B (n_42_45), .C1 (n_46_45), .C2 (n_52_42) );
AOI211_X1 g_30_51 (.ZN (n_30_51), .A (n_34_49), .B (n_40_46), .C1 (n_44_46), .C2 (n_50_43) );
AOI211_X1 g_28_52 (.ZN (n_28_52), .A (n_32_50), .B (n_38_47), .C1 (n_42_45), .C2 (n_48_44) );
AOI211_X1 g_26_53 (.ZN (n_26_53), .A (n_30_51), .B (n_36_48), .C1 (n_40_46), .C2 (n_46_45) );
AOI211_X1 g_24_54 (.ZN (n_24_54), .A (n_28_52), .B (n_34_49), .C1 (n_38_47), .C2 (n_44_46) );
AOI211_X1 g_22_55 (.ZN (n_22_55), .A (n_26_53), .B (n_32_50), .C1 (n_36_48), .C2 (n_42_45) );
AOI211_X1 g_20_56 (.ZN (n_20_56), .A (n_24_54), .B (n_30_51), .C1 (n_34_49), .C2 (n_40_46) );
AOI211_X1 g_18_57 (.ZN (n_18_57), .A (n_22_55), .B (n_28_52), .C1 (n_32_50), .C2 (n_38_47) );
AOI211_X1 g_16_58 (.ZN (n_16_58), .A (n_20_56), .B (n_26_53), .C1 (n_30_51), .C2 (n_36_48) );
AOI211_X1 g_14_59 (.ZN (n_14_59), .A (n_18_57), .B (n_24_54), .C1 (n_28_52), .C2 (n_34_49) );
AOI211_X1 g_12_58 (.ZN (n_12_58), .A (n_16_58), .B (n_22_55), .C1 (n_26_53), .C2 (n_32_50) );
AOI211_X1 g_10_59 (.ZN (n_10_59), .A (n_14_59), .B (n_20_56), .C1 (n_24_54), .C2 (n_30_51) );
AOI211_X1 g_9_61 (.ZN (n_9_61), .A (n_12_58), .B (n_18_57), .C1 (n_22_55), .C2 (n_28_52) );
AOI211_X1 g_11_60 (.ZN (n_11_60), .A (n_10_59), .B (n_16_58), .C1 (n_20_56), .C2 (n_26_53) );
AOI211_X1 g_13_59 (.ZN (n_13_59), .A (n_9_61), .B (n_14_59), .C1 (n_18_57), .C2 (n_24_54) );
AOI211_X1 g_15_58 (.ZN (n_15_58), .A (n_11_60), .B (n_12_58), .C1 (n_16_58), .C2 (n_22_55) );
AOI211_X1 g_17_57 (.ZN (n_17_57), .A (n_13_59), .B (n_10_59), .C1 (n_14_59), .C2 (n_20_56) );
AOI211_X1 g_19_56 (.ZN (n_19_56), .A (n_15_58), .B (n_9_61), .C1 (n_12_58), .C2 (n_18_57) );
AOI211_X1 g_21_55 (.ZN (n_21_55), .A (n_17_57), .B (n_11_60), .C1 (n_10_59), .C2 (n_16_58) );
AOI211_X1 g_20_57 (.ZN (n_20_57), .A (n_19_56), .B (n_13_59), .C1 (n_9_61), .C2 (n_14_59) );
AOI211_X1 g_22_56 (.ZN (n_22_56), .A (n_21_55), .B (n_15_58), .C1 (n_11_60), .C2 (n_12_58) );
AOI211_X1 g_24_55 (.ZN (n_24_55), .A (n_20_57), .B (n_17_57), .C1 (n_13_59), .C2 (n_10_59) );
AOI211_X1 g_26_54 (.ZN (n_26_54), .A (n_22_56), .B (n_19_56), .C1 (n_15_58), .C2 (n_9_61) );
AOI211_X1 g_28_53 (.ZN (n_28_53), .A (n_24_55), .B (n_21_55), .C1 (n_17_57), .C2 (n_11_60) );
AOI211_X1 g_29_51 (.ZN (n_29_51), .A (n_26_54), .B (n_20_57), .C1 (n_19_56), .C2 (n_13_59) );
AOI211_X1 g_31_50 (.ZN (n_31_50), .A (n_28_53), .B (n_22_56), .C1 (n_21_55), .C2 (n_15_58) );
AOI211_X1 g_33_49 (.ZN (n_33_49), .A (n_29_51), .B (n_24_55), .C1 (n_20_57), .C2 (n_17_57) );
AOI211_X1 g_35_48 (.ZN (n_35_48), .A (n_31_50), .B (n_26_54), .C1 (n_22_56), .C2 (n_19_56) );
AOI211_X1 g_34_50 (.ZN (n_34_50), .A (n_33_49), .B (n_28_53), .C1 (n_24_55), .C2 (n_21_55) );
AOI211_X1 g_36_49 (.ZN (n_36_49), .A (n_35_48), .B (n_29_51), .C1 (n_26_54), .C2 (n_20_57) );
AOI211_X1 g_38_48 (.ZN (n_38_48), .A (n_34_50), .B (n_31_50), .C1 (n_28_53), .C2 (n_22_56) );
AOI211_X1 g_40_47 (.ZN (n_40_47), .A (n_36_49), .B (n_33_49), .C1 (n_29_51), .C2 (n_24_55) );
AOI211_X1 g_42_46 (.ZN (n_42_46), .A (n_38_48), .B (n_35_48), .C1 (n_31_50), .C2 (n_26_54) );
AOI211_X1 g_44_45 (.ZN (n_44_45), .A (n_40_47), .B (n_34_50), .C1 (n_33_49), .C2 (n_28_53) );
AOI211_X1 g_46_44 (.ZN (n_46_44), .A (n_42_46), .B (n_36_49), .C1 (n_35_48), .C2 (n_29_51) );
AOI211_X1 g_48_43 (.ZN (n_48_43), .A (n_44_45), .B (n_38_48), .C1 (n_34_50), .C2 (n_31_50) );
AOI211_X1 g_50_42 (.ZN (n_50_42), .A (n_46_44), .B (n_40_47), .C1 (n_36_49), .C2 (n_33_49) );
AOI211_X1 g_52_41 (.ZN (n_52_41), .A (n_48_43), .B (n_42_46), .C1 (n_38_48), .C2 (n_35_48) );
AOI211_X1 g_54_40 (.ZN (n_54_40), .A (n_50_42), .B (n_44_45), .C1 (n_40_47), .C2 (n_34_50) );
AOI211_X1 g_56_39 (.ZN (n_56_39), .A (n_52_41), .B (n_46_44), .C1 (n_42_46), .C2 (n_36_49) );
AOI211_X1 g_58_38 (.ZN (n_58_38), .A (n_54_40), .B (n_48_43), .C1 (n_44_45), .C2 (n_38_48) );
AOI211_X1 g_60_37 (.ZN (n_60_37), .A (n_56_39), .B (n_50_42), .C1 (n_46_44), .C2 (n_40_47) );
AOI211_X1 g_62_36 (.ZN (n_62_36), .A (n_58_38), .B (n_52_41), .C1 (n_48_43), .C2 (n_42_46) );
AOI211_X1 g_64_35 (.ZN (n_64_35), .A (n_60_37), .B (n_54_40), .C1 (n_50_42), .C2 (n_44_45) );
AOI211_X1 g_63_37 (.ZN (n_63_37), .A (n_62_36), .B (n_56_39), .C1 (n_52_41), .C2 (n_46_44) );
AOI211_X1 g_61_38 (.ZN (n_61_38), .A (n_64_35), .B (n_58_38), .C1 (n_54_40), .C2 (n_48_43) );
AOI211_X1 g_59_39 (.ZN (n_59_39), .A (n_63_37), .B (n_60_37), .C1 (n_56_39), .C2 (n_50_42) );
AOI211_X1 g_57_40 (.ZN (n_57_40), .A (n_61_38), .B (n_62_36), .C1 (n_58_38), .C2 (n_52_41) );
AOI211_X1 g_55_41 (.ZN (n_55_41), .A (n_59_39), .B (n_64_35), .C1 (n_60_37), .C2 (n_54_40) );
AOI211_X1 g_53_42 (.ZN (n_53_42), .A (n_57_40), .B (n_63_37), .C1 (n_62_36), .C2 (n_56_39) );
AOI211_X1 g_51_43 (.ZN (n_51_43), .A (n_55_41), .B (n_61_38), .C1 (n_64_35), .C2 (n_58_38) );
AOI211_X1 g_49_44 (.ZN (n_49_44), .A (n_53_42), .B (n_59_39), .C1 (n_63_37), .C2 (n_60_37) );
AOI211_X1 g_47_45 (.ZN (n_47_45), .A (n_51_43), .B (n_57_40), .C1 (n_61_38), .C2 (n_62_36) );
AOI211_X1 g_45_46 (.ZN (n_45_46), .A (n_49_44), .B (n_55_41), .C1 (n_59_39), .C2 (n_64_35) );
AOI211_X1 g_43_47 (.ZN (n_43_47), .A (n_47_45), .B (n_53_42), .C1 (n_57_40), .C2 (n_63_37) );
AOI211_X1 g_41_48 (.ZN (n_41_48), .A (n_45_46), .B (n_51_43), .C1 (n_55_41), .C2 (n_61_38) );
AOI211_X1 g_39_49 (.ZN (n_39_49), .A (n_43_47), .B (n_49_44), .C1 (n_53_42), .C2 (n_59_39) );
AOI211_X1 g_37_50 (.ZN (n_37_50), .A (n_41_48), .B (n_47_45), .C1 (n_51_43), .C2 (n_57_40) );
AOI211_X1 g_35_51 (.ZN (n_35_51), .A (n_39_49), .B (n_45_46), .C1 (n_49_44), .C2 (n_55_41) );
AOI211_X1 g_33_52 (.ZN (n_33_52), .A (n_37_50), .B (n_43_47), .C1 (n_47_45), .C2 (n_53_42) );
AOI211_X1 g_31_53 (.ZN (n_31_53), .A (n_35_51), .B (n_41_48), .C1 (n_45_46), .C2 (n_51_43) );
AOI211_X1 g_32_51 (.ZN (n_32_51), .A (n_33_52), .B (n_39_49), .C1 (n_43_47), .C2 (n_49_44) );
AOI211_X1 g_30_52 (.ZN (n_30_52), .A (n_31_53), .B (n_37_50), .C1 (n_41_48), .C2 (n_47_45) );
AOI211_X1 g_29_54 (.ZN (n_29_54), .A (n_32_51), .B (n_35_51), .C1 (n_39_49), .C2 (n_45_46) );
AOI211_X1 g_27_55 (.ZN (n_27_55), .A (n_30_52), .B (n_33_52), .C1 (n_37_50), .C2 (n_43_47) );
AOI211_X1 g_25_54 (.ZN (n_25_54), .A (n_29_54), .B (n_31_53), .C1 (n_35_51), .C2 (n_41_48) );
AOI211_X1 g_23_55 (.ZN (n_23_55), .A (n_27_55), .B (n_32_51), .C1 (n_33_52), .C2 (n_39_49) );
AOI211_X1 g_21_56 (.ZN (n_21_56), .A (n_25_54), .B (n_30_52), .C1 (n_31_53), .C2 (n_37_50) );
AOI211_X1 g_19_57 (.ZN (n_19_57), .A (n_23_55), .B (n_29_54), .C1 (n_32_51), .C2 (n_35_51) );
AOI211_X1 g_17_58 (.ZN (n_17_58), .A (n_21_56), .B (n_27_55), .C1 (n_30_52), .C2 (n_33_52) );
AOI211_X1 g_16_60 (.ZN (n_16_60), .A (n_19_57), .B (n_25_54), .C1 (n_29_54), .C2 (n_31_53) );
AOI211_X1 g_18_59 (.ZN (n_18_59), .A (n_17_58), .B (n_23_55), .C1 (n_27_55), .C2 (n_32_51) );
AOI211_X1 g_20_58 (.ZN (n_20_58), .A (n_16_60), .B (n_21_56), .C1 (n_25_54), .C2 (n_30_52) );
AOI211_X1 g_22_57 (.ZN (n_22_57), .A (n_18_59), .B (n_19_57), .C1 (n_23_55), .C2 (n_29_54) );
AOI211_X1 g_24_56 (.ZN (n_24_56), .A (n_20_58), .B (n_17_58), .C1 (n_21_56), .C2 (n_27_55) );
AOI211_X1 g_26_55 (.ZN (n_26_55), .A (n_22_57), .B (n_16_60), .C1 (n_19_57), .C2 (n_25_54) );
AOI211_X1 g_28_54 (.ZN (n_28_54), .A (n_24_56), .B (n_18_59), .C1 (n_17_58), .C2 (n_23_55) );
AOI211_X1 g_30_53 (.ZN (n_30_53), .A (n_26_55), .B (n_20_58), .C1 (n_16_60), .C2 (n_21_56) );
AOI211_X1 g_32_52 (.ZN (n_32_52), .A (n_28_54), .B (n_22_57), .C1 (n_18_59), .C2 (n_19_57) );
AOI211_X1 g_34_51 (.ZN (n_34_51), .A (n_30_53), .B (n_24_56), .C1 (n_20_58), .C2 (n_17_58) );
AOI211_X1 g_36_50 (.ZN (n_36_50), .A (n_32_52), .B (n_26_55), .C1 (n_22_57), .C2 (n_16_60) );
AOI211_X1 g_38_49 (.ZN (n_38_49), .A (n_34_51), .B (n_28_54), .C1 (n_24_56), .C2 (n_18_59) );
AOI211_X1 g_40_48 (.ZN (n_40_48), .A (n_36_50), .B (n_30_53), .C1 (n_26_55), .C2 (n_20_58) );
AOI211_X1 g_42_47 (.ZN (n_42_47), .A (n_38_49), .B (n_32_52), .C1 (n_28_54), .C2 (n_22_57) );
AOI211_X1 g_41_49 (.ZN (n_41_49), .A (n_40_48), .B (n_34_51), .C1 (n_30_53), .C2 (n_24_56) );
AOI211_X1 g_39_48 (.ZN (n_39_48), .A (n_42_47), .B (n_36_50), .C1 (n_32_52), .C2 (n_26_55) );
AOI211_X1 g_41_47 (.ZN (n_41_47), .A (n_41_49), .B (n_38_49), .C1 (n_34_51), .C2 (n_28_54) );
AOI211_X1 g_43_46 (.ZN (n_43_46), .A (n_39_48), .B (n_40_48), .C1 (n_36_50), .C2 (n_30_53) );
AOI211_X1 g_45_45 (.ZN (n_45_45), .A (n_41_47), .B (n_42_47), .C1 (n_38_49), .C2 (n_32_52) );
AOI211_X1 g_47_44 (.ZN (n_47_44), .A (n_43_46), .B (n_41_49), .C1 (n_40_48), .C2 (n_34_51) );
AOI211_X1 g_49_43 (.ZN (n_49_43), .A (n_45_45), .B (n_39_48), .C1 (n_42_47), .C2 (n_36_50) );
AOI211_X1 g_51_42 (.ZN (n_51_42), .A (n_47_44), .B (n_41_47), .C1 (n_41_49), .C2 (n_38_49) );
AOI211_X1 g_53_41 (.ZN (n_53_41), .A (n_49_43), .B (n_43_46), .C1 (n_39_48), .C2 (n_40_48) );
AOI211_X1 g_55_40 (.ZN (n_55_40), .A (n_51_42), .B (n_45_45), .C1 (n_41_47), .C2 (n_42_47) );
AOI211_X1 g_57_39 (.ZN (n_57_39), .A (n_53_41), .B (n_47_44), .C1 (n_43_46), .C2 (n_41_49) );
AOI211_X1 g_59_38 (.ZN (n_59_38), .A (n_55_40), .B (n_49_43), .C1 (n_45_45), .C2 (n_39_48) );
AOI211_X1 g_61_37 (.ZN (n_61_37), .A (n_57_39), .B (n_51_42), .C1 (n_47_44), .C2 (n_41_47) );
AOI211_X1 g_60_39 (.ZN (n_60_39), .A (n_59_38), .B (n_53_41), .C1 (n_49_43), .C2 (n_43_46) );
AOI211_X1 g_62_38 (.ZN (n_62_38), .A (n_61_37), .B (n_55_40), .C1 (n_51_42), .C2 (n_45_45) );
AOI211_X1 g_64_37 (.ZN (n_64_37), .A (n_60_39), .B (n_57_39), .C1 (n_53_41), .C2 (n_47_44) );
AOI211_X1 g_66_36 (.ZN (n_66_36), .A (n_62_38), .B (n_59_38), .C1 (n_55_40), .C2 (n_49_43) );
AOI211_X1 g_68_35 (.ZN (n_68_35), .A (n_64_37), .B (n_61_37), .C1 (n_57_39), .C2 (n_51_42) );
AOI211_X1 g_70_34 (.ZN (n_70_34), .A (n_66_36), .B (n_60_39), .C1 (n_59_38), .C2 (n_53_41) );
AOI211_X1 g_69_36 (.ZN (n_69_36), .A (n_68_35), .B (n_62_38), .C1 (n_61_37), .C2 (n_55_40) );
AOI211_X1 g_71_35 (.ZN (n_71_35), .A (n_70_34), .B (n_64_37), .C1 (n_60_39), .C2 (n_57_39) );
AOI211_X1 g_70_37 (.ZN (n_70_37), .A (n_69_36), .B (n_66_36), .C1 (n_62_38), .C2 (n_59_38) );
AOI211_X1 g_69_35 (.ZN (n_69_35), .A (n_71_35), .B (n_68_35), .C1 (n_64_37), .C2 (n_61_37) );
AOI211_X1 g_71_34 (.ZN (n_71_34), .A (n_70_37), .B (n_70_34), .C1 (n_66_36), .C2 (n_60_39) );
AOI211_X1 g_73_33 (.ZN (n_73_33), .A (n_69_35), .B (n_69_36), .C1 (n_68_35), .C2 (n_62_38) );
AOI211_X1 g_75_32 (.ZN (n_75_32), .A (n_71_34), .B (n_71_35), .C1 (n_70_34), .C2 (n_64_37) );
AOI211_X1 g_77_31 (.ZN (n_77_31), .A (n_73_33), .B (n_70_37), .C1 (n_69_36), .C2 (n_66_36) );
AOI211_X1 g_79_30 (.ZN (n_79_30), .A (n_75_32), .B (n_69_35), .C1 (n_71_35), .C2 (n_68_35) );
AOI211_X1 g_81_29 (.ZN (n_81_29), .A (n_77_31), .B (n_71_34), .C1 (n_70_37), .C2 (n_70_34) );
AOI211_X1 g_83_28 (.ZN (n_83_28), .A (n_79_30), .B (n_73_33), .C1 (n_69_35), .C2 (n_69_36) );
AOI211_X1 g_85_27 (.ZN (n_85_27), .A (n_81_29), .B (n_75_32), .C1 (n_71_34), .C2 (n_71_35) );
AOI211_X1 g_87_26 (.ZN (n_87_26), .A (n_83_28), .B (n_77_31), .C1 (n_73_33), .C2 (n_70_37) );
AOI211_X1 g_89_25 (.ZN (n_89_25), .A (n_85_27), .B (n_79_30), .C1 (n_75_32), .C2 (n_69_35) );
AOI211_X1 g_91_24 (.ZN (n_91_24), .A (n_87_26), .B (n_81_29), .C1 (n_77_31), .C2 (n_71_34) );
AOI211_X1 g_93_23 (.ZN (n_93_23), .A (n_89_25), .B (n_83_28), .C1 (n_79_30), .C2 (n_73_33) );
AOI211_X1 g_92_25 (.ZN (n_92_25), .A (n_91_24), .B (n_85_27), .C1 (n_81_29), .C2 (n_75_32) );
AOI211_X1 g_90_26 (.ZN (n_90_26), .A (n_93_23), .B (n_87_26), .C1 (n_83_28), .C2 (n_77_31) );
AOI211_X1 g_88_27 (.ZN (n_88_27), .A (n_92_25), .B (n_89_25), .C1 (n_85_27), .C2 (n_79_30) );
AOI211_X1 g_86_28 (.ZN (n_86_28), .A (n_90_26), .B (n_91_24), .C1 (n_87_26), .C2 (n_81_29) );
AOI211_X1 g_84_29 (.ZN (n_84_29), .A (n_88_27), .B (n_93_23), .C1 (n_89_25), .C2 (n_83_28) );
AOI211_X1 g_82_30 (.ZN (n_82_30), .A (n_86_28), .B (n_92_25), .C1 (n_91_24), .C2 (n_85_27) );
AOI211_X1 g_80_31 (.ZN (n_80_31), .A (n_84_29), .B (n_90_26), .C1 (n_93_23), .C2 (n_87_26) );
AOI211_X1 g_78_32 (.ZN (n_78_32), .A (n_82_30), .B (n_88_27), .C1 (n_92_25), .C2 (n_89_25) );
AOI211_X1 g_76_33 (.ZN (n_76_33), .A (n_80_31), .B (n_86_28), .C1 (n_90_26), .C2 (n_91_24) );
AOI211_X1 g_74_34 (.ZN (n_74_34), .A (n_78_32), .B (n_84_29), .C1 (n_88_27), .C2 (n_93_23) );
AOI211_X1 g_72_35 (.ZN (n_72_35), .A (n_76_33), .B (n_82_30), .C1 (n_86_28), .C2 (n_92_25) );
AOI211_X1 g_70_36 (.ZN (n_70_36), .A (n_74_34), .B (n_80_31), .C1 (n_84_29), .C2 (n_90_26) );
AOI211_X1 g_68_37 (.ZN (n_68_37), .A (n_72_35), .B (n_78_32), .C1 (n_82_30), .C2 (n_88_27) );
AOI211_X1 g_66_38 (.ZN (n_66_38), .A (n_70_36), .B (n_76_33), .C1 (n_80_31), .C2 (n_86_28) );
AOI211_X1 g_67_36 (.ZN (n_67_36), .A (n_68_37), .B (n_74_34), .C1 (n_78_32), .C2 (n_84_29) );
AOI211_X1 g_65_37 (.ZN (n_65_37), .A (n_66_38), .B (n_72_35), .C1 (n_76_33), .C2 (n_82_30) );
AOI211_X1 g_63_38 (.ZN (n_63_38), .A (n_67_36), .B (n_70_36), .C1 (n_74_34), .C2 (n_80_31) );
AOI211_X1 g_61_39 (.ZN (n_61_39), .A (n_65_37), .B (n_68_37), .C1 (n_72_35), .C2 (n_78_32) );
AOI211_X1 g_59_40 (.ZN (n_59_40), .A (n_63_38), .B (n_66_38), .C1 (n_70_36), .C2 (n_76_33) );
AOI211_X1 g_57_41 (.ZN (n_57_41), .A (n_61_39), .B (n_67_36), .C1 (n_68_37), .C2 (n_74_34) );
AOI211_X1 g_55_42 (.ZN (n_55_42), .A (n_59_40), .B (n_65_37), .C1 (n_66_38), .C2 (n_72_35) );
AOI211_X1 g_53_43 (.ZN (n_53_43), .A (n_57_41), .B (n_63_38), .C1 (n_67_36), .C2 (n_70_36) );
AOI211_X1 g_51_44 (.ZN (n_51_44), .A (n_55_42), .B (n_61_39), .C1 (n_65_37), .C2 (n_68_37) );
AOI211_X1 g_49_45 (.ZN (n_49_45), .A (n_53_43), .B (n_59_40), .C1 (n_63_38), .C2 (n_66_38) );
AOI211_X1 g_47_46 (.ZN (n_47_46), .A (n_51_44), .B (n_57_41), .C1 (n_61_39), .C2 (n_67_36) );
AOI211_X1 g_45_47 (.ZN (n_45_47), .A (n_49_45), .B (n_55_42), .C1 (n_59_40), .C2 (n_65_37) );
AOI211_X1 g_43_48 (.ZN (n_43_48), .A (n_47_46), .B (n_53_43), .C1 (n_57_41), .C2 (n_63_38) );
AOI211_X1 g_42_50 (.ZN (n_42_50), .A (n_45_47), .B (n_51_44), .C1 (n_55_42), .C2 (n_61_39) );
AOI211_X1 g_40_49 (.ZN (n_40_49), .A (n_43_48), .B (n_49_45), .C1 (n_53_43), .C2 (n_59_40) );
AOI211_X1 g_42_48 (.ZN (n_42_48), .A (n_42_50), .B (n_47_46), .C1 (n_51_44), .C2 (n_57_41) );
AOI211_X1 g_44_47 (.ZN (n_44_47), .A (n_40_49), .B (n_45_47), .C1 (n_49_45), .C2 (n_55_42) );
AOI211_X1 g_46_46 (.ZN (n_46_46), .A (n_42_48), .B (n_43_48), .C1 (n_47_46), .C2 (n_53_43) );
AOI211_X1 g_48_45 (.ZN (n_48_45), .A (n_44_47), .B (n_42_50), .C1 (n_45_47), .C2 (n_51_44) );
AOI211_X1 g_50_44 (.ZN (n_50_44), .A (n_46_46), .B (n_40_49), .C1 (n_43_48), .C2 (n_49_45) );
AOI211_X1 g_52_43 (.ZN (n_52_43), .A (n_48_45), .B (n_42_48), .C1 (n_42_50), .C2 (n_47_46) );
AOI211_X1 g_54_42 (.ZN (n_54_42), .A (n_50_44), .B (n_44_47), .C1 (n_40_49), .C2 (n_45_47) );
AOI211_X1 g_56_41 (.ZN (n_56_41), .A (n_52_43), .B (n_46_46), .C1 (n_42_48), .C2 (n_43_48) );
AOI211_X1 g_58_40 (.ZN (n_58_40), .A (n_54_42), .B (n_48_45), .C1 (n_44_47), .C2 (n_42_50) );
AOI211_X1 g_57_42 (.ZN (n_57_42), .A (n_56_41), .B (n_50_44), .C1 (n_46_46), .C2 (n_40_49) );
AOI211_X1 g_59_41 (.ZN (n_59_41), .A (n_58_40), .B (n_52_43), .C1 (n_48_45), .C2 (n_42_48) );
AOI211_X1 g_61_40 (.ZN (n_61_40), .A (n_57_42), .B (n_54_42), .C1 (n_50_44), .C2 (n_44_47) );
AOI211_X1 g_63_39 (.ZN (n_63_39), .A (n_59_41), .B (n_56_41), .C1 (n_52_43), .C2 (n_46_46) );
AOI211_X1 g_65_38 (.ZN (n_65_38), .A (n_61_40), .B (n_58_40), .C1 (n_54_42), .C2 (n_48_45) );
AOI211_X1 g_67_37 (.ZN (n_67_37), .A (n_63_39), .B (n_57_42), .C1 (n_56_41), .C2 (n_50_44) );
AOI211_X1 g_66_39 (.ZN (n_66_39), .A (n_65_38), .B (n_59_41), .C1 (n_58_40), .C2 (n_52_43) );
AOI211_X1 g_68_38 (.ZN (n_68_38), .A (n_67_37), .B (n_61_40), .C1 (n_57_42), .C2 (n_54_42) );
AOI211_X1 g_66_37 (.ZN (n_66_37), .A (n_66_39), .B (n_63_39), .C1 (n_59_41), .C2 (n_56_41) );
AOI211_X1 g_68_36 (.ZN (n_68_36), .A (n_68_38), .B (n_65_38), .C1 (n_61_40), .C2 (n_58_40) );
AOI211_X1 g_70_35 (.ZN (n_70_35), .A (n_66_37), .B (n_67_37), .C1 (n_63_39), .C2 (n_57_42) );
AOI211_X1 g_72_34 (.ZN (n_72_34), .A (n_68_36), .B (n_66_39), .C1 (n_65_38), .C2 (n_59_41) );
AOI211_X1 g_74_33 (.ZN (n_74_33), .A (n_70_35), .B (n_68_38), .C1 (n_67_37), .C2 (n_61_40) );
AOI211_X1 g_73_35 (.ZN (n_73_35), .A (n_72_34), .B (n_66_37), .C1 (n_66_39), .C2 (n_63_39) );
AOI211_X1 g_75_34 (.ZN (n_75_34), .A (n_74_33), .B (n_68_36), .C1 (n_68_38), .C2 (n_65_38) );
AOI211_X1 g_74_36 (.ZN (n_74_36), .A (n_73_35), .B (n_70_35), .C1 (n_66_37), .C2 (n_67_37) );
AOI211_X1 g_76_35 (.ZN (n_76_35), .A (n_75_34), .B (n_72_34), .C1 (n_68_36), .C2 (n_66_39) );
AOI211_X1 g_78_34 (.ZN (n_78_34), .A (n_74_36), .B (n_74_33), .C1 (n_70_35), .C2 (n_68_38) );
AOI211_X1 g_79_32 (.ZN (n_79_32), .A (n_76_35), .B (n_73_35), .C1 (n_72_34), .C2 (n_66_37) );
AOI211_X1 g_81_31 (.ZN (n_81_31), .A (n_78_34), .B (n_75_34), .C1 (n_74_33), .C2 (n_68_36) );
AOI211_X1 g_83_30 (.ZN (n_83_30), .A (n_79_32), .B (n_74_36), .C1 (n_73_35), .C2 (n_70_35) );
AOI211_X1 g_85_29 (.ZN (n_85_29), .A (n_81_31), .B (n_76_35), .C1 (n_75_34), .C2 (n_72_34) );
AOI211_X1 g_87_28 (.ZN (n_87_28), .A (n_83_30), .B (n_78_34), .C1 (n_74_36), .C2 (n_74_33) );
AOI211_X1 g_89_27 (.ZN (n_89_27), .A (n_85_29), .B (n_79_32), .C1 (n_76_35), .C2 (n_73_35) );
AOI211_X1 g_91_26 (.ZN (n_91_26), .A (n_87_28), .B (n_81_31), .C1 (n_78_34), .C2 (n_75_34) );
AOI211_X1 g_93_25 (.ZN (n_93_25), .A (n_89_27), .B (n_83_30), .C1 (n_79_32), .C2 (n_74_36) );
AOI211_X1 g_95_24 (.ZN (n_95_24), .A (n_91_26), .B (n_85_29), .C1 (n_81_31), .C2 (n_76_35) );
AOI211_X1 g_94_26 (.ZN (n_94_26), .A (n_93_25), .B (n_87_28), .C1 (n_83_30), .C2 (n_78_34) );
AOI211_X1 g_92_27 (.ZN (n_92_27), .A (n_95_24), .B (n_89_27), .C1 (n_85_29), .C2 (n_79_32) );
AOI211_X1 g_90_28 (.ZN (n_90_28), .A (n_94_26), .B (n_91_26), .C1 (n_87_28), .C2 (n_81_31) );
AOI211_X1 g_88_29 (.ZN (n_88_29), .A (n_92_27), .B (n_93_25), .C1 (n_89_27), .C2 (n_83_30) );
AOI211_X1 g_86_30 (.ZN (n_86_30), .A (n_90_28), .B (n_95_24), .C1 (n_91_26), .C2 (n_85_29) );
AOI211_X1 g_84_31 (.ZN (n_84_31), .A (n_88_29), .B (n_94_26), .C1 (n_93_25), .C2 (n_87_28) );
AOI211_X1 g_82_32 (.ZN (n_82_32), .A (n_86_30), .B (n_92_27), .C1 (n_95_24), .C2 (n_89_27) );
AOI211_X1 g_80_33 (.ZN (n_80_33), .A (n_84_31), .B (n_90_28), .C1 (n_94_26), .C2 (n_91_26) );
AOI211_X1 g_79_35 (.ZN (n_79_35), .A (n_82_32), .B (n_88_29), .C1 (n_92_27), .C2 (n_93_25) );
AOI211_X1 g_78_33 (.ZN (n_78_33), .A (n_80_33), .B (n_86_30), .C1 (n_90_28), .C2 (n_95_24) );
AOI211_X1 g_80_32 (.ZN (n_80_32), .A (n_79_35), .B (n_84_31), .C1 (n_88_29), .C2 (n_94_26) );
AOI211_X1 g_82_31 (.ZN (n_82_31), .A (n_78_33), .B (n_82_32), .C1 (n_86_30), .C2 (n_92_27) );
AOI211_X1 g_84_30 (.ZN (n_84_30), .A (n_80_32), .B (n_80_33), .C1 (n_84_31), .C2 (n_90_28) );
AOI211_X1 g_86_29 (.ZN (n_86_29), .A (n_82_31), .B (n_79_35), .C1 (n_82_32), .C2 (n_88_29) );
AOI211_X1 g_88_28 (.ZN (n_88_28), .A (n_84_30), .B (n_78_33), .C1 (n_80_33), .C2 (n_86_30) );
AOI211_X1 g_90_27 (.ZN (n_90_27), .A (n_86_29), .B (n_80_32), .C1 (n_79_35), .C2 (n_84_31) );
AOI211_X1 g_92_26 (.ZN (n_92_26), .A (n_88_28), .B (n_82_31), .C1 (n_78_33), .C2 (n_82_32) );
AOI211_X1 g_94_25 (.ZN (n_94_25), .A (n_90_27), .B (n_84_30), .C1 (n_80_32), .C2 (n_80_33) );
AOI211_X1 g_96_24 (.ZN (n_96_24), .A (n_92_26), .B (n_86_29), .C1 (n_82_31), .C2 (n_79_35) );
AOI211_X1 g_98_23 (.ZN (n_98_23), .A (n_94_25), .B (n_88_28), .C1 (n_84_30), .C2 (n_78_33) );
AOI211_X1 g_100_24 (.ZN (n_100_24), .A (n_96_24), .B (n_90_27), .C1 (n_86_29), .C2 (n_80_32) );
AOI211_X1 g_98_25 (.ZN (n_98_25), .A (n_98_23), .B (n_92_26), .C1 (n_88_28), .C2 (n_82_31) );
AOI211_X1 g_96_26 (.ZN (n_96_26), .A (n_100_24), .B (n_94_25), .C1 (n_90_27), .C2 (n_84_30) );
AOI211_X1 g_94_27 (.ZN (n_94_27), .A (n_98_25), .B (n_96_24), .C1 (n_92_26), .C2 (n_86_29) );
AOI211_X1 g_92_28 (.ZN (n_92_28), .A (n_96_26), .B (n_98_23), .C1 (n_94_25), .C2 (n_88_28) );
AOI211_X1 g_90_29 (.ZN (n_90_29), .A (n_94_27), .B (n_100_24), .C1 (n_96_24), .C2 (n_90_27) );
AOI211_X1 g_88_30 (.ZN (n_88_30), .A (n_92_28), .B (n_98_25), .C1 (n_98_23), .C2 (n_92_26) );
AOI211_X1 g_89_28 (.ZN (n_89_28), .A (n_90_29), .B (n_96_26), .C1 (n_100_24), .C2 (n_94_25) );
AOI211_X1 g_87_29 (.ZN (n_87_29), .A (n_88_30), .B (n_94_27), .C1 (n_98_25), .C2 (n_96_24) );
AOI211_X1 g_85_30 (.ZN (n_85_30), .A (n_89_28), .B (n_92_28), .C1 (n_96_26), .C2 (n_98_23) );
AOI211_X1 g_83_31 (.ZN (n_83_31), .A (n_87_29), .B (n_90_29), .C1 (n_94_27), .C2 (n_100_24) );
AOI211_X1 g_81_32 (.ZN (n_81_32), .A (n_85_30), .B (n_88_30), .C1 (n_92_28), .C2 (n_98_25) );
AOI211_X1 g_79_33 (.ZN (n_79_33), .A (n_83_31), .B (n_89_28), .C1 (n_90_29), .C2 (n_96_26) );
AOI211_X1 g_77_34 (.ZN (n_77_34), .A (n_81_32), .B (n_87_29), .C1 (n_88_30), .C2 (n_94_27) );
AOI211_X1 g_75_35 (.ZN (n_75_35), .A (n_79_33), .B (n_85_30), .C1 (n_89_28), .C2 (n_92_28) );
AOI211_X1 g_73_36 (.ZN (n_73_36), .A (n_77_34), .B (n_83_31), .C1 (n_87_29), .C2 (n_90_29) );
AOI211_X1 g_71_37 (.ZN (n_71_37), .A (n_75_35), .B (n_81_32), .C1 (n_85_30), .C2 (n_88_30) );
AOI211_X1 g_69_38 (.ZN (n_69_38), .A (n_73_36), .B (n_79_33), .C1 (n_83_31), .C2 (n_89_28) );
AOI211_X1 g_67_39 (.ZN (n_67_39), .A (n_71_37), .B (n_77_34), .C1 (n_81_32), .C2 (n_87_29) );
AOI211_X1 g_65_40 (.ZN (n_65_40), .A (n_69_38), .B (n_75_35), .C1 (n_79_33), .C2 (n_85_30) );
AOI211_X1 g_64_38 (.ZN (n_64_38), .A (n_67_39), .B (n_73_36), .C1 (n_77_34), .C2 (n_83_31) );
AOI211_X1 g_62_39 (.ZN (n_62_39), .A (n_65_40), .B (n_71_37), .C1 (n_75_35), .C2 (n_81_32) );
AOI211_X1 g_60_40 (.ZN (n_60_40), .A (n_64_38), .B (n_69_38), .C1 (n_73_36), .C2 (n_79_33) );
AOI211_X1 g_58_41 (.ZN (n_58_41), .A (n_62_39), .B (n_67_39), .C1 (n_71_37), .C2 (n_77_34) );
AOI211_X1 g_56_42 (.ZN (n_56_42), .A (n_60_40), .B (n_65_40), .C1 (n_69_38), .C2 (n_75_35) );
AOI211_X1 g_54_43 (.ZN (n_54_43), .A (n_58_41), .B (n_64_38), .C1 (n_67_39), .C2 (n_73_36) );
AOI211_X1 g_52_44 (.ZN (n_52_44), .A (n_56_42), .B (n_62_39), .C1 (n_65_40), .C2 (n_71_37) );
AOI211_X1 g_50_45 (.ZN (n_50_45), .A (n_54_43), .B (n_60_40), .C1 (n_64_38), .C2 (n_69_38) );
AOI211_X1 g_48_46 (.ZN (n_48_46), .A (n_52_44), .B (n_58_41), .C1 (n_62_39), .C2 (n_67_39) );
AOI211_X1 g_46_47 (.ZN (n_46_47), .A (n_50_45), .B (n_56_42), .C1 (n_60_40), .C2 (n_65_40) );
AOI211_X1 g_44_48 (.ZN (n_44_48), .A (n_48_46), .B (n_54_43), .C1 (n_58_41), .C2 (n_64_38) );
AOI211_X1 g_42_49 (.ZN (n_42_49), .A (n_46_47), .B (n_52_44), .C1 (n_56_42), .C2 (n_62_39) );
AOI211_X1 g_40_50 (.ZN (n_40_50), .A (n_44_48), .B (n_50_45), .C1 (n_54_43), .C2 (n_60_40) );
AOI211_X1 g_38_51 (.ZN (n_38_51), .A (n_42_49), .B (n_48_46), .C1 (n_52_44), .C2 (n_58_41) );
AOI211_X1 g_37_49 (.ZN (n_37_49), .A (n_40_50), .B (n_46_47), .C1 (n_50_45), .C2 (n_56_42) );
AOI211_X1 g_35_50 (.ZN (n_35_50), .A (n_38_51), .B (n_44_48), .C1 (n_48_46), .C2 (n_54_43) );
AOI211_X1 g_33_51 (.ZN (n_33_51), .A (n_37_49), .B (n_42_49), .C1 (n_46_47), .C2 (n_52_44) );
AOI211_X1 g_31_52 (.ZN (n_31_52), .A (n_35_50), .B (n_40_50), .C1 (n_44_48), .C2 (n_50_45) );
AOI211_X1 g_29_53 (.ZN (n_29_53), .A (n_33_51), .B (n_38_51), .C1 (n_42_49), .C2 (n_48_46) );
AOI211_X1 g_27_54 (.ZN (n_27_54), .A (n_31_52), .B (n_37_49), .C1 (n_40_50), .C2 (n_46_47) );
AOI211_X1 g_25_55 (.ZN (n_25_55), .A (n_29_53), .B (n_35_50), .C1 (n_38_51), .C2 (n_44_48) );
AOI211_X1 g_23_56 (.ZN (n_23_56), .A (n_27_54), .B (n_33_51), .C1 (n_37_49), .C2 (n_42_49) );
AOI211_X1 g_21_57 (.ZN (n_21_57), .A (n_25_55), .B (n_31_52), .C1 (n_35_50), .C2 (n_40_50) );
AOI211_X1 g_19_58 (.ZN (n_19_58), .A (n_23_56), .B (n_29_53), .C1 (n_33_51), .C2 (n_38_51) );
AOI211_X1 g_17_59 (.ZN (n_17_59), .A (n_21_57), .B (n_27_54), .C1 (n_31_52), .C2 (n_37_49) );
AOI211_X1 g_15_60 (.ZN (n_15_60), .A (n_19_58), .B (n_25_55), .C1 (n_29_53), .C2 (n_35_50) );
AOI211_X1 g_13_61 (.ZN (n_13_61), .A (n_17_59), .B (n_23_56), .C1 (n_27_54), .C2 (n_33_51) );
AOI211_X1 g_11_62 (.ZN (n_11_62), .A (n_15_60), .B (n_21_57), .C1 (n_25_55), .C2 (n_31_52) );
AOI211_X1 g_12_60 (.ZN (n_12_60), .A (n_13_61), .B (n_19_58), .C1 (n_23_56), .C2 (n_29_53) );
AOI211_X1 g_10_61 (.ZN (n_10_61), .A (n_11_62), .B (n_17_59), .C1 (n_21_57), .C2 (n_27_54) );
AOI211_X1 g_8_62 (.ZN (n_8_62), .A (n_12_60), .B (n_15_60), .C1 (n_19_58), .C2 (n_25_55) );
AOI211_X1 g_6_63 (.ZN (n_6_63), .A (n_10_61), .B (n_13_61), .C1 (n_17_59), .C2 (n_23_56) );
AOI211_X1 g_7_61 (.ZN (n_7_61), .A (n_8_62), .B (n_11_62), .C1 (n_15_60), .C2 (n_21_57) );
AOI211_X1 g_8_63 (.ZN (n_8_63), .A (n_6_63), .B (n_12_60), .C1 (n_13_61), .C2 (n_19_58) );
AOI211_X1 g_6_62 (.ZN (n_6_62), .A (n_7_61), .B (n_10_61), .C1 (n_11_62), .C2 (n_17_59) );
AOI211_X1 g_8_61 (.ZN (n_8_61), .A (n_8_63), .B (n_8_62), .C1 (n_12_60), .C2 (n_15_60) );
AOI211_X1 g_10_60 (.ZN (n_10_60), .A (n_6_62), .B (n_6_63), .C1 (n_10_61), .C2 (n_13_61) );
AOI211_X1 g_9_62 (.ZN (n_9_62), .A (n_8_61), .B (n_7_61), .C1 (n_8_62), .C2 (n_11_62) );
AOI211_X1 g_11_61 (.ZN (n_11_61), .A (n_10_60), .B (n_8_63), .C1 (n_6_63), .C2 (n_12_60) );
AOI211_X1 g_13_60 (.ZN (n_13_60), .A (n_9_62), .B (n_6_62), .C1 (n_7_61), .C2 (n_10_61) );
AOI211_X1 g_12_62 (.ZN (n_12_62), .A (n_11_61), .B (n_8_61), .C1 (n_8_63), .C2 (n_8_62) );
AOI211_X1 g_14_61 (.ZN (n_14_61), .A (n_13_60), .B (n_10_60), .C1 (n_6_62), .C2 (n_6_63) );
AOI211_X1 g_13_63 (.ZN (n_13_63), .A (n_12_62), .B (n_9_62), .C1 (n_8_61), .C2 (n_7_61) );
AOI211_X1 g_12_61 (.ZN (n_12_61), .A (n_14_61), .B (n_11_61), .C1 (n_10_60), .C2 (n_8_63) );
AOI211_X1 g_10_62 (.ZN (n_10_62), .A (n_13_63), .B (n_13_60), .C1 (n_9_62), .C2 (n_6_62) );
AOI211_X1 g_11_64 (.ZN (n_11_64), .A (n_12_61), .B (n_12_62), .C1 (n_11_61), .C2 (n_8_61) );
AOI211_X1 g_9_63 (.ZN (n_9_63), .A (n_10_62), .B (n_14_61), .C1 (n_13_60), .C2 (n_10_60) );
AOI211_X1 g_7_64 (.ZN (n_7_64), .A (n_11_64), .B (n_13_63), .C1 (n_12_62), .C2 (n_9_62) );
AOI211_X1 g_5_65 (.ZN (n_5_65), .A (n_9_63), .B (n_12_61), .C1 (n_14_61), .C2 (n_11_61) );
AOI211_X1 g_4_67 (.ZN (n_4_67), .A (n_7_64), .B (n_10_62), .C1 (n_13_63), .C2 (n_13_60) );
AOI211_X1 g_6_66 (.ZN (n_6_66), .A (n_5_65), .B (n_11_64), .C1 (n_12_61), .C2 (n_12_62) );
AOI211_X1 g_5_64 (.ZN (n_5_64), .A (n_4_67), .B (n_9_63), .C1 (n_10_62), .C2 (n_14_61) );
AOI211_X1 g_7_63 (.ZN (n_7_63), .A (n_6_66), .B (n_7_64), .C1 (n_11_64), .C2 (n_13_63) );
AOI211_X1 g_8_65 (.ZN (n_8_65), .A (n_5_64), .B (n_5_65), .C1 (n_9_63), .C2 (n_12_61) );
AOI211_X1 g_10_64 (.ZN (n_10_64), .A (n_7_63), .B (n_4_67), .C1 (n_7_64), .C2 (n_10_62) );
AOI211_X1 g_12_63 (.ZN (n_12_63), .A (n_8_65), .B (n_6_66), .C1 (n_5_65), .C2 (n_11_64) );
AOI211_X1 g_14_62 (.ZN (n_14_62), .A (n_10_64), .B (n_5_64), .C1 (n_4_67), .C2 (n_9_63) );
AOI211_X1 g_16_61 (.ZN (n_16_61), .A (n_12_63), .B (n_7_63), .C1 (n_6_66), .C2 (n_7_64) );
AOI211_X1 g_14_60 (.ZN (n_14_60), .A (n_14_62), .B (n_8_65), .C1 (n_5_64), .C2 (n_5_65) );
AOI211_X1 g_16_59 (.ZN (n_16_59), .A (n_16_61), .B (n_10_64), .C1 (n_7_63), .C2 (n_4_67) );
AOI211_X1 g_18_58 (.ZN (n_18_58), .A (n_14_60), .B (n_12_63), .C1 (n_8_65), .C2 (n_6_66) );
AOI211_X1 g_17_60 (.ZN (n_17_60), .A (n_16_59), .B (n_14_62), .C1 (n_10_64), .C2 (n_5_64) );
AOI211_X1 g_19_59 (.ZN (n_19_59), .A (n_18_58), .B (n_16_61), .C1 (n_12_63), .C2 (n_7_63) );
AOI211_X1 g_21_58 (.ZN (n_21_58), .A (n_17_60), .B (n_14_60), .C1 (n_14_62), .C2 (n_8_65) );
AOI211_X1 g_23_57 (.ZN (n_23_57), .A (n_19_59), .B (n_16_59), .C1 (n_16_61), .C2 (n_10_64) );
AOI211_X1 g_25_56 (.ZN (n_25_56), .A (n_21_58), .B (n_18_58), .C1 (n_14_60), .C2 (n_12_63) );
AOI211_X1 g_24_58 (.ZN (n_24_58), .A (n_23_57), .B (n_17_60), .C1 (n_16_59), .C2 (n_14_62) );
AOI211_X1 g_26_57 (.ZN (n_26_57), .A (n_25_56), .B (n_19_59), .C1 (n_18_58), .C2 (n_16_61) );
AOI211_X1 g_28_56 (.ZN (n_28_56), .A (n_24_58), .B (n_21_58), .C1 (n_17_60), .C2 (n_14_60) );
AOI211_X1 g_30_55 (.ZN (n_30_55), .A (n_26_57), .B (n_23_57), .C1 (n_19_59), .C2 (n_16_59) );
AOI211_X1 g_32_54 (.ZN (n_32_54), .A (n_28_56), .B (n_25_56), .C1 (n_21_58), .C2 (n_18_58) );
AOI211_X1 g_34_53 (.ZN (n_34_53), .A (n_30_55), .B (n_24_58), .C1 (n_23_57), .C2 (n_17_60) );
AOI211_X1 g_36_52 (.ZN (n_36_52), .A (n_32_54), .B (n_26_57), .C1 (n_25_56), .C2 (n_19_59) );
AOI211_X1 g_35_54 (.ZN (n_35_54), .A (n_34_53), .B (n_28_56), .C1 (n_24_58), .C2 (n_21_58) );
AOI211_X1 g_34_52 (.ZN (n_34_52), .A (n_36_52), .B (n_30_55), .C1 (n_26_57), .C2 (n_23_57) );
AOI211_X1 g_36_51 (.ZN (n_36_51), .A (n_35_54), .B (n_32_54), .C1 (n_28_56), .C2 (n_25_56) );
AOI211_X1 g_38_50 (.ZN (n_38_50), .A (n_34_52), .B (n_34_53), .C1 (n_30_55), .C2 (n_24_58) );
AOI211_X1 g_40_51 (.ZN (n_40_51), .A (n_36_51), .B (n_36_52), .C1 (n_32_54), .C2 (n_26_57) );
AOI211_X1 g_38_52 (.ZN (n_38_52), .A (n_38_50), .B (n_35_54), .C1 (n_34_53), .C2 (n_28_56) );
AOI211_X1 g_39_50 (.ZN (n_39_50), .A (n_40_51), .B (n_34_52), .C1 (n_36_52), .C2 (n_30_55) );
AOI211_X1 g_37_51 (.ZN (n_37_51), .A (n_38_52), .B (n_36_51), .C1 (n_35_54), .C2 (n_32_54) );
AOI211_X1 g_35_52 (.ZN (n_35_52), .A (n_39_50), .B (n_38_50), .C1 (n_34_52), .C2 (n_34_53) );
AOI211_X1 g_33_53 (.ZN (n_33_53), .A (n_37_51), .B (n_40_51), .C1 (n_36_51), .C2 (n_36_52) );
AOI211_X1 g_31_54 (.ZN (n_31_54), .A (n_35_52), .B (n_38_52), .C1 (n_38_50), .C2 (n_35_54) );
AOI211_X1 g_29_55 (.ZN (n_29_55), .A (n_33_53), .B (n_39_50), .C1 (n_40_51), .C2 (n_34_52) );
AOI211_X1 g_27_56 (.ZN (n_27_56), .A (n_31_54), .B (n_37_51), .C1 (n_38_52), .C2 (n_36_51) );
AOI211_X1 g_25_57 (.ZN (n_25_57), .A (n_29_55), .B (n_35_52), .C1 (n_39_50), .C2 (n_38_50) );
AOI211_X1 g_23_58 (.ZN (n_23_58), .A (n_27_56), .B (n_33_53), .C1 (n_37_51), .C2 (n_40_51) );
AOI211_X1 g_21_59 (.ZN (n_21_59), .A (n_25_57), .B (n_31_54), .C1 (n_35_52), .C2 (n_38_52) );
AOI211_X1 g_19_60 (.ZN (n_19_60), .A (n_23_58), .B (n_29_55), .C1 (n_33_53), .C2 (n_39_50) );
AOI211_X1 g_17_61 (.ZN (n_17_61), .A (n_21_59), .B (n_27_56), .C1 (n_31_54), .C2 (n_37_51) );
AOI211_X1 g_15_62 (.ZN (n_15_62), .A (n_19_60), .B (n_25_57), .C1 (n_29_55), .C2 (n_35_52) );
AOI211_X1 g_14_64 (.ZN (n_14_64), .A (n_17_61), .B (n_23_58), .C1 (n_27_56), .C2 (n_33_53) );
AOI211_X1 g_13_62 (.ZN (n_13_62), .A (n_15_62), .B (n_21_59), .C1 (n_25_57), .C2 (n_31_54) );
AOI211_X1 g_15_61 (.ZN (n_15_61), .A (n_14_64), .B (n_19_60), .C1 (n_23_58), .C2 (n_29_55) );
AOI211_X1 g_16_63 (.ZN (n_16_63), .A (n_13_62), .B (n_17_61), .C1 (n_21_59), .C2 (n_27_56) );
AOI211_X1 g_18_62 (.ZN (n_18_62), .A (n_15_61), .B (n_15_62), .C1 (n_19_60), .C2 (n_25_57) );
AOI211_X1 g_20_61 (.ZN (n_20_61), .A (n_16_63), .B (n_14_64), .C1 (n_17_61), .C2 (n_23_58) );
AOI211_X1 g_18_60 (.ZN (n_18_60), .A (n_18_62), .B (n_13_62), .C1 (n_15_62), .C2 (n_21_59) );
AOI211_X1 g_20_59 (.ZN (n_20_59), .A (n_20_61), .B (n_15_61), .C1 (n_14_64), .C2 (n_19_60) );
AOI211_X1 g_22_58 (.ZN (n_22_58), .A (n_18_60), .B (n_16_63), .C1 (n_13_62), .C2 (n_17_61) );
AOI211_X1 g_24_57 (.ZN (n_24_57), .A (n_20_59), .B (n_18_62), .C1 (n_15_61), .C2 (n_15_62) );
AOI211_X1 g_26_56 (.ZN (n_26_56), .A (n_22_58), .B (n_20_61), .C1 (n_16_63), .C2 (n_14_64) );
AOI211_X1 g_28_55 (.ZN (n_28_55), .A (n_24_57), .B (n_18_60), .C1 (n_18_62), .C2 (n_13_62) );
AOI211_X1 g_30_54 (.ZN (n_30_54), .A (n_26_56), .B (n_20_59), .C1 (n_20_61), .C2 (n_15_61) );
AOI211_X1 g_32_53 (.ZN (n_32_53), .A (n_28_55), .B (n_22_58), .C1 (n_18_60), .C2 (n_16_63) );
AOI211_X1 g_33_55 (.ZN (n_33_55), .A (n_30_54), .B (n_24_57), .C1 (n_20_59), .C2 (n_18_62) );
AOI211_X1 g_31_56 (.ZN (n_31_56), .A (n_32_53), .B (n_26_56), .C1 (n_22_58), .C2 (n_20_61) );
AOI211_X1 g_29_57 (.ZN (n_29_57), .A (n_33_55), .B (n_28_55), .C1 (n_24_57), .C2 (n_18_60) );
AOI211_X1 g_27_58 (.ZN (n_27_58), .A (n_31_56), .B (n_30_54), .C1 (n_26_56), .C2 (n_20_59) );
AOI211_X1 g_25_59 (.ZN (n_25_59), .A (n_29_57), .B (n_32_53), .C1 (n_28_55), .C2 (n_22_58) );
AOI211_X1 g_23_60 (.ZN (n_23_60), .A (n_27_58), .B (n_33_55), .C1 (n_30_54), .C2 (n_24_57) );
AOI211_X1 g_21_61 (.ZN (n_21_61), .A (n_25_59), .B (n_31_56), .C1 (n_32_53), .C2 (n_26_56) );
AOI211_X1 g_22_59 (.ZN (n_22_59), .A (n_23_60), .B (n_29_57), .C1 (n_33_55), .C2 (n_28_55) );
AOI211_X1 g_20_60 (.ZN (n_20_60), .A (n_21_61), .B (n_27_58), .C1 (n_31_56), .C2 (n_30_54) );
AOI211_X1 g_18_61 (.ZN (n_18_61), .A (n_22_59), .B (n_25_59), .C1 (n_29_57), .C2 (n_32_53) );
AOI211_X1 g_16_62 (.ZN (n_16_62), .A (n_20_60), .B (n_23_60), .C1 (n_27_58), .C2 (n_33_55) );
AOI211_X1 g_14_63 (.ZN (n_14_63), .A (n_18_61), .B (n_21_61), .C1 (n_25_59), .C2 (n_31_56) );
AOI211_X1 g_12_64 (.ZN (n_12_64), .A (n_16_62), .B (n_22_59), .C1 (n_23_60), .C2 (n_29_57) );
AOI211_X1 g_10_63 (.ZN (n_10_63), .A (n_14_63), .B (n_20_60), .C1 (n_21_61), .C2 (n_27_58) );
AOI211_X1 g_8_64 (.ZN (n_8_64), .A (n_12_64), .B (n_18_61), .C1 (n_22_59), .C2 (n_25_59) );
AOI211_X1 g_6_65 (.ZN (n_6_65), .A (n_10_63), .B (n_16_62), .C1 (n_20_60), .C2 (n_23_60) );
AOI211_X1 g_4_66 (.ZN (n_4_66), .A (n_8_64), .B (n_14_63), .C1 (n_18_61), .C2 (n_21_61) );
AOI211_X1 g_3_68 (.ZN (n_3_68), .A (n_6_65), .B (n_12_64), .C1 (n_16_62), .C2 (n_22_59) );
AOI211_X1 g_2_70 (.ZN (n_2_70), .A (n_4_66), .B (n_10_63), .C1 (n_14_63), .C2 (n_20_60) );
AOI211_X1 g_4_69 (.ZN (n_4_69), .A (n_3_68), .B (n_8_64), .C1 (n_12_64), .C2 (n_18_61) );
AOI211_X1 g_5_67 (.ZN (n_5_67), .A (n_2_70), .B (n_6_65), .C1 (n_10_63), .C2 (n_16_62) );
AOI211_X1 g_7_66 (.ZN (n_7_66), .A (n_4_69), .B (n_4_66), .C1 (n_8_64), .C2 (n_14_63) );
AOI211_X1 g_9_65 (.ZN (n_9_65), .A (n_5_67), .B (n_3_68), .C1 (n_6_65), .C2 (n_12_64) );
AOI211_X1 g_11_66 (.ZN (n_11_66), .A (n_7_66), .B (n_2_70), .C1 (n_4_66), .C2 (n_10_63) );
AOI211_X1 g_13_65 (.ZN (n_13_65), .A (n_9_65), .B (n_4_69), .C1 (n_3_68), .C2 (n_8_64) );
AOI211_X1 g_15_64 (.ZN (n_15_64), .A (n_11_66), .B (n_5_67), .C1 (n_2_70), .C2 (n_6_65) );
AOI211_X1 g_17_63 (.ZN (n_17_63), .A (n_13_65), .B (n_7_66), .C1 (n_4_69), .C2 (n_4_66) );
AOI211_X1 g_19_62 (.ZN (n_19_62), .A (n_15_64), .B (n_9_65), .C1 (n_5_67), .C2 (n_3_68) );
AOI211_X1 g_18_64 (.ZN (n_18_64), .A (n_17_63), .B (n_11_66), .C1 (n_7_66), .C2 (n_2_70) );
AOI211_X1 g_17_62 (.ZN (n_17_62), .A (n_19_62), .B (n_13_65), .C1 (n_9_65), .C2 (n_4_69) );
AOI211_X1 g_19_61 (.ZN (n_19_61), .A (n_18_64), .B (n_15_64), .C1 (n_11_66), .C2 (n_5_67) );
AOI211_X1 g_21_60 (.ZN (n_21_60), .A (n_17_62), .B (n_17_63), .C1 (n_13_65), .C2 (n_7_66) );
AOI211_X1 g_23_59 (.ZN (n_23_59), .A (n_19_61), .B (n_19_62), .C1 (n_15_64), .C2 (n_9_65) );
AOI211_X1 g_25_58 (.ZN (n_25_58), .A (n_21_60), .B (n_18_64), .C1 (n_17_63), .C2 (n_11_66) );
AOI211_X1 g_27_57 (.ZN (n_27_57), .A (n_23_59), .B (n_17_62), .C1 (n_19_62), .C2 (n_13_65) );
AOI211_X1 g_29_56 (.ZN (n_29_56), .A (n_25_58), .B (n_19_61), .C1 (n_18_64), .C2 (n_15_64) );
AOI211_X1 g_31_55 (.ZN (n_31_55), .A (n_27_57), .B (n_21_60), .C1 (n_17_62), .C2 (n_17_63) );
AOI211_X1 g_33_54 (.ZN (n_33_54), .A (n_29_56), .B (n_23_59), .C1 (n_19_61), .C2 (n_19_62) );
AOI211_X1 g_35_53 (.ZN (n_35_53), .A (n_31_55), .B (n_25_58), .C1 (n_21_60), .C2 (n_18_64) );
AOI211_X1 g_37_52 (.ZN (n_37_52), .A (n_33_54), .B (n_27_57), .C1 (n_23_59), .C2 (n_17_62) );
AOI211_X1 g_39_51 (.ZN (n_39_51), .A (n_35_53), .B (n_29_56), .C1 (n_25_58), .C2 (n_19_61) );
AOI211_X1 g_41_50 (.ZN (n_41_50), .A (n_37_52), .B (n_31_55), .C1 (n_27_57), .C2 (n_21_60) );
AOI211_X1 g_43_49 (.ZN (n_43_49), .A (n_39_51), .B (n_33_54), .C1 (n_29_56), .C2 (n_23_59) );
AOI211_X1 g_45_48 (.ZN (n_45_48), .A (n_41_50), .B (n_35_53), .C1 (n_31_55), .C2 (n_25_58) );
AOI211_X1 g_47_47 (.ZN (n_47_47), .A (n_43_49), .B (n_37_52), .C1 (n_33_54), .C2 (n_27_57) );
AOI211_X1 g_49_46 (.ZN (n_49_46), .A (n_45_48), .B (n_39_51), .C1 (n_35_53), .C2 (n_29_56) );
AOI211_X1 g_51_45 (.ZN (n_51_45), .A (n_47_47), .B (n_41_50), .C1 (n_37_52), .C2 (n_31_55) );
AOI211_X1 g_53_44 (.ZN (n_53_44), .A (n_49_46), .B (n_43_49), .C1 (n_39_51), .C2 (n_33_54) );
AOI211_X1 g_55_43 (.ZN (n_55_43), .A (n_51_45), .B (n_45_48), .C1 (n_41_50), .C2 (n_35_53) );
AOI211_X1 g_54_45 (.ZN (n_54_45), .A (n_53_44), .B (n_47_47), .C1 (n_43_49), .C2 (n_37_52) );
AOI211_X1 g_56_44 (.ZN (n_56_44), .A (n_55_43), .B (n_49_46), .C1 (n_45_48), .C2 (n_39_51) );
AOI211_X1 g_58_43 (.ZN (n_58_43), .A (n_54_45), .B (n_51_45), .C1 (n_47_47), .C2 (n_41_50) );
AOI211_X1 g_60_42 (.ZN (n_60_42), .A (n_56_44), .B (n_53_44), .C1 (n_49_46), .C2 (n_43_49) );
AOI211_X1 g_62_41 (.ZN (n_62_41), .A (n_58_43), .B (n_55_43), .C1 (n_51_45), .C2 (n_45_48) );
AOI211_X1 g_64_40 (.ZN (n_64_40), .A (n_60_42), .B (n_54_45), .C1 (n_53_44), .C2 (n_47_47) );
AOI211_X1 g_66_41 (.ZN (n_66_41), .A (n_62_41), .B (n_56_44), .C1 (n_55_43), .C2 (n_49_46) );
AOI211_X1 g_65_39 (.ZN (n_65_39), .A (n_64_40), .B (n_58_43), .C1 (n_54_45), .C2 (n_51_45) );
AOI211_X1 g_67_38 (.ZN (n_67_38), .A (n_66_41), .B (n_60_42), .C1 (n_56_44), .C2 (n_53_44) );
AOI211_X1 g_69_37 (.ZN (n_69_37), .A (n_65_39), .B (n_62_41), .C1 (n_58_43), .C2 (n_55_43) );
AOI211_X1 g_71_36 (.ZN (n_71_36), .A (n_67_38), .B (n_64_40), .C1 (n_60_42), .C2 (n_54_45) );
AOI211_X1 g_70_38 (.ZN (n_70_38), .A (n_69_37), .B (n_66_41), .C1 (n_62_41), .C2 (n_56_44) );
AOI211_X1 g_72_37 (.ZN (n_72_37), .A (n_71_36), .B (n_65_39), .C1 (n_64_40), .C2 (n_58_43) );
AOI211_X1 g_71_39 (.ZN (n_71_39), .A (n_70_38), .B (n_67_38), .C1 (n_66_41), .C2 (n_60_42) );
AOI211_X1 g_69_40 (.ZN (n_69_40), .A (n_72_37), .B (n_69_37), .C1 (n_65_39), .C2 (n_62_41) );
AOI211_X1 g_67_41 (.ZN (n_67_41), .A (n_71_39), .B (n_71_36), .C1 (n_67_38), .C2 (n_64_40) );
AOI211_X1 g_68_39 (.ZN (n_68_39), .A (n_69_40), .B (n_70_38), .C1 (n_69_37), .C2 (n_66_41) );
AOI211_X1 g_66_40 (.ZN (n_66_40), .A (n_67_41), .B (n_72_37), .C1 (n_71_36), .C2 (n_65_39) );
AOI211_X1 g_64_39 (.ZN (n_64_39), .A (n_68_39), .B (n_71_39), .C1 (n_70_38), .C2 (n_67_38) );
AOI211_X1 g_62_40 (.ZN (n_62_40), .A (n_66_40), .B (n_69_40), .C1 (n_72_37), .C2 (n_69_37) );
AOI211_X1 g_60_41 (.ZN (n_60_41), .A (n_64_39), .B (n_67_41), .C1 (n_71_39), .C2 (n_71_36) );
AOI211_X1 g_58_42 (.ZN (n_58_42), .A (n_62_40), .B (n_68_39), .C1 (n_69_40), .C2 (n_70_38) );
AOI211_X1 g_56_43 (.ZN (n_56_43), .A (n_60_41), .B (n_66_40), .C1 (n_67_41), .C2 (n_72_37) );
AOI211_X1 g_54_44 (.ZN (n_54_44), .A (n_58_42), .B (n_64_39), .C1 (n_68_39), .C2 (n_71_39) );
AOI211_X1 g_52_45 (.ZN (n_52_45), .A (n_56_43), .B (n_62_40), .C1 (n_66_40), .C2 (n_69_40) );
AOI211_X1 g_50_46 (.ZN (n_50_46), .A (n_54_44), .B (n_60_41), .C1 (n_64_39), .C2 (n_67_41) );
AOI211_X1 g_48_47 (.ZN (n_48_47), .A (n_52_45), .B (n_58_42), .C1 (n_62_40), .C2 (n_68_39) );
AOI211_X1 g_46_48 (.ZN (n_46_48), .A (n_50_46), .B (n_56_43), .C1 (n_60_41), .C2 (n_66_40) );
AOI211_X1 g_44_49 (.ZN (n_44_49), .A (n_48_47), .B (n_54_44), .C1 (n_58_42), .C2 (n_64_39) );
AOI211_X1 g_43_51 (.ZN (n_43_51), .A (n_46_48), .B (n_52_45), .C1 (n_56_43), .C2 (n_62_40) );
AOI211_X1 g_45_50 (.ZN (n_45_50), .A (n_44_49), .B (n_50_46), .C1 (n_54_44), .C2 (n_60_41) );
AOI211_X1 g_47_49 (.ZN (n_47_49), .A (n_43_51), .B (n_48_47), .C1 (n_52_45), .C2 (n_58_42) );
AOI211_X1 g_49_48 (.ZN (n_49_48), .A (n_45_50), .B (n_46_48), .C1 (n_50_46), .C2 (n_56_43) );
AOI211_X1 g_51_47 (.ZN (n_51_47), .A (n_47_49), .B (n_44_49), .C1 (n_48_47), .C2 (n_54_44) );
AOI211_X1 g_53_46 (.ZN (n_53_46), .A (n_49_48), .B (n_43_51), .C1 (n_46_48), .C2 (n_52_45) );
AOI211_X1 g_55_45 (.ZN (n_55_45), .A (n_51_47), .B (n_45_50), .C1 (n_44_49), .C2 (n_50_46) );
AOI211_X1 g_57_44 (.ZN (n_57_44), .A (n_53_46), .B (n_47_49), .C1 (n_43_51), .C2 (n_48_47) );
AOI211_X1 g_59_43 (.ZN (n_59_43), .A (n_55_45), .B (n_49_48), .C1 (n_45_50), .C2 (n_46_48) );
AOI211_X1 g_61_42 (.ZN (n_61_42), .A (n_57_44), .B (n_51_47), .C1 (n_47_49), .C2 (n_44_49) );
AOI211_X1 g_63_41 (.ZN (n_63_41), .A (n_59_43), .B (n_53_46), .C1 (n_49_48), .C2 (n_43_51) );
AOI211_X1 g_65_42 (.ZN (n_65_42), .A (n_61_42), .B (n_55_45), .C1 (n_51_47), .C2 (n_45_50) );
AOI211_X1 g_63_43 (.ZN (n_63_43), .A (n_63_41), .B (n_57_44), .C1 (n_53_46), .C2 (n_47_49) );
AOI211_X1 g_64_41 (.ZN (n_64_41), .A (n_65_42), .B (n_59_43), .C1 (n_55_45), .C2 (n_49_48) );
AOI211_X1 g_62_42 (.ZN (n_62_42), .A (n_63_43), .B (n_61_42), .C1 (n_57_44), .C2 (n_51_47) );
AOI211_X1 g_63_40 (.ZN (n_63_40), .A (n_64_41), .B (n_63_41), .C1 (n_59_43), .C2 (n_53_46) );
AOI211_X1 g_61_41 (.ZN (n_61_41), .A (n_62_42), .B (n_65_42), .C1 (n_61_42), .C2 (n_55_45) );
AOI211_X1 g_59_42 (.ZN (n_59_42), .A (n_63_40), .B (n_63_43), .C1 (n_63_41), .C2 (n_57_44) );
AOI211_X1 g_57_43 (.ZN (n_57_43), .A (n_61_41), .B (n_64_41), .C1 (n_65_42), .C2 (n_59_43) );
AOI211_X1 g_55_44 (.ZN (n_55_44), .A (n_59_42), .B (n_62_42), .C1 (n_63_43), .C2 (n_61_42) );
AOI211_X1 g_53_45 (.ZN (n_53_45), .A (n_57_43), .B (n_63_40), .C1 (n_64_41), .C2 (n_63_41) );
AOI211_X1 g_51_46 (.ZN (n_51_46), .A (n_55_44), .B (n_61_41), .C1 (n_62_42), .C2 (n_65_42) );
AOI211_X1 g_49_47 (.ZN (n_49_47), .A (n_53_45), .B (n_59_42), .C1 (n_63_40), .C2 (n_63_43) );
AOI211_X1 g_47_48 (.ZN (n_47_48), .A (n_51_46), .B (n_57_43), .C1 (n_61_41), .C2 (n_64_41) );
AOI211_X1 g_45_49 (.ZN (n_45_49), .A (n_49_47), .B (n_55_44), .C1 (n_59_42), .C2 (n_62_42) );
AOI211_X1 g_43_50 (.ZN (n_43_50), .A (n_47_48), .B (n_53_45), .C1 (n_57_43), .C2 (n_63_40) );
AOI211_X1 g_41_51 (.ZN (n_41_51), .A (n_45_49), .B (n_51_46), .C1 (n_55_44), .C2 (n_61_41) );
AOI211_X1 g_39_52 (.ZN (n_39_52), .A (n_43_50), .B (n_49_47), .C1 (n_53_45), .C2 (n_59_42) );
AOI211_X1 g_37_53 (.ZN (n_37_53), .A (n_41_51), .B (n_47_48), .C1 (n_51_46), .C2 (n_57_43) );
AOI211_X1 g_36_55 (.ZN (n_36_55), .A (n_39_52), .B (n_45_49), .C1 (n_49_47), .C2 (n_55_44) );
AOI211_X1 g_34_54 (.ZN (n_34_54), .A (n_37_53), .B (n_43_50), .C1 (n_47_48), .C2 (n_53_45) );
AOI211_X1 g_36_53 (.ZN (n_36_53), .A (n_36_55), .B (n_41_51), .C1 (n_45_49), .C2 (n_51_46) );
AOI211_X1 g_38_54 (.ZN (n_38_54), .A (n_34_54), .B (n_39_52), .C1 (n_43_50), .C2 (n_49_47) );
AOI211_X1 g_40_53 (.ZN (n_40_53), .A (n_36_53), .B (n_37_53), .C1 (n_41_51), .C2 (n_47_48) );
AOI211_X1 g_42_52 (.ZN (n_42_52), .A (n_38_54), .B (n_36_55), .C1 (n_39_52), .C2 (n_45_49) );
AOI211_X1 g_44_51 (.ZN (n_44_51), .A (n_40_53), .B (n_34_54), .C1 (n_37_53), .C2 (n_43_50) );
AOI211_X1 g_46_50 (.ZN (n_46_50), .A (n_42_52), .B (n_36_53), .C1 (n_36_55), .C2 (n_41_51) );
AOI211_X1 g_48_49 (.ZN (n_48_49), .A (n_44_51), .B (n_38_54), .C1 (n_34_54), .C2 (n_39_52) );
AOI211_X1 g_50_48 (.ZN (n_50_48), .A (n_46_50), .B (n_40_53), .C1 (n_36_53), .C2 (n_37_53) );
AOI211_X1 g_52_47 (.ZN (n_52_47), .A (n_48_49), .B (n_42_52), .C1 (n_38_54), .C2 (n_36_55) );
AOI211_X1 g_54_46 (.ZN (n_54_46), .A (n_50_48), .B (n_44_51), .C1 (n_40_53), .C2 (n_34_54) );
AOI211_X1 g_56_45 (.ZN (n_56_45), .A (n_52_47), .B (n_46_50), .C1 (n_42_52), .C2 (n_36_53) );
AOI211_X1 g_58_44 (.ZN (n_58_44), .A (n_54_46), .B (n_48_49), .C1 (n_44_51), .C2 (n_38_54) );
AOI211_X1 g_60_43 (.ZN (n_60_43), .A (n_56_45), .B (n_50_48), .C1 (n_46_50), .C2 (n_40_53) );
AOI211_X1 g_59_45 (.ZN (n_59_45), .A (n_58_44), .B (n_52_47), .C1 (n_48_49), .C2 (n_42_52) );
AOI211_X1 g_61_44 (.ZN (n_61_44), .A (n_60_43), .B (n_54_46), .C1 (n_50_48), .C2 (n_44_51) );
AOI211_X1 g_60_46 (.ZN (n_60_46), .A (n_59_45), .B (n_56_45), .C1 (n_52_47), .C2 (n_46_50) );
AOI211_X1 g_59_44 (.ZN (n_59_44), .A (n_61_44), .B (n_58_44), .C1 (n_54_46), .C2 (n_48_49) );
AOI211_X1 g_61_43 (.ZN (n_61_43), .A (n_60_46), .B (n_60_43), .C1 (n_56_45), .C2 (n_50_48) );
AOI211_X1 g_63_42 (.ZN (n_63_42), .A (n_59_44), .B (n_59_45), .C1 (n_58_44), .C2 (n_52_47) );
AOI211_X1 g_65_41 (.ZN (n_65_41), .A (n_61_43), .B (n_61_44), .C1 (n_60_43), .C2 (n_54_46) );
AOI211_X1 g_67_40 (.ZN (n_67_40), .A (n_63_42), .B (n_60_46), .C1 (n_59_45), .C2 (n_56_45) );
AOI211_X1 g_69_39 (.ZN (n_69_39), .A (n_65_41), .B (n_59_44), .C1 (n_61_44), .C2 (n_58_44) );
AOI211_X1 g_71_38 (.ZN (n_71_38), .A (n_67_40), .B (n_61_43), .C1 (n_60_46), .C2 (n_60_43) );
AOI211_X1 g_72_36 (.ZN (n_72_36), .A (n_69_39), .B (n_63_42), .C1 (n_59_44), .C2 (n_59_45) );
AOI211_X1 g_74_35 (.ZN (n_74_35), .A (n_71_38), .B (n_65_41), .C1 (n_61_43), .C2 (n_61_44) );
AOI211_X1 g_76_34 (.ZN (n_76_34), .A (n_72_36), .B (n_67_40), .C1 (n_63_42), .C2 (n_60_46) );
AOI211_X1 g_77_36 (.ZN (n_77_36), .A (n_74_35), .B (n_69_39), .C1 (n_65_41), .C2 (n_59_44) );
AOI211_X1 g_75_37 (.ZN (n_75_37), .A (n_76_34), .B (n_71_38), .C1 (n_67_40), .C2 (n_61_43) );
AOI211_X1 g_73_38 (.ZN (n_73_38), .A (n_77_36), .B (n_72_36), .C1 (n_69_39), .C2 (n_63_42) );
AOI211_X1 g_72_40 (.ZN (n_72_40), .A (n_75_37), .B (n_74_35), .C1 (n_71_38), .C2 (n_65_41) );
AOI211_X1 g_70_39 (.ZN (n_70_39), .A (n_73_38), .B (n_76_34), .C1 (n_72_36), .C2 (n_67_40) );
AOI211_X1 g_68_40 (.ZN (n_68_40), .A (n_72_40), .B (n_77_36), .C1 (n_74_35), .C2 (n_69_39) );
AOI211_X1 g_70_41 (.ZN (n_70_41), .A (n_70_39), .B (n_75_37), .C1 (n_76_34), .C2 (n_71_38) );
AOI211_X1 g_68_42 (.ZN (n_68_42), .A (n_68_40), .B (n_73_38), .C1 (n_77_36), .C2 (n_72_36) );
AOI211_X1 g_66_43 (.ZN (n_66_43), .A (n_70_41), .B (n_72_40), .C1 (n_75_37), .C2 (n_74_35) );
AOI211_X1 g_64_42 (.ZN (n_64_42), .A (n_68_42), .B (n_70_39), .C1 (n_73_38), .C2 (n_76_34) );
AOI211_X1 g_62_43 (.ZN (n_62_43), .A (n_66_43), .B (n_68_40), .C1 (n_72_40), .C2 (n_77_36) );
AOI211_X1 g_60_44 (.ZN (n_60_44), .A (n_64_42), .B (n_70_41), .C1 (n_70_39), .C2 (n_75_37) );
AOI211_X1 g_58_45 (.ZN (n_58_45), .A (n_62_43), .B (n_68_42), .C1 (n_68_40), .C2 (n_73_38) );
AOI211_X1 g_56_46 (.ZN (n_56_46), .A (n_60_44), .B (n_66_43), .C1 (n_70_41), .C2 (n_72_40) );
AOI211_X1 g_54_47 (.ZN (n_54_47), .A (n_58_45), .B (n_64_42), .C1 (n_68_42), .C2 (n_70_39) );
AOI211_X1 g_52_46 (.ZN (n_52_46), .A (n_56_46), .B (n_62_43), .C1 (n_66_43), .C2 (n_68_40) );
AOI211_X1 g_50_47 (.ZN (n_50_47), .A (n_54_47), .B (n_60_44), .C1 (n_64_42), .C2 (n_70_41) );
AOI211_X1 g_48_48 (.ZN (n_48_48), .A (n_52_46), .B (n_58_45), .C1 (n_62_43), .C2 (n_68_42) );
AOI211_X1 g_46_49 (.ZN (n_46_49), .A (n_50_47), .B (n_56_46), .C1 (n_60_44), .C2 (n_66_43) );
AOI211_X1 g_44_50 (.ZN (n_44_50), .A (n_48_48), .B (n_54_47), .C1 (n_58_45), .C2 (n_64_42) );
AOI211_X1 g_42_51 (.ZN (n_42_51), .A (n_46_49), .B (n_52_46), .C1 (n_56_46), .C2 (n_62_43) );
AOI211_X1 g_40_52 (.ZN (n_40_52), .A (n_44_50), .B (n_50_47), .C1 (n_54_47), .C2 (n_60_44) );
AOI211_X1 g_38_53 (.ZN (n_38_53), .A (n_42_51), .B (n_48_48), .C1 (n_52_46), .C2 (n_58_45) );
AOI211_X1 g_36_54 (.ZN (n_36_54), .A (n_40_52), .B (n_46_49), .C1 (n_50_47), .C2 (n_56_46) );
AOI211_X1 g_34_55 (.ZN (n_34_55), .A (n_38_53), .B (n_44_50), .C1 (n_48_48), .C2 (n_54_47) );
AOI211_X1 g_32_56 (.ZN (n_32_56), .A (n_36_54), .B (n_42_51), .C1 (n_46_49), .C2 (n_52_46) );
AOI211_X1 g_30_57 (.ZN (n_30_57), .A (n_34_55), .B (n_40_52), .C1 (n_44_50), .C2 (n_50_47) );
AOI211_X1 g_28_58 (.ZN (n_28_58), .A (n_32_56), .B (n_38_53), .C1 (n_42_51), .C2 (n_48_48) );
AOI211_X1 g_26_59 (.ZN (n_26_59), .A (n_30_57), .B (n_36_54), .C1 (n_40_52), .C2 (n_46_49) );
AOI211_X1 g_24_60 (.ZN (n_24_60), .A (n_28_58), .B (n_34_55), .C1 (n_38_53), .C2 (n_44_50) );
AOI211_X1 g_22_61 (.ZN (n_22_61), .A (n_26_59), .B (n_32_56), .C1 (n_36_54), .C2 (n_42_51) );
AOI211_X1 g_20_62 (.ZN (n_20_62), .A (n_24_60), .B (n_30_57), .C1 (n_34_55), .C2 (n_40_52) );
AOI211_X1 g_18_63 (.ZN (n_18_63), .A (n_22_61), .B (n_28_58), .C1 (n_32_56), .C2 (n_38_53) );
AOI211_X1 g_16_64 (.ZN (n_16_64), .A (n_20_62), .B (n_26_59), .C1 (n_30_57), .C2 (n_36_54) );
AOI211_X1 g_14_65 (.ZN (n_14_65), .A (n_18_63), .B (n_24_60), .C1 (n_28_58), .C2 (n_34_55) );
AOI211_X1 g_15_63 (.ZN (n_15_63), .A (n_16_64), .B (n_22_61), .C1 (n_26_59), .C2 (n_32_56) );
AOI211_X1 g_16_65 (.ZN (n_16_65), .A (n_14_65), .B (n_20_62), .C1 (n_24_60), .C2 (n_30_57) );
AOI211_X1 g_14_66 (.ZN (n_14_66), .A (n_15_63), .B (n_18_63), .C1 (n_22_61), .C2 (n_28_58) );
AOI211_X1 g_13_64 (.ZN (n_13_64), .A (n_16_65), .B (n_16_64), .C1 (n_20_62), .C2 (n_26_59) );
AOI211_X1 g_11_63 (.ZN (n_11_63), .A (n_14_66), .B (n_14_65), .C1 (n_18_63), .C2 (n_24_60) );
AOI211_X1 g_12_65 (.ZN (n_12_65), .A (n_13_64), .B (n_15_63), .C1 (n_16_64), .C2 (n_22_61) );
AOI211_X1 g_10_66 (.ZN (n_10_66), .A (n_11_63), .B (n_16_65), .C1 (n_14_65), .C2 (n_20_62) );
AOI211_X1 g_9_64 (.ZN (n_9_64), .A (n_12_65), .B (n_14_66), .C1 (n_15_63), .C2 (n_18_63) );
AOI211_X1 g_7_65 (.ZN (n_7_65), .A (n_10_66), .B (n_13_64), .C1 (n_16_65), .C2 (n_16_64) );
AOI211_X1 g_6_67 (.ZN (n_6_67), .A (n_9_64), .B (n_11_63), .C1 (n_14_66), .C2 (n_14_65) );
AOI211_X1 g_8_66 (.ZN (n_8_66), .A (n_7_65), .B (n_12_65), .C1 (n_13_64), .C2 (n_15_63) );
AOI211_X1 g_10_65 (.ZN (n_10_65), .A (n_6_67), .B (n_10_66), .C1 (n_11_63), .C2 (n_16_65) );
AOI211_X1 g_9_67 (.ZN (n_9_67), .A (n_8_66), .B (n_9_64), .C1 (n_12_65), .C2 (n_14_66) );
AOI211_X1 g_7_68 (.ZN (n_7_68), .A (n_10_65), .B (n_7_65), .C1 (n_10_66), .C2 (n_13_64) );
AOI211_X1 g_5_69 (.ZN (n_5_69), .A (n_9_67), .B (n_6_67), .C1 (n_9_64), .C2 (n_11_63) );
AOI211_X1 g_4_71 (.ZN (n_4_71), .A (n_7_68), .B (n_8_66), .C1 (n_7_65), .C2 (n_12_65) );
AOI211_X1 g_6_70 (.ZN (n_6_70), .A (n_5_69), .B (n_10_65), .C1 (n_6_67), .C2 (n_10_66) );
AOI211_X1 g_5_68 (.ZN (n_5_68), .A (n_4_71), .B (n_9_67), .C1 (n_8_66), .C2 (n_9_64) );
AOI211_X1 g_7_67 (.ZN (n_7_67), .A (n_6_70), .B (n_7_68), .C1 (n_10_65), .C2 (n_7_65) );
AOI211_X1 g_9_66 (.ZN (n_9_66), .A (n_5_68), .B (n_5_69), .C1 (n_9_67), .C2 (n_6_67) );
AOI211_X1 g_11_65 (.ZN (n_11_65), .A (n_7_67), .B (n_4_71), .C1 (n_7_68), .C2 (n_8_66) );
AOI211_X1 g_12_67 (.ZN (n_12_67), .A (n_9_66), .B (n_6_70), .C1 (n_5_69), .C2 (n_10_65) );
AOI211_X1 g_10_68 (.ZN (n_10_68), .A (n_11_65), .B (n_5_68), .C1 (n_4_71), .C2 (n_9_67) );
AOI211_X1 g_8_67 (.ZN (n_8_67), .A (n_12_67), .B (n_7_67), .C1 (n_6_70), .C2 (n_7_68) );
AOI211_X1 g_6_68 (.ZN (n_6_68), .A (n_10_68), .B (n_9_66), .C1 (n_5_68), .C2 (n_5_69) );
AOI211_X1 g_8_69 (.ZN (n_8_69), .A (n_8_67), .B (n_11_65), .C1 (n_7_67), .C2 (n_4_71) );
AOI211_X1 g_7_71 (.ZN (n_7_71), .A (n_6_68), .B (n_12_67), .C1 (n_9_66), .C2 (n_6_70) );
AOI211_X1 g_6_69 (.ZN (n_6_69), .A (n_8_69), .B (n_10_68), .C1 (n_11_65), .C2 (n_5_68) );
AOI211_X1 g_4_70 (.ZN (n_4_70), .A (n_7_71), .B (n_8_67), .C1 (n_12_67), .C2 (n_7_67) );
AOI211_X1 g_5_72 (.ZN (n_5_72), .A (n_6_69), .B (n_6_68), .C1 (n_10_68), .C2 (n_9_66) );
AOI211_X1 g_4_74 (.ZN (n_4_74), .A (n_4_70), .B (n_8_69), .C1 (n_8_67), .C2 (n_11_65) );
AOI211_X1 g_3_72 (.ZN (n_3_72), .A (n_5_72), .B (n_7_71), .C1 (n_6_68), .C2 (n_12_67) );
AOI211_X1 g_2_74 (.ZN (n_2_74), .A (n_4_74), .B (n_6_69), .C1 (n_8_69), .C2 (n_10_68) );
AOI211_X1 g_4_73 (.ZN (n_4_73), .A (n_3_72), .B (n_4_70), .C1 (n_7_71), .C2 (n_8_67) );
AOI211_X1 g_5_71 (.ZN (n_5_71), .A (n_2_74), .B (n_5_72), .C1 (n_6_69), .C2 (n_6_68) );
AOI211_X1 g_6_73 (.ZN (n_6_73), .A (n_4_73), .B (n_4_74), .C1 (n_4_70), .C2 (n_8_69) );
AOI211_X1 g_5_75 (.ZN (n_5_75), .A (n_5_71), .B (n_3_72), .C1 (n_5_72), .C2 (n_7_71) );
AOI211_X1 g_3_76 (.ZN (n_3_76), .A (n_6_73), .B (n_2_74), .C1 (n_4_74), .C2 (n_6_69) );
AOI211_X1 g_2_78 (.ZN (n_2_78), .A (n_5_75), .B (n_4_73), .C1 (n_3_72), .C2 (n_4_70) );
AOI211_X1 g_4_77 (.ZN (n_4_77), .A (n_3_76), .B (n_5_71), .C1 (n_2_74), .C2 (n_5_72) );
AOI211_X1 g_6_76 (.ZN (n_6_76), .A (n_2_78), .B (n_6_73), .C1 (n_4_73), .C2 (n_4_74) );
AOI211_X1 g_4_75 (.ZN (n_4_75), .A (n_4_77), .B (n_5_75), .C1 (n_5_71), .C2 (n_3_72) );
AOI211_X1 g_5_73 (.ZN (n_5_73), .A (n_6_76), .B (n_3_76), .C1 (n_6_73), .C2 (n_2_74) );
AOI211_X1 g_6_71 (.ZN (n_6_71), .A (n_4_75), .B (n_2_78), .C1 (n_5_75), .C2 (n_4_73) );
AOI211_X1 g_7_69 (.ZN (n_7_69), .A (n_5_73), .B (n_4_77), .C1 (n_3_76), .C2 (n_5_71) );
AOI211_X1 g_9_68 (.ZN (n_9_68), .A (n_6_71), .B (n_6_76), .C1 (n_2_78), .C2 (n_6_73) );
AOI211_X1 g_11_67 (.ZN (n_11_67), .A (n_7_69), .B (n_4_75), .C1 (n_4_77), .C2 (n_5_75) );
AOI211_X1 g_13_66 (.ZN (n_13_66), .A (n_9_68), .B (n_5_73), .C1 (n_6_76), .C2 (n_3_76) );
AOI211_X1 g_15_65 (.ZN (n_15_65), .A (n_11_67), .B (n_6_71), .C1 (n_4_75), .C2 (n_2_78) );
AOI211_X1 g_17_64 (.ZN (n_17_64), .A (n_13_66), .B (n_7_69), .C1 (n_5_73), .C2 (n_4_77) );
AOI211_X1 g_19_63 (.ZN (n_19_63), .A (n_15_65), .B (n_9_68), .C1 (n_6_71), .C2 (n_6_76) );
AOI211_X1 g_21_62 (.ZN (n_21_62), .A (n_17_64), .B (n_11_67), .C1 (n_7_69), .C2 (n_4_75) );
AOI211_X1 g_22_60 (.ZN (n_22_60), .A (n_19_63), .B (n_13_66), .C1 (n_9_68), .C2 (n_5_73) );
AOI211_X1 g_24_59 (.ZN (n_24_59), .A (n_21_62), .B (n_15_65), .C1 (n_11_67), .C2 (n_6_71) );
AOI211_X1 g_26_58 (.ZN (n_26_58), .A (n_22_60), .B (n_17_64), .C1 (n_13_66), .C2 (n_7_69) );
AOI211_X1 g_28_57 (.ZN (n_28_57), .A (n_24_59), .B (n_19_63), .C1 (n_15_65), .C2 (n_9_68) );
AOI211_X1 g_30_56 (.ZN (n_30_56), .A (n_26_58), .B (n_21_62), .C1 (n_17_64), .C2 (n_11_67) );
AOI211_X1 g_32_55 (.ZN (n_32_55), .A (n_28_57), .B (n_22_60), .C1 (n_19_63), .C2 (n_13_66) );
AOI211_X1 g_34_56 (.ZN (n_34_56), .A (n_30_56), .B (n_24_59), .C1 (n_21_62), .C2 (n_15_65) );
AOI211_X1 g_32_57 (.ZN (n_32_57), .A (n_32_55), .B (n_26_58), .C1 (n_22_60), .C2 (n_17_64) );
AOI211_X1 g_30_58 (.ZN (n_30_58), .A (n_34_56), .B (n_28_57), .C1 (n_24_59), .C2 (n_19_63) );
AOI211_X1 g_28_59 (.ZN (n_28_59), .A (n_32_57), .B (n_30_56), .C1 (n_26_58), .C2 (n_21_62) );
AOI211_X1 g_26_60 (.ZN (n_26_60), .A (n_30_58), .B (n_32_55), .C1 (n_28_57), .C2 (n_22_60) );
AOI211_X1 g_24_61 (.ZN (n_24_61), .A (n_28_59), .B (n_34_56), .C1 (n_30_56), .C2 (n_24_59) );
AOI211_X1 g_22_62 (.ZN (n_22_62), .A (n_26_60), .B (n_32_57), .C1 (n_32_55), .C2 (n_26_58) );
AOI211_X1 g_20_63 (.ZN (n_20_63), .A (n_24_61), .B (n_30_58), .C1 (n_34_56), .C2 (n_28_57) );
AOI211_X1 g_19_65 (.ZN (n_19_65), .A (n_22_62), .B (n_28_59), .C1 (n_32_57), .C2 (n_30_56) );
AOI211_X1 g_21_64 (.ZN (n_21_64), .A (n_20_63), .B (n_26_60), .C1 (n_30_58), .C2 (n_32_55) );
AOI211_X1 g_23_63 (.ZN (n_23_63), .A (n_19_65), .B (n_24_61), .C1 (n_28_59), .C2 (n_34_56) );
AOI211_X1 g_25_62 (.ZN (n_25_62), .A (n_21_64), .B (n_22_62), .C1 (n_26_60), .C2 (n_32_57) );
AOI211_X1 g_23_61 (.ZN (n_23_61), .A (n_23_63), .B (n_20_63), .C1 (n_24_61), .C2 (n_30_58) );
AOI211_X1 g_25_60 (.ZN (n_25_60), .A (n_25_62), .B (n_19_65), .C1 (n_22_62), .C2 (n_28_59) );
AOI211_X1 g_27_59 (.ZN (n_27_59), .A (n_23_61), .B (n_21_64), .C1 (n_20_63), .C2 (n_26_60) );
AOI211_X1 g_29_58 (.ZN (n_29_58), .A (n_25_60), .B (n_23_63), .C1 (n_19_65), .C2 (n_24_61) );
AOI211_X1 g_31_57 (.ZN (n_31_57), .A (n_27_59), .B (n_25_62), .C1 (n_21_64), .C2 (n_22_62) );
AOI211_X1 g_33_56 (.ZN (n_33_56), .A (n_29_58), .B (n_23_61), .C1 (n_23_63), .C2 (n_20_63) );
AOI211_X1 g_35_55 (.ZN (n_35_55), .A (n_31_57), .B (n_25_60), .C1 (n_25_62), .C2 (n_19_65) );
AOI211_X1 g_37_54 (.ZN (n_37_54), .A (n_33_56), .B (n_27_59), .C1 (n_23_61), .C2 (n_21_64) );
AOI211_X1 g_39_53 (.ZN (n_39_53), .A (n_35_55), .B (n_29_58), .C1 (n_25_60), .C2 (n_23_63) );
AOI211_X1 g_41_52 (.ZN (n_41_52), .A (n_37_54), .B (n_31_57), .C1 (n_27_59), .C2 (n_25_62) );
AOI211_X1 g_40_54 (.ZN (n_40_54), .A (n_39_53), .B (n_33_56), .C1 (n_29_58), .C2 (n_23_61) );
AOI211_X1 g_42_53 (.ZN (n_42_53), .A (n_41_52), .B (n_35_55), .C1 (n_31_57), .C2 (n_25_60) );
AOI211_X1 g_44_52 (.ZN (n_44_52), .A (n_40_54), .B (n_37_54), .C1 (n_33_56), .C2 (n_27_59) );
AOI211_X1 g_46_51 (.ZN (n_46_51), .A (n_42_53), .B (n_39_53), .C1 (n_35_55), .C2 (n_29_58) );
AOI211_X1 g_48_50 (.ZN (n_48_50), .A (n_44_52), .B (n_41_52), .C1 (n_37_54), .C2 (n_31_57) );
AOI211_X1 g_50_49 (.ZN (n_50_49), .A (n_46_51), .B (n_40_54), .C1 (n_39_53), .C2 (n_33_56) );
AOI211_X1 g_52_48 (.ZN (n_52_48), .A (n_48_50), .B (n_42_53), .C1 (n_41_52), .C2 (n_35_55) );
AOI211_X1 g_51_50 (.ZN (n_51_50), .A (n_50_49), .B (n_44_52), .C1 (n_40_54), .C2 (n_37_54) );
AOI211_X1 g_49_49 (.ZN (n_49_49), .A (n_52_48), .B (n_46_51), .C1 (n_42_53), .C2 (n_39_53) );
AOI211_X1 g_51_48 (.ZN (n_51_48), .A (n_51_50), .B (n_48_50), .C1 (n_44_52), .C2 (n_41_52) );
AOI211_X1 g_53_47 (.ZN (n_53_47), .A (n_49_49), .B (n_50_49), .C1 (n_46_51), .C2 (n_40_54) );
AOI211_X1 g_55_46 (.ZN (n_55_46), .A (n_51_48), .B (n_52_48), .C1 (n_48_50), .C2 (n_42_53) );
AOI211_X1 g_57_45 (.ZN (n_57_45), .A (n_53_47), .B (n_51_50), .C1 (n_50_49), .C2 (n_44_52) );
AOI211_X1 g_58_47 (.ZN (n_58_47), .A (n_55_46), .B (n_49_49), .C1 (n_52_48), .C2 (n_46_51) );
AOI211_X1 g_56_48 (.ZN (n_56_48), .A (n_57_45), .B (n_51_48), .C1 (n_51_50), .C2 (n_48_50) );
AOI211_X1 g_57_46 (.ZN (n_57_46), .A (n_58_47), .B (n_53_47), .C1 (n_49_49), .C2 (n_50_49) );
AOI211_X1 g_55_47 (.ZN (n_55_47), .A (n_56_48), .B (n_55_46), .C1 (n_51_48), .C2 (n_52_48) );
AOI211_X1 g_53_48 (.ZN (n_53_48), .A (n_57_46), .B (n_57_45), .C1 (n_53_47), .C2 (n_51_50) );
AOI211_X1 g_51_49 (.ZN (n_51_49), .A (n_55_47), .B (n_58_47), .C1 (n_55_46), .C2 (n_49_49) );
AOI211_X1 g_49_50 (.ZN (n_49_50), .A (n_53_48), .B (n_56_48), .C1 (n_57_45), .C2 (n_51_48) );
AOI211_X1 g_47_51 (.ZN (n_47_51), .A (n_51_49), .B (n_57_46), .C1 (n_58_47), .C2 (n_53_47) );
AOI211_X1 g_45_52 (.ZN (n_45_52), .A (n_49_50), .B (n_55_47), .C1 (n_56_48), .C2 (n_55_46) );
AOI211_X1 g_43_53 (.ZN (n_43_53), .A (n_47_51), .B (n_53_48), .C1 (n_57_46), .C2 (n_57_45) );
AOI211_X1 g_41_54 (.ZN (n_41_54), .A (n_45_52), .B (n_51_49), .C1 (n_55_47), .C2 (n_58_47) );
AOI211_X1 g_39_55 (.ZN (n_39_55), .A (n_43_53), .B (n_49_50), .C1 (n_53_48), .C2 (n_56_48) );
AOI211_X1 g_37_56 (.ZN (n_37_56), .A (n_41_54), .B (n_47_51), .C1 (n_51_49), .C2 (n_57_46) );
AOI211_X1 g_35_57 (.ZN (n_35_57), .A (n_39_55), .B (n_45_52), .C1 (n_49_50), .C2 (n_55_47) );
AOI211_X1 g_33_58 (.ZN (n_33_58), .A (n_37_56), .B (n_43_53), .C1 (n_47_51), .C2 (n_53_48) );
AOI211_X1 g_31_59 (.ZN (n_31_59), .A (n_35_57), .B (n_41_54), .C1 (n_45_52), .C2 (n_51_49) );
AOI211_X1 g_29_60 (.ZN (n_29_60), .A (n_33_58), .B (n_39_55), .C1 (n_43_53), .C2 (n_49_50) );
AOI211_X1 g_27_61 (.ZN (n_27_61), .A (n_31_59), .B (n_37_56), .C1 (n_41_54), .C2 (n_47_51) );
AOI211_X1 g_26_63 (.ZN (n_26_63), .A (n_29_60), .B (n_35_57), .C1 (n_39_55), .C2 (n_45_52) );
AOI211_X1 g_25_61 (.ZN (n_25_61), .A (n_27_61), .B (n_33_58), .C1 (n_37_56), .C2 (n_43_53) );
AOI211_X1 g_27_60 (.ZN (n_27_60), .A (n_26_63), .B (n_31_59), .C1 (n_35_57), .C2 (n_41_54) );
AOI211_X1 g_29_59 (.ZN (n_29_59), .A (n_25_61), .B (n_29_60), .C1 (n_33_58), .C2 (n_39_55) );
AOI211_X1 g_31_58 (.ZN (n_31_58), .A (n_27_60), .B (n_27_61), .C1 (n_31_59), .C2 (n_37_56) );
AOI211_X1 g_33_57 (.ZN (n_33_57), .A (n_29_59), .B (n_26_63), .C1 (n_29_60), .C2 (n_35_57) );
AOI211_X1 g_35_56 (.ZN (n_35_56), .A (n_31_58), .B (n_25_61), .C1 (n_27_61), .C2 (n_33_58) );
AOI211_X1 g_37_55 (.ZN (n_37_55), .A (n_33_57), .B (n_27_60), .C1 (n_26_63), .C2 (n_31_59) );
AOI211_X1 g_39_54 (.ZN (n_39_54), .A (n_35_56), .B (n_29_59), .C1 (n_25_61), .C2 (n_29_60) );
AOI211_X1 g_41_53 (.ZN (n_41_53), .A (n_37_55), .B (n_31_58), .C1 (n_27_60), .C2 (n_27_61) );
AOI211_X1 g_43_52 (.ZN (n_43_52), .A (n_39_54), .B (n_33_57), .C1 (n_29_59), .C2 (n_26_63) );
AOI211_X1 g_45_51 (.ZN (n_45_51), .A (n_41_53), .B (n_35_56), .C1 (n_31_58), .C2 (n_25_61) );
AOI211_X1 g_47_50 (.ZN (n_47_50), .A (n_43_52), .B (n_37_55), .C1 (n_33_57), .C2 (n_27_60) );
AOI211_X1 g_49_51 (.ZN (n_49_51), .A (n_45_51), .B (n_39_54), .C1 (n_35_56), .C2 (n_29_59) );
AOI211_X1 g_47_52 (.ZN (n_47_52), .A (n_47_50), .B (n_41_53), .C1 (n_37_55), .C2 (n_31_58) );
AOI211_X1 g_45_53 (.ZN (n_45_53), .A (n_49_51), .B (n_43_52), .C1 (n_39_54), .C2 (n_33_57) );
AOI211_X1 g_43_54 (.ZN (n_43_54), .A (n_47_52), .B (n_45_51), .C1 (n_41_53), .C2 (n_35_56) );
AOI211_X1 g_41_55 (.ZN (n_41_55), .A (n_45_53), .B (n_47_50), .C1 (n_43_52), .C2 (n_37_55) );
AOI211_X1 g_39_56 (.ZN (n_39_56), .A (n_43_54), .B (n_49_51), .C1 (n_45_51), .C2 (n_39_54) );
AOI211_X1 g_37_57 (.ZN (n_37_57), .A (n_41_55), .B (n_47_52), .C1 (n_47_50), .C2 (n_41_53) );
AOI211_X1 g_38_55 (.ZN (n_38_55), .A (n_39_56), .B (n_45_53), .C1 (n_49_51), .C2 (n_43_52) );
AOI211_X1 g_36_56 (.ZN (n_36_56), .A (n_37_57), .B (n_43_54), .C1 (n_47_52), .C2 (n_45_51) );
AOI211_X1 g_34_57 (.ZN (n_34_57), .A (n_38_55), .B (n_41_55), .C1 (n_45_53), .C2 (n_47_50) );
AOI211_X1 g_32_58 (.ZN (n_32_58), .A (n_36_56), .B (n_39_56), .C1 (n_43_54), .C2 (n_49_51) );
AOI211_X1 g_30_59 (.ZN (n_30_59), .A (n_34_57), .B (n_37_57), .C1 (n_41_55), .C2 (n_47_52) );
AOI211_X1 g_28_60 (.ZN (n_28_60), .A (n_32_58), .B (n_38_55), .C1 (n_39_56), .C2 (n_45_53) );
AOI211_X1 g_26_61 (.ZN (n_26_61), .A (n_30_59), .B (n_36_56), .C1 (n_37_57), .C2 (n_43_54) );
AOI211_X1 g_24_62 (.ZN (n_24_62), .A (n_28_60), .B (n_34_57), .C1 (n_38_55), .C2 (n_41_55) );
AOI211_X1 g_22_63 (.ZN (n_22_63), .A (n_26_61), .B (n_32_58), .C1 (n_36_56), .C2 (n_39_56) );
AOI211_X1 g_20_64 (.ZN (n_20_64), .A (n_24_62), .B (n_30_59), .C1 (n_34_57), .C2 (n_37_57) );
AOI211_X1 g_18_65 (.ZN (n_18_65), .A (n_22_63), .B (n_28_60), .C1 (n_32_58), .C2 (n_38_55) );
AOI211_X1 g_16_66 (.ZN (n_16_66), .A (n_20_64), .B (n_26_61), .C1 (n_30_59), .C2 (n_36_56) );
AOI211_X1 g_14_67 (.ZN (n_14_67), .A (n_18_65), .B (n_24_62), .C1 (n_28_60), .C2 (n_34_57) );
AOI211_X1 g_12_66 (.ZN (n_12_66), .A (n_16_66), .B (n_22_63), .C1 (n_26_61), .C2 (n_32_58) );
AOI211_X1 g_10_67 (.ZN (n_10_67), .A (n_14_67), .B (n_20_64), .C1 (n_24_62), .C2 (n_30_59) );
AOI211_X1 g_8_68 (.ZN (n_8_68), .A (n_12_66), .B (n_18_65), .C1 (n_22_63), .C2 (n_28_60) );
AOI211_X1 g_7_70 (.ZN (n_7_70), .A (n_10_67), .B (n_16_66), .C1 (n_20_64), .C2 (n_26_61) );
AOI211_X1 g_6_72 (.ZN (n_6_72), .A (n_8_68), .B (n_14_67), .C1 (n_18_65), .C2 (n_24_62) );
AOI211_X1 g_7_74 (.ZN (n_7_74), .A (n_7_70), .B (n_12_66), .C1 (n_16_66), .C2 (n_22_63) );
AOI211_X1 g_8_72 (.ZN (n_8_72), .A (n_6_72), .B (n_10_67), .C1 (n_14_67), .C2 (n_20_64) );
AOI211_X1 g_9_70 (.ZN (n_9_70), .A (n_7_74), .B (n_8_68), .C1 (n_12_66), .C2 (n_18_65) );
AOI211_X1 g_11_69 (.ZN (n_11_69), .A (n_8_72), .B (n_7_70), .C1 (n_10_67), .C2 (n_16_66) );
AOI211_X1 g_13_68 (.ZN (n_13_68), .A (n_9_70), .B (n_6_72), .C1 (n_8_68), .C2 (n_14_67) );
AOI211_X1 g_15_67 (.ZN (n_15_67), .A (n_11_69), .B (n_7_74), .C1 (n_7_70), .C2 (n_12_66) );
AOI211_X1 g_17_66 (.ZN (n_17_66), .A (n_13_68), .B (n_8_72), .C1 (n_6_72), .C2 (n_10_67) );
AOI211_X1 g_16_68 (.ZN (n_16_68), .A (n_15_67), .B (n_9_70), .C1 (n_7_74), .C2 (n_8_68) );
AOI211_X1 g_15_66 (.ZN (n_15_66), .A (n_17_66), .B (n_11_69), .C1 (n_8_72), .C2 (n_7_70) );
AOI211_X1 g_17_65 (.ZN (n_17_65), .A (n_16_68), .B (n_13_68), .C1 (n_9_70), .C2 (n_6_72) );
AOI211_X1 g_19_64 (.ZN (n_19_64), .A (n_15_66), .B (n_15_67), .C1 (n_11_69), .C2 (n_7_74) );
AOI211_X1 g_21_63 (.ZN (n_21_63), .A (n_17_65), .B (n_17_66), .C1 (n_13_68), .C2 (n_8_72) );
AOI211_X1 g_23_62 (.ZN (n_23_62), .A (n_19_64), .B (n_16_68), .C1 (n_15_67), .C2 (n_9_70) );
AOI211_X1 g_24_64 (.ZN (n_24_64), .A (n_21_63), .B (n_15_66), .C1 (n_17_66), .C2 (n_11_69) );
AOI211_X1 g_22_65 (.ZN (n_22_65), .A (n_23_62), .B (n_17_65), .C1 (n_16_68), .C2 (n_13_68) );
AOI211_X1 g_20_66 (.ZN (n_20_66), .A (n_24_64), .B (n_19_64), .C1 (n_15_66), .C2 (n_15_67) );
AOI211_X1 g_18_67 (.ZN (n_18_67), .A (n_22_65), .B (n_21_63), .C1 (n_17_65), .C2 (n_17_66) );
AOI211_X1 g_17_69 (.ZN (n_17_69), .A (n_20_66), .B (n_23_62), .C1 (n_19_64), .C2 (n_16_68) );
AOI211_X1 g_16_67 (.ZN (n_16_67), .A (n_18_67), .B (n_24_64), .C1 (n_21_63), .C2 (n_15_66) );
AOI211_X1 g_18_66 (.ZN (n_18_66), .A (n_17_69), .B (n_22_65), .C1 (n_23_62), .C2 (n_17_65) );
AOI211_X1 g_20_65 (.ZN (n_20_65), .A (n_16_67), .B (n_20_66), .C1 (n_24_64), .C2 (n_19_64) );
AOI211_X1 g_22_64 (.ZN (n_22_64), .A (n_18_66), .B (n_18_67), .C1 (n_22_65), .C2 (n_21_63) );
AOI211_X1 g_24_63 (.ZN (n_24_63), .A (n_20_65), .B (n_17_69), .C1 (n_20_66), .C2 (n_23_62) );
AOI211_X1 g_26_62 (.ZN (n_26_62), .A (n_22_64), .B (n_16_67), .C1 (n_18_67), .C2 (n_24_64) );
AOI211_X1 g_28_61 (.ZN (n_28_61), .A (n_24_63), .B (n_18_66), .C1 (n_17_69), .C2 (n_22_65) );
AOI211_X1 g_30_60 (.ZN (n_30_60), .A (n_26_62), .B (n_20_65), .C1 (n_16_67), .C2 (n_20_66) );
AOI211_X1 g_32_59 (.ZN (n_32_59), .A (n_28_61), .B (n_22_64), .C1 (n_18_66), .C2 (n_18_67) );
AOI211_X1 g_34_58 (.ZN (n_34_58), .A (n_30_60), .B (n_24_63), .C1 (n_20_65), .C2 (n_17_69) );
AOI211_X1 g_36_57 (.ZN (n_36_57), .A (n_32_59), .B (n_26_62), .C1 (n_22_64), .C2 (n_16_67) );
AOI211_X1 g_38_56 (.ZN (n_38_56), .A (n_34_58), .B (n_28_61), .C1 (n_24_63), .C2 (n_18_66) );
AOI211_X1 g_40_55 (.ZN (n_40_55), .A (n_36_57), .B (n_30_60), .C1 (n_26_62), .C2 (n_20_65) );
AOI211_X1 g_42_54 (.ZN (n_42_54), .A (n_38_56), .B (n_32_59), .C1 (n_28_61), .C2 (n_22_64) );
AOI211_X1 g_44_53 (.ZN (n_44_53), .A (n_40_55), .B (n_34_58), .C1 (n_30_60), .C2 (n_24_63) );
AOI211_X1 g_46_52 (.ZN (n_46_52), .A (n_42_54), .B (n_36_57), .C1 (n_32_59), .C2 (n_26_62) );
AOI211_X1 g_48_51 (.ZN (n_48_51), .A (n_44_53), .B (n_38_56), .C1 (n_34_58), .C2 (n_28_61) );
AOI211_X1 g_50_50 (.ZN (n_50_50), .A (n_46_52), .B (n_40_55), .C1 (n_36_57), .C2 (n_30_60) );
AOI211_X1 g_52_49 (.ZN (n_52_49), .A (n_48_51), .B (n_42_54), .C1 (n_38_56), .C2 (n_32_59) );
AOI211_X1 g_54_48 (.ZN (n_54_48), .A (n_50_50), .B (n_44_53), .C1 (n_40_55), .C2 (n_34_58) );
AOI211_X1 g_56_47 (.ZN (n_56_47), .A (n_52_49), .B (n_46_52), .C1 (n_42_54), .C2 (n_36_57) );
AOI211_X1 g_58_46 (.ZN (n_58_46), .A (n_54_48), .B (n_48_51), .C1 (n_44_53), .C2 (n_38_56) );
AOI211_X1 g_60_45 (.ZN (n_60_45), .A (n_56_47), .B (n_50_50), .C1 (n_46_52), .C2 (n_40_55) );
AOI211_X1 g_62_44 (.ZN (n_62_44), .A (n_58_46), .B (n_52_49), .C1 (n_48_51), .C2 (n_42_54) );
AOI211_X1 g_64_43 (.ZN (n_64_43), .A (n_60_45), .B (n_54_48), .C1 (n_50_50), .C2 (n_44_53) );
AOI211_X1 g_66_42 (.ZN (n_66_42), .A (n_62_44), .B (n_56_47), .C1 (n_52_49), .C2 (n_46_52) );
AOI211_X1 g_68_41 (.ZN (n_68_41), .A (n_64_43), .B (n_58_46), .C1 (n_54_48), .C2 (n_48_51) );
AOI211_X1 g_70_40 (.ZN (n_70_40), .A (n_66_42), .B (n_60_45), .C1 (n_56_47), .C2 (n_50_50) );
AOI211_X1 g_72_39 (.ZN (n_72_39), .A (n_68_41), .B (n_62_44), .C1 (n_58_46), .C2 (n_52_49) );
AOI211_X1 g_73_37 (.ZN (n_73_37), .A (n_70_40), .B (n_64_43), .C1 (n_60_45), .C2 (n_54_48) );
AOI211_X1 g_75_36 (.ZN (n_75_36), .A (n_72_39), .B (n_66_42), .C1 (n_62_44), .C2 (n_56_47) );
AOI211_X1 g_77_35 (.ZN (n_77_35), .A (n_73_37), .B (n_68_41), .C1 (n_64_43), .C2 (n_58_46) );
AOI211_X1 g_79_34 (.ZN (n_79_34), .A (n_75_36), .B (n_70_40), .C1 (n_66_42), .C2 (n_60_45) );
AOI211_X1 g_81_33 (.ZN (n_81_33), .A (n_77_35), .B (n_72_39), .C1 (n_68_41), .C2 (n_62_44) );
AOI211_X1 g_83_32 (.ZN (n_83_32), .A (n_79_34), .B (n_73_37), .C1 (n_70_40), .C2 (n_64_43) );
AOI211_X1 g_85_31 (.ZN (n_85_31), .A (n_81_33), .B (n_75_36), .C1 (n_72_39), .C2 (n_66_42) );
AOI211_X1 g_87_30 (.ZN (n_87_30), .A (n_83_32), .B (n_77_35), .C1 (n_73_37), .C2 (n_68_41) );
AOI211_X1 g_89_29 (.ZN (n_89_29), .A (n_85_31), .B (n_79_34), .C1 (n_75_36), .C2 (n_70_40) );
AOI211_X1 g_91_28 (.ZN (n_91_28), .A (n_87_30), .B (n_81_33), .C1 (n_77_35), .C2 (n_72_39) );
AOI211_X1 g_93_27 (.ZN (n_93_27), .A (n_89_29), .B (n_83_32), .C1 (n_79_34), .C2 (n_73_37) );
AOI211_X1 g_95_26 (.ZN (n_95_26), .A (n_91_28), .B (n_85_31), .C1 (n_81_33), .C2 (n_75_36) );
AOI211_X1 g_97_25 (.ZN (n_97_25), .A (n_93_27), .B (n_87_30), .C1 (n_83_32), .C2 (n_77_35) );
AOI211_X1 g_99_26 (.ZN (n_99_26), .A (n_95_26), .B (n_89_29), .C1 (n_85_31), .C2 (n_79_34) );
AOI211_X1 g_97_27 (.ZN (n_97_27), .A (n_97_25), .B (n_91_28), .C1 (n_87_30), .C2 (n_81_33) );
AOI211_X1 g_95_28 (.ZN (n_95_28), .A (n_99_26), .B (n_93_27), .C1 (n_89_29), .C2 (n_83_32) );
AOI211_X1 g_93_29 (.ZN (n_93_29), .A (n_97_27), .B (n_95_26), .C1 (n_91_28), .C2 (n_85_31) );
AOI211_X1 g_91_30 (.ZN (n_91_30), .A (n_95_28), .B (n_97_25), .C1 (n_93_27), .C2 (n_87_30) );
AOI211_X1 g_89_31 (.ZN (n_89_31), .A (n_93_29), .B (n_99_26), .C1 (n_95_26), .C2 (n_89_29) );
AOI211_X1 g_87_32 (.ZN (n_87_32), .A (n_91_30), .B (n_97_27), .C1 (n_97_25), .C2 (n_91_28) );
AOI211_X1 g_85_33 (.ZN (n_85_33), .A (n_89_31), .B (n_95_28), .C1 (n_99_26), .C2 (n_93_27) );
AOI211_X1 g_86_31 (.ZN (n_86_31), .A (n_87_32), .B (n_93_29), .C1 (n_97_27), .C2 (n_95_26) );
AOI211_X1 g_84_32 (.ZN (n_84_32), .A (n_85_33), .B (n_91_30), .C1 (n_95_28), .C2 (n_97_25) );
AOI211_X1 g_82_33 (.ZN (n_82_33), .A (n_86_31), .B (n_89_31), .C1 (n_93_29), .C2 (n_99_26) );
AOI211_X1 g_80_34 (.ZN (n_80_34), .A (n_84_32), .B (n_87_32), .C1 (n_91_30), .C2 (n_97_27) );
AOI211_X1 g_78_35 (.ZN (n_78_35), .A (n_82_33), .B (n_85_33), .C1 (n_89_31), .C2 (n_95_28) );
AOI211_X1 g_76_36 (.ZN (n_76_36), .A (n_80_34), .B (n_86_31), .C1 (n_87_32), .C2 (n_93_29) );
AOI211_X1 g_74_37 (.ZN (n_74_37), .A (n_78_35), .B (n_84_32), .C1 (n_85_33), .C2 (n_91_30) );
AOI211_X1 g_72_38 (.ZN (n_72_38), .A (n_76_36), .B (n_82_33), .C1 (n_86_31), .C2 (n_89_31) );
AOI211_X1 g_74_39 (.ZN (n_74_39), .A (n_74_37), .B (n_80_34), .C1 (n_84_32), .C2 (n_87_32) );
AOI211_X1 g_76_38 (.ZN (n_76_38), .A (n_72_38), .B (n_78_35), .C1 (n_82_33), .C2 (n_85_33) );
AOI211_X1 g_78_37 (.ZN (n_78_37), .A (n_74_39), .B (n_76_36), .C1 (n_80_34), .C2 (n_86_31) );
AOI211_X1 g_80_36 (.ZN (n_80_36), .A (n_76_38), .B (n_74_37), .C1 (n_78_35), .C2 (n_84_32) );
AOI211_X1 g_81_34 (.ZN (n_81_34), .A (n_78_37), .B (n_72_38), .C1 (n_76_36), .C2 (n_82_33) );
AOI211_X1 g_83_33 (.ZN (n_83_33), .A (n_80_36), .B (n_74_39), .C1 (n_74_37), .C2 (n_80_34) );
AOI211_X1 g_85_32 (.ZN (n_85_32), .A (n_81_34), .B (n_76_38), .C1 (n_72_38), .C2 (n_78_35) );
AOI211_X1 g_87_31 (.ZN (n_87_31), .A (n_83_33), .B (n_78_37), .C1 (n_74_39), .C2 (n_76_36) );
AOI211_X1 g_89_30 (.ZN (n_89_30), .A (n_85_32), .B (n_80_36), .C1 (n_76_38), .C2 (n_74_37) );
AOI211_X1 g_91_29 (.ZN (n_91_29), .A (n_87_31), .B (n_81_34), .C1 (n_78_37), .C2 (n_72_38) );
AOI211_X1 g_93_28 (.ZN (n_93_28), .A (n_89_30), .B (n_83_33), .C1 (n_80_36), .C2 (n_74_39) );
AOI211_X1 g_95_27 (.ZN (n_95_27), .A (n_91_29), .B (n_85_32), .C1 (n_81_34), .C2 (n_76_38) );
AOI211_X1 g_97_26 (.ZN (n_97_26), .A (n_93_28), .B (n_87_31), .C1 (n_83_33), .C2 (n_78_37) );
AOI211_X1 g_99_25 (.ZN (n_99_25), .A (n_95_27), .B (n_89_30), .C1 (n_85_32), .C2 (n_80_36) );
AOI211_X1 g_100_27 (.ZN (n_100_27), .A (n_97_26), .B (n_91_29), .C1 (n_87_31), .C2 (n_81_34) );
AOI211_X1 g_98_28 (.ZN (n_98_28), .A (n_99_25), .B (n_93_28), .C1 (n_89_30), .C2 (n_83_33) );
AOI211_X1 g_96_27 (.ZN (n_96_27), .A (n_100_27), .B (n_95_27), .C1 (n_91_29), .C2 (n_85_32) );
AOI211_X1 g_94_28 (.ZN (n_94_28), .A (n_98_28), .B (n_97_26), .C1 (n_93_28), .C2 (n_87_31) );
AOI211_X1 g_92_29 (.ZN (n_92_29), .A (n_96_27), .B (n_99_25), .C1 (n_95_27), .C2 (n_89_30) );
AOI211_X1 g_90_30 (.ZN (n_90_30), .A (n_94_28), .B (n_100_27), .C1 (n_97_26), .C2 (n_91_29) );
AOI211_X1 g_88_31 (.ZN (n_88_31), .A (n_92_29), .B (n_98_28), .C1 (n_99_25), .C2 (n_93_28) );
AOI211_X1 g_86_32 (.ZN (n_86_32), .A (n_90_30), .B (n_96_27), .C1 (n_100_27), .C2 (n_95_27) );
AOI211_X1 g_84_33 (.ZN (n_84_33), .A (n_88_31), .B (n_94_28), .C1 (n_98_28), .C2 (n_97_26) );
AOI211_X1 g_82_34 (.ZN (n_82_34), .A (n_86_32), .B (n_92_29), .C1 (n_96_27), .C2 (n_99_25) );
AOI211_X1 g_80_35 (.ZN (n_80_35), .A (n_84_33), .B (n_90_30), .C1 (n_94_28), .C2 (n_100_27) );
AOI211_X1 g_78_36 (.ZN (n_78_36), .A (n_82_34), .B (n_88_31), .C1 (n_92_29), .C2 (n_98_28) );
AOI211_X1 g_76_37 (.ZN (n_76_37), .A (n_80_35), .B (n_86_32), .C1 (n_90_30), .C2 (n_96_27) );
AOI211_X1 g_74_38 (.ZN (n_74_38), .A (n_78_36), .B (n_84_33), .C1 (n_88_31), .C2 (n_94_28) );
AOI211_X1 g_73_40 (.ZN (n_73_40), .A (n_76_37), .B (n_82_34), .C1 (n_86_32), .C2 (n_92_29) );
AOI211_X1 g_75_39 (.ZN (n_75_39), .A (n_74_38), .B (n_80_35), .C1 (n_84_33), .C2 (n_90_30) );
AOI211_X1 g_77_38 (.ZN (n_77_38), .A (n_73_40), .B (n_78_36), .C1 (n_82_34), .C2 (n_88_31) );
AOI211_X1 g_79_37 (.ZN (n_79_37), .A (n_75_39), .B (n_76_37), .C1 (n_80_35), .C2 (n_86_32) );
AOI211_X1 g_81_36 (.ZN (n_81_36), .A (n_77_38), .B (n_74_38), .C1 (n_78_36), .C2 (n_84_33) );
AOI211_X1 g_83_35 (.ZN (n_83_35), .A (n_79_37), .B (n_73_40), .C1 (n_76_37), .C2 (n_82_34) );
AOI211_X1 g_85_34 (.ZN (n_85_34), .A (n_81_36), .B (n_75_39), .C1 (n_74_38), .C2 (n_80_35) );
AOI211_X1 g_87_33 (.ZN (n_87_33), .A (n_83_35), .B (n_77_38), .C1 (n_73_40), .C2 (n_78_36) );
AOI211_X1 g_89_32 (.ZN (n_89_32), .A (n_85_34), .B (n_79_37), .C1 (n_75_39), .C2 (n_76_37) );
AOI211_X1 g_91_31 (.ZN (n_91_31), .A (n_87_33), .B (n_81_36), .C1 (n_77_38), .C2 (n_74_38) );
AOI211_X1 g_93_30 (.ZN (n_93_30), .A (n_89_32), .B (n_83_35), .C1 (n_79_37), .C2 (n_73_40) );
AOI211_X1 g_95_29 (.ZN (n_95_29), .A (n_91_31), .B (n_85_34), .C1 (n_81_36), .C2 (n_75_39) );
AOI211_X1 g_97_28 (.ZN (n_97_28), .A (n_93_30), .B (n_87_33), .C1 (n_83_35), .C2 (n_77_38) );
AOI211_X1 g_99_27 (.ZN (n_99_27), .A (n_95_29), .B (n_89_32), .C1 (n_85_34), .C2 (n_79_37) );
AOI211_X1 g_100_29 (.ZN (n_100_29), .A (n_97_28), .B (n_91_31), .C1 (n_87_33), .C2 (n_81_36) );
AOI211_X1 g_98_30 (.ZN (n_98_30), .A (n_99_27), .B (n_93_30), .C1 (n_89_32), .C2 (n_83_35) );
AOI211_X1 g_96_29 (.ZN (n_96_29), .A (n_100_29), .B (n_95_29), .C1 (n_91_31), .C2 (n_85_34) );
AOI211_X1 g_94_30 (.ZN (n_94_30), .A (n_98_30), .B (n_97_28), .C1 (n_93_30), .C2 (n_87_33) );
AOI211_X1 g_92_31 (.ZN (n_92_31), .A (n_96_29), .B (n_99_27), .C1 (n_95_29), .C2 (n_89_32) );
AOI211_X1 g_90_32 (.ZN (n_90_32), .A (n_94_30), .B (n_100_29), .C1 (n_97_28), .C2 (n_91_31) );
AOI211_X1 g_88_33 (.ZN (n_88_33), .A (n_92_31), .B (n_98_30), .C1 (n_99_27), .C2 (n_93_30) );
AOI211_X1 g_86_34 (.ZN (n_86_34), .A (n_90_32), .B (n_96_29), .C1 (n_100_29), .C2 (n_95_29) );
AOI211_X1 g_84_35 (.ZN (n_84_35), .A (n_88_33), .B (n_94_30), .C1 (n_98_30), .C2 (n_97_28) );
AOI211_X1 g_82_36 (.ZN (n_82_36), .A (n_86_34), .B (n_92_31), .C1 (n_96_29), .C2 (n_99_27) );
AOI211_X1 g_83_34 (.ZN (n_83_34), .A (n_84_35), .B (n_90_32), .C1 (n_94_30), .C2 (n_100_29) );
AOI211_X1 g_81_35 (.ZN (n_81_35), .A (n_82_36), .B (n_88_33), .C1 (n_92_31), .C2 (n_98_30) );
AOI211_X1 g_79_36 (.ZN (n_79_36), .A (n_83_34), .B (n_86_34), .C1 (n_90_32), .C2 (n_96_29) );
AOI211_X1 g_77_37 (.ZN (n_77_37), .A (n_81_35), .B (n_84_35), .C1 (n_88_33), .C2 (n_94_30) );
AOI211_X1 g_75_38 (.ZN (n_75_38), .A (n_79_36), .B (n_82_36), .C1 (n_86_34), .C2 (n_92_31) );
AOI211_X1 g_73_39 (.ZN (n_73_39), .A (n_77_37), .B (n_83_34), .C1 (n_84_35), .C2 (n_90_32) );
AOI211_X1 g_71_40 (.ZN (n_71_40), .A (n_75_38), .B (n_81_35), .C1 (n_82_36), .C2 (n_88_33) );
AOI211_X1 g_69_41 (.ZN (n_69_41), .A (n_73_39), .B (n_79_36), .C1 (n_83_34), .C2 (n_86_34) );
AOI211_X1 g_67_42 (.ZN (n_67_42), .A (n_71_40), .B (n_77_37), .C1 (n_81_35), .C2 (n_84_35) );
AOI211_X1 g_65_43 (.ZN (n_65_43), .A (n_69_41), .B (n_75_38), .C1 (n_79_36), .C2 (n_82_36) );
AOI211_X1 g_63_44 (.ZN (n_63_44), .A (n_67_42), .B (n_73_39), .C1 (n_77_37), .C2 (n_83_34) );
AOI211_X1 g_61_45 (.ZN (n_61_45), .A (n_65_43), .B (n_71_40), .C1 (n_75_38), .C2 (n_81_35) );
AOI211_X1 g_59_46 (.ZN (n_59_46), .A (n_63_44), .B (n_69_41), .C1 (n_73_39), .C2 (n_79_36) );
AOI211_X1 g_57_47 (.ZN (n_57_47), .A (n_61_45), .B (n_67_42), .C1 (n_71_40), .C2 (n_77_37) );
AOI211_X1 g_55_48 (.ZN (n_55_48), .A (n_59_46), .B (n_65_43), .C1 (n_69_41), .C2 (n_75_38) );
AOI211_X1 g_53_49 (.ZN (n_53_49), .A (n_57_47), .B (n_63_44), .C1 (n_67_42), .C2 (n_73_39) );
AOI211_X1 g_52_51 (.ZN (n_52_51), .A (n_55_48), .B (n_61_45), .C1 (n_65_43), .C2 (n_71_40) );
AOI211_X1 g_54_50 (.ZN (n_54_50), .A (n_53_49), .B (n_59_46), .C1 (n_63_44), .C2 (n_69_41) );
AOI211_X1 g_56_49 (.ZN (n_56_49), .A (n_52_51), .B (n_57_47), .C1 (n_61_45), .C2 (n_67_42) );
AOI211_X1 g_58_48 (.ZN (n_58_48), .A (n_54_50), .B (n_55_48), .C1 (n_59_46), .C2 (n_65_43) );
AOI211_X1 g_60_47 (.ZN (n_60_47), .A (n_56_49), .B (n_53_49), .C1 (n_57_47), .C2 (n_63_44) );
AOI211_X1 g_62_46 (.ZN (n_62_46), .A (n_58_48), .B (n_52_51), .C1 (n_55_48), .C2 (n_61_45) );
AOI211_X1 g_64_45 (.ZN (n_64_45), .A (n_60_47), .B (n_54_50), .C1 (n_53_49), .C2 (n_59_46) );
AOI211_X1 g_66_44 (.ZN (n_66_44), .A (n_62_46), .B (n_56_49), .C1 (n_52_51), .C2 (n_57_47) );
AOI211_X1 g_68_43 (.ZN (n_68_43), .A (n_64_45), .B (n_58_48), .C1 (n_54_50), .C2 (n_55_48) );
AOI211_X1 g_70_42 (.ZN (n_70_42), .A (n_66_44), .B (n_60_47), .C1 (n_56_49), .C2 (n_53_49) );
AOI211_X1 g_72_41 (.ZN (n_72_41), .A (n_68_43), .B (n_62_46), .C1 (n_58_48), .C2 (n_52_51) );
AOI211_X1 g_74_40 (.ZN (n_74_40), .A (n_70_42), .B (n_64_45), .C1 (n_60_47), .C2 (n_54_50) );
AOI211_X1 g_76_39 (.ZN (n_76_39), .A (n_72_41), .B (n_66_44), .C1 (n_62_46), .C2 (n_56_49) );
AOI211_X1 g_78_38 (.ZN (n_78_38), .A (n_74_40), .B (n_68_43), .C1 (n_64_45), .C2 (n_58_48) );
AOI211_X1 g_80_37 (.ZN (n_80_37), .A (n_76_39), .B (n_70_42), .C1 (n_66_44), .C2 (n_60_47) );
AOI211_X1 g_79_39 (.ZN (n_79_39), .A (n_78_38), .B (n_72_41), .C1 (n_68_43), .C2 (n_62_46) );
AOI211_X1 g_81_38 (.ZN (n_81_38), .A (n_80_37), .B (n_74_40), .C1 (n_70_42), .C2 (n_64_45) );
AOI211_X1 g_83_37 (.ZN (n_83_37), .A (n_79_39), .B (n_76_39), .C1 (n_72_41), .C2 (n_66_44) );
AOI211_X1 g_82_35 (.ZN (n_82_35), .A (n_81_38), .B (n_78_38), .C1 (n_74_40), .C2 (n_68_43) );
AOI211_X1 g_84_34 (.ZN (n_84_34), .A (n_83_37), .B (n_80_37), .C1 (n_76_39), .C2 (n_70_42) );
AOI211_X1 g_86_33 (.ZN (n_86_33), .A (n_82_35), .B (n_79_39), .C1 (n_78_38), .C2 (n_72_41) );
AOI211_X1 g_88_32 (.ZN (n_88_32), .A (n_84_34), .B (n_81_38), .C1 (n_80_37), .C2 (n_74_40) );
AOI211_X1 g_90_31 (.ZN (n_90_31), .A (n_86_33), .B (n_83_37), .C1 (n_79_39), .C2 (n_76_39) );
AOI211_X1 g_92_30 (.ZN (n_92_30), .A (n_88_32), .B (n_82_35), .C1 (n_81_38), .C2 (n_78_38) );
AOI211_X1 g_94_29 (.ZN (n_94_29), .A (n_90_31), .B (n_84_34), .C1 (n_83_37), .C2 (n_80_37) );
AOI211_X1 g_96_28 (.ZN (n_96_28), .A (n_92_30), .B (n_86_33), .C1 (n_82_35), .C2 (n_79_39) );
AOI211_X1 g_98_27 (.ZN (n_98_27), .A (n_94_29), .B (n_88_32), .C1 (n_84_34), .C2 (n_81_38) );
AOI211_X1 g_100_28 (.ZN (n_100_28), .A (n_96_28), .B (n_90_31), .C1 (n_86_33), .C2 (n_83_37) );
AOI211_X1 g_98_29 (.ZN (n_98_29), .A (n_98_27), .B (n_92_30), .C1 (n_88_32), .C2 (n_82_35) );
AOI211_X1 g_96_30 (.ZN (n_96_30), .A (n_100_28), .B (n_94_29), .C1 (n_90_31), .C2 (n_84_34) );
AOI211_X1 g_94_31 (.ZN (n_94_31), .A (n_98_29), .B (n_96_28), .C1 (n_92_30), .C2 (n_86_33) );
AOI211_X1 g_92_32 (.ZN (n_92_32), .A (n_96_30), .B (n_98_27), .C1 (n_94_29), .C2 (n_88_32) );
AOI211_X1 g_90_33 (.ZN (n_90_33), .A (n_94_31), .B (n_100_28), .C1 (n_96_28), .C2 (n_90_31) );
AOI211_X1 g_88_34 (.ZN (n_88_34), .A (n_92_32), .B (n_98_29), .C1 (n_98_27), .C2 (n_92_30) );
AOI211_X1 g_86_35 (.ZN (n_86_35), .A (n_90_33), .B (n_96_30), .C1 (n_100_28), .C2 (n_94_29) );
AOI211_X1 g_84_36 (.ZN (n_84_36), .A (n_88_34), .B (n_94_31), .C1 (n_98_29), .C2 (n_96_28) );
AOI211_X1 g_82_37 (.ZN (n_82_37), .A (n_86_35), .B (n_92_32), .C1 (n_96_30), .C2 (n_98_27) );
AOI211_X1 g_80_38 (.ZN (n_80_38), .A (n_84_36), .B (n_90_33), .C1 (n_94_31), .C2 (n_100_28) );
AOI211_X1 g_78_39 (.ZN (n_78_39), .A (n_82_37), .B (n_88_34), .C1 (n_92_32), .C2 (n_98_29) );
AOI211_X1 g_76_40 (.ZN (n_76_40), .A (n_80_38), .B (n_86_35), .C1 (n_90_33), .C2 (n_96_30) );
AOI211_X1 g_74_41 (.ZN (n_74_41), .A (n_78_39), .B (n_84_36), .C1 (n_88_34), .C2 (n_94_31) );
AOI211_X1 g_72_42 (.ZN (n_72_42), .A (n_76_40), .B (n_82_37), .C1 (n_86_35), .C2 (n_92_32) );
AOI211_X1 g_70_43 (.ZN (n_70_43), .A (n_74_41), .B (n_80_38), .C1 (n_84_36), .C2 (n_90_33) );
AOI211_X1 g_71_41 (.ZN (n_71_41), .A (n_72_42), .B (n_78_39), .C1 (n_82_37), .C2 (n_88_34) );
AOI211_X1 g_69_42 (.ZN (n_69_42), .A (n_70_43), .B (n_76_40), .C1 (n_80_38), .C2 (n_86_35) );
AOI211_X1 g_67_43 (.ZN (n_67_43), .A (n_71_41), .B (n_74_41), .C1 (n_78_39), .C2 (n_84_36) );
AOI211_X1 g_65_44 (.ZN (n_65_44), .A (n_69_42), .B (n_72_42), .C1 (n_76_40), .C2 (n_82_37) );
AOI211_X1 g_63_45 (.ZN (n_63_45), .A (n_67_43), .B (n_70_43), .C1 (n_74_41), .C2 (n_80_38) );
AOI211_X1 g_61_46 (.ZN (n_61_46), .A (n_65_44), .B (n_71_41), .C1 (n_72_42), .C2 (n_78_39) );
AOI211_X1 g_59_47 (.ZN (n_59_47), .A (n_63_45), .B (n_69_42), .C1 (n_70_43), .C2 (n_76_40) );
AOI211_X1 g_57_48 (.ZN (n_57_48), .A (n_61_46), .B (n_67_43), .C1 (n_71_41), .C2 (n_74_41) );
AOI211_X1 g_55_49 (.ZN (n_55_49), .A (n_59_47), .B (n_65_44), .C1 (n_69_42), .C2 (n_72_42) );
AOI211_X1 g_53_50 (.ZN (n_53_50), .A (n_57_48), .B (n_63_45), .C1 (n_67_43), .C2 (n_70_43) );
AOI211_X1 g_51_51 (.ZN (n_51_51), .A (n_55_49), .B (n_61_46), .C1 (n_65_44), .C2 (n_71_41) );
AOI211_X1 g_49_52 (.ZN (n_49_52), .A (n_53_50), .B (n_59_47), .C1 (n_63_45), .C2 (n_69_42) );
AOI211_X1 g_47_53 (.ZN (n_47_53), .A (n_51_51), .B (n_57_48), .C1 (n_61_46), .C2 (n_67_43) );
AOI211_X1 g_45_54 (.ZN (n_45_54), .A (n_49_52), .B (n_55_49), .C1 (n_59_47), .C2 (n_65_44) );
AOI211_X1 g_43_55 (.ZN (n_43_55), .A (n_47_53), .B (n_53_50), .C1 (n_57_48), .C2 (n_63_45) );
AOI211_X1 g_41_56 (.ZN (n_41_56), .A (n_45_54), .B (n_51_51), .C1 (n_55_49), .C2 (n_61_46) );
AOI211_X1 g_39_57 (.ZN (n_39_57), .A (n_43_55), .B (n_49_52), .C1 (n_53_50), .C2 (n_59_47) );
AOI211_X1 g_37_58 (.ZN (n_37_58), .A (n_41_56), .B (n_47_53), .C1 (n_51_51), .C2 (n_57_48) );
AOI211_X1 g_35_59 (.ZN (n_35_59), .A (n_39_57), .B (n_45_54), .C1 (n_49_52), .C2 (n_55_49) );
AOI211_X1 g_33_60 (.ZN (n_33_60), .A (n_37_58), .B (n_43_55), .C1 (n_47_53), .C2 (n_53_50) );
AOI211_X1 g_31_61 (.ZN (n_31_61), .A (n_35_59), .B (n_41_56), .C1 (n_45_54), .C2 (n_51_51) );
AOI211_X1 g_29_62 (.ZN (n_29_62), .A (n_33_60), .B (n_39_57), .C1 (n_43_55), .C2 (n_49_52) );
AOI211_X1 g_27_63 (.ZN (n_27_63), .A (n_31_61), .B (n_37_58), .C1 (n_41_56), .C2 (n_47_53) );
AOI211_X1 g_25_64 (.ZN (n_25_64), .A (n_29_62), .B (n_35_59), .C1 (n_39_57), .C2 (n_45_54) );
AOI211_X1 g_23_65 (.ZN (n_23_65), .A (n_27_63), .B (n_33_60), .C1 (n_37_58), .C2 (n_43_55) );
AOI211_X1 g_21_66 (.ZN (n_21_66), .A (n_25_64), .B (n_31_61), .C1 (n_35_59), .C2 (n_41_56) );
AOI211_X1 g_19_67 (.ZN (n_19_67), .A (n_23_65), .B (n_29_62), .C1 (n_33_60), .C2 (n_39_57) );
AOI211_X1 g_17_68 (.ZN (n_17_68), .A (n_21_66), .B (n_27_63), .C1 (n_31_61), .C2 (n_37_58) );
AOI211_X1 g_15_69 (.ZN (n_15_69), .A (n_19_67), .B (n_25_64), .C1 (n_29_62), .C2 (n_35_59) );
AOI211_X1 g_13_70 (.ZN (n_13_70), .A (n_17_68), .B (n_23_65), .C1 (n_27_63), .C2 (n_33_60) );
AOI211_X1 g_14_68 (.ZN (n_14_68), .A (n_15_69), .B (n_21_66), .C1 (n_25_64), .C2 (n_31_61) );
AOI211_X1 g_12_69 (.ZN (n_12_69), .A (n_13_70), .B (n_19_67), .C1 (n_23_65), .C2 (n_29_62) );
AOI211_X1 g_13_67 (.ZN (n_13_67), .A (n_14_68), .B (n_17_68), .C1 (n_21_66), .C2 (n_27_63) );
AOI211_X1 g_11_68 (.ZN (n_11_68), .A (n_12_69), .B (n_15_69), .C1 (n_19_67), .C2 (n_25_64) );
AOI211_X1 g_9_69 (.ZN (n_9_69), .A (n_13_67), .B (n_13_70), .C1 (n_17_68), .C2 (n_23_65) );
AOI211_X1 g_8_71 (.ZN (n_8_71), .A (n_11_68), .B (n_14_68), .C1 (n_15_69), .C2 (n_21_66) );
AOI211_X1 g_10_70 (.ZN (n_10_70), .A (n_9_69), .B (n_12_69), .C1 (n_13_70), .C2 (n_19_67) );
AOI211_X1 g_9_72 (.ZN (n_9_72), .A (n_8_71), .B (n_13_67), .C1 (n_14_68), .C2 (n_17_68) );
AOI211_X1 g_8_70 (.ZN (n_8_70), .A (n_10_70), .B (n_11_68), .C1 (n_12_69), .C2 (n_15_69) );
AOI211_X1 g_10_69 (.ZN (n_10_69), .A (n_9_72), .B (n_9_69), .C1 (n_13_67), .C2 (n_13_70) );
AOI211_X1 g_12_68 (.ZN (n_12_68), .A (n_8_70), .B (n_8_71), .C1 (n_11_68), .C2 (n_14_68) );
AOI211_X1 g_14_69 (.ZN (n_14_69), .A (n_10_69), .B (n_10_70), .C1 (n_9_69), .C2 (n_12_69) );
AOI211_X1 g_12_70 (.ZN (n_12_70), .A (n_12_68), .B (n_9_72), .C1 (n_8_71), .C2 (n_13_67) );
AOI211_X1 g_10_71 (.ZN (n_10_71), .A (n_14_69), .B (n_8_70), .C1 (n_10_70), .C2 (n_11_68) );
AOI211_X1 g_9_73 (.ZN (n_9_73), .A (n_12_70), .B (n_10_69), .C1 (n_9_72), .C2 (n_9_69) );
AOI211_X1 g_7_72 (.ZN (n_7_72), .A (n_10_71), .B (n_12_68), .C1 (n_8_70), .C2 (n_8_71) );
AOI211_X1 g_9_71 (.ZN (n_9_71), .A (n_9_73), .B (n_14_69), .C1 (n_10_69), .C2 (n_10_70) );
AOI211_X1 g_11_70 (.ZN (n_11_70), .A (n_7_72), .B (n_12_70), .C1 (n_12_68), .C2 (n_9_72) );
AOI211_X1 g_13_69 (.ZN (n_13_69), .A (n_9_71), .B (n_10_71), .C1 (n_14_69), .C2 (n_8_70) );
AOI211_X1 g_15_68 (.ZN (n_15_68), .A (n_11_70), .B (n_9_73), .C1 (n_12_70), .C2 (n_10_69) );
AOI211_X1 g_17_67 (.ZN (n_17_67), .A (n_13_69), .B (n_7_72), .C1 (n_10_71), .C2 (n_12_68) );
AOI211_X1 g_19_66 (.ZN (n_19_66), .A (n_15_68), .B (n_9_71), .C1 (n_9_73), .C2 (n_14_69) );
AOI211_X1 g_21_65 (.ZN (n_21_65), .A (n_17_67), .B (n_11_70), .C1 (n_7_72), .C2 (n_12_70) );
AOI211_X1 g_23_64 (.ZN (n_23_64), .A (n_19_66), .B (n_13_69), .C1 (n_9_71), .C2 (n_10_71) );
AOI211_X1 g_25_63 (.ZN (n_25_63), .A (n_21_65), .B (n_15_68), .C1 (n_11_70), .C2 (n_9_73) );
AOI211_X1 g_27_62 (.ZN (n_27_62), .A (n_23_64), .B (n_17_67), .C1 (n_13_69), .C2 (n_7_72) );
AOI211_X1 g_29_61 (.ZN (n_29_61), .A (n_25_63), .B (n_19_66), .C1 (n_15_68), .C2 (n_9_71) );
AOI211_X1 g_31_60 (.ZN (n_31_60), .A (n_27_62), .B (n_21_65), .C1 (n_17_67), .C2 (n_11_70) );
AOI211_X1 g_33_59 (.ZN (n_33_59), .A (n_29_61), .B (n_23_64), .C1 (n_19_66), .C2 (n_13_69) );
AOI211_X1 g_35_58 (.ZN (n_35_58), .A (n_31_60), .B (n_25_63), .C1 (n_21_65), .C2 (n_15_68) );
AOI211_X1 g_34_60 (.ZN (n_34_60), .A (n_33_59), .B (n_27_62), .C1 (n_23_64), .C2 (n_17_67) );
AOI211_X1 g_36_59 (.ZN (n_36_59), .A (n_35_58), .B (n_29_61), .C1 (n_25_63), .C2 (n_19_66) );
AOI211_X1 g_38_58 (.ZN (n_38_58), .A (n_34_60), .B (n_31_60), .C1 (n_27_62), .C2 (n_21_65) );
AOI211_X1 g_40_57 (.ZN (n_40_57), .A (n_36_59), .B (n_33_59), .C1 (n_29_61), .C2 (n_23_64) );
AOI211_X1 g_42_56 (.ZN (n_42_56), .A (n_38_58), .B (n_35_58), .C1 (n_31_60), .C2 (n_25_63) );
AOI211_X1 g_44_55 (.ZN (n_44_55), .A (n_40_57), .B (n_34_60), .C1 (n_33_59), .C2 (n_27_62) );
AOI211_X1 g_46_54 (.ZN (n_46_54), .A (n_42_56), .B (n_36_59), .C1 (n_35_58), .C2 (n_29_61) );
AOI211_X1 g_48_53 (.ZN (n_48_53), .A (n_44_55), .B (n_38_58), .C1 (n_34_60), .C2 (n_31_60) );
AOI211_X1 g_50_52 (.ZN (n_50_52), .A (n_46_54), .B (n_40_57), .C1 (n_36_59), .C2 (n_33_59) );
AOI211_X1 g_49_54 (.ZN (n_49_54), .A (n_48_53), .B (n_42_56), .C1 (n_38_58), .C2 (n_35_58) );
AOI211_X1 g_48_52 (.ZN (n_48_52), .A (n_50_52), .B (n_44_55), .C1 (n_40_57), .C2 (n_34_60) );
AOI211_X1 g_50_51 (.ZN (n_50_51), .A (n_49_54), .B (n_46_54), .C1 (n_42_56), .C2 (n_36_59) );
AOI211_X1 g_52_50 (.ZN (n_52_50), .A (n_48_52), .B (n_48_53), .C1 (n_44_55), .C2 (n_38_58) );
AOI211_X1 g_54_49 (.ZN (n_54_49), .A (n_50_51), .B (n_50_52), .C1 (n_46_54), .C2 (n_40_57) );
AOI211_X1 g_53_51 (.ZN (n_53_51), .A (n_52_50), .B (n_49_54), .C1 (n_48_53), .C2 (n_42_56) );
AOI211_X1 g_55_50 (.ZN (n_55_50), .A (n_54_49), .B (n_48_52), .C1 (n_50_52), .C2 (n_44_55) );
AOI211_X1 g_57_49 (.ZN (n_57_49), .A (n_53_51), .B (n_50_51), .C1 (n_49_54), .C2 (n_46_54) );
AOI211_X1 g_59_48 (.ZN (n_59_48), .A (n_55_50), .B (n_52_50), .C1 (n_48_52), .C2 (n_48_53) );
AOI211_X1 g_61_47 (.ZN (n_61_47), .A (n_57_49), .B (n_54_49), .C1 (n_50_51), .C2 (n_50_52) );
AOI211_X1 g_62_45 (.ZN (n_62_45), .A (n_59_48), .B (n_53_51), .C1 (n_52_50), .C2 (n_49_54) );
AOI211_X1 g_64_44 (.ZN (n_64_44), .A (n_61_47), .B (n_55_50), .C1 (n_54_49), .C2 (n_48_52) );
AOI211_X1 g_63_46 (.ZN (n_63_46), .A (n_62_45), .B (n_57_49), .C1 (n_53_51), .C2 (n_50_51) );
AOI211_X1 g_65_45 (.ZN (n_65_45), .A (n_64_44), .B (n_59_48), .C1 (n_55_50), .C2 (n_52_50) );
AOI211_X1 g_67_44 (.ZN (n_67_44), .A (n_63_46), .B (n_61_47), .C1 (n_57_49), .C2 (n_54_49) );
AOI211_X1 g_69_43 (.ZN (n_69_43), .A (n_65_45), .B (n_62_45), .C1 (n_59_48), .C2 (n_53_51) );
AOI211_X1 g_71_42 (.ZN (n_71_42), .A (n_67_44), .B (n_64_44), .C1 (n_61_47), .C2 (n_55_50) );
AOI211_X1 g_73_41 (.ZN (n_73_41), .A (n_69_43), .B (n_63_46), .C1 (n_62_45), .C2 (n_57_49) );
AOI211_X1 g_75_40 (.ZN (n_75_40), .A (n_71_42), .B (n_65_45), .C1 (n_64_44), .C2 (n_59_48) );
AOI211_X1 g_77_39 (.ZN (n_77_39), .A (n_73_41), .B (n_67_44), .C1 (n_63_46), .C2 (n_61_47) );
AOI211_X1 g_79_38 (.ZN (n_79_38), .A (n_75_40), .B (n_69_43), .C1 (n_65_45), .C2 (n_62_45) );
AOI211_X1 g_81_37 (.ZN (n_81_37), .A (n_77_39), .B (n_71_42), .C1 (n_67_44), .C2 (n_64_44) );
AOI211_X1 g_83_36 (.ZN (n_83_36), .A (n_79_38), .B (n_73_41), .C1 (n_69_43), .C2 (n_63_46) );
AOI211_X1 g_85_35 (.ZN (n_85_35), .A (n_81_37), .B (n_75_40), .C1 (n_71_42), .C2 (n_65_45) );
AOI211_X1 g_87_34 (.ZN (n_87_34), .A (n_83_36), .B (n_77_39), .C1 (n_73_41), .C2 (n_67_44) );
AOI211_X1 g_89_33 (.ZN (n_89_33), .A (n_85_35), .B (n_79_38), .C1 (n_75_40), .C2 (n_69_43) );
AOI211_X1 g_91_32 (.ZN (n_91_32), .A (n_87_34), .B (n_81_37), .C1 (n_77_39), .C2 (n_71_42) );
AOI211_X1 g_93_31 (.ZN (n_93_31), .A (n_89_33), .B (n_83_36), .C1 (n_79_38), .C2 (n_73_41) );
AOI211_X1 g_95_30 (.ZN (n_95_30), .A (n_91_32), .B (n_85_35), .C1 (n_81_37), .C2 (n_75_40) );
AOI211_X1 g_97_29 (.ZN (n_97_29), .A (n_93_31), .B (n_87_34), .C1 (n_83_36), .C2 (n_77_39) );
AOI211_X1 g_99_30 (.ZN (n_99_30), .A (n_95_30), .B (n_89_33), .C1 (n_85_35), .C2 (n_79_38) );
AOI211_X1 g_97_31 (.ZN (n_97_31), .A (n_97_29), .B (n_91_32), .C1 (n_87_34), .C2 (n_81_37) );
AOI211_X1 g_95_32 (.ZN (n_95_32), .A (n_99_30), .B (n_93_31), .C1 (n_89_33), .C2 (n_83_36) );
AOI211_X1 g_93_33 (.ZN (n_93_33), .A (n_97_31), .B (n_95_30), .C1 (n_91_32), .C2 (n_85_35) );
AOI211_X1 g_91_34 (.ZN (n_91_34), .A (n_95_32), .B (n_97_29), .C1 (n_93_31), .C2 (n_87_34) );
AOI211_X1 g_89_35 (.ZN (n_89_35), .A (n_93_33), .B (n_99_30), .C1 (n_95_30), .C2 (n_89_33) );
AOI211_X1 g_87_36 (.ZN (n_87_36), .A (n_91_34), .B (n_97_31), .C1 (n_97_29), .C2 (n_91_32) );
AOI211_X1 g_85_37 (.ZN (n_85_37), .A (n_89_35), .B (n_95_32), .C1 (n_99_30), .C2 (n_93_31) );
AOI211_X1 g_83_38 (.ZN (n_83_38), .A (n_87_36), .B (n_93_33), .C1 (n_97_31), .C2 (n_95_30) );
AOI211_X1 g_81_39 (.ZN (n_81_39), .A (n_85_37), .B (n_91_34), .C1 (n_95_32), .C2 (n_97_29) );
AOI211_X1 g_79_40 (.ZN (n_79_40), .A (n_83_38), .B (n_89_35), .C1 (n_93_33), .C2 (n_99_30) );
AOI211_X1 g_77_41 (.ZN (n_77_41), .A (n_81_39), .B (n_87_36), .C1 (n_91_34), .C2 (n_97_31) );
AOI211_X1 g_75_42 (.ZN (n_75_42), .A (n_79_40), .B (n_85_37), .C1 (n_89_35), .C2 (n_95_32) );
AOI211_X1 g_73_43 (.ZN (n_73_43), .A (n_77_41), .B (n_83_38), .C1 (n_87_36), .C2 (n_93_33) );
AOI211_X1 g_71_44 (.ZN (n_71_44), .A (n_75_42), .B (n_81_39), .C1 (n_85_37), .C2 (n_91_34) );
AOI211_X1 g_69_45 (.ZN (n_69_45), .A (n_73_43), .B (n_79_40), .C1 (n_83_38), .C2 (n_89_35) );
AOI211_X1 g_67_46 (.ZN (n_67_46), .A (n_71_44), .B (n_77_41), .C1 (n_81_39), .C2 (n_87_36) );
AOI211_X1 g_68_44 (.ZN (n_68_44), .A (n_69_45), .B (n_75_42), .C1 (n_79_40), .C2 (n_85_37) );
AOI211_X1 g_66_45 (.ZN (n_66_45), .A (n_67_46), .B (n_73_43), .C1 (n_77_41), .C2 (n_83_38) );
AOI211_X1 g_64_46 (.ZN (n_64_46), .A (n_68_44), .B (n_71_44), .C1 (n_75_42), .C2 (n_81_39) );
AOI211_X1 g_62_47 (.ZN (n_62_47), .A (n_66_45), .B (n_69_45), .C1 (n_73_43), .C2 (n_79_40) );
AOI211_X1 g_60_48 (.ZN (n_60_48), .A (n_64_46), .B (n_67_46), .C1 (n_71_44), .C2 (n_77_41) );
AOI211_X1 g_58_49 (.ZN (n_58_49), .A (n_62_47), .B (n_68_44), .C1 (n_69_45), .C2 (n_75_42) );
AOI211_X1 g_56_50 (.ZN (n_56_50), .A (n_60_48), .B (n_66_45), .C1 (n_67_46), .C2 (n_73_43) );
AOI211_X1 g_54_51 (.ZN (n_54_51), .A (n_58_49), .B (n_64_46), .C1 (n_68_44), .C2 (n_71_44) );
AOI211_X1 g_52_52 (.ZN (n_52_52), .A (n_56_50), .B (n_62_47), .C1 (n_66_45), .C2 (n_69_45) );
AOI211_X1 g_50_53 (.ZN (n_50_53), .A (n_54_51), .B (n_60_48), .C1 (n_64_46), .C2 (n_67_46) );
AOI211_X1 g_48_54 (.ZN (n_48_54), .A (n_52_52), .B (n_58_49), .C1 (n_62_47), .C2 (n_68_44) );
AOI211_X1 g_46_53 (.ZN (n_46_53), .A (n_50_53), .B (n_56_50), .C1 (n_60_48), .C2 (n_66_45) );
AOI211_X1 g_44_54 (.ZN (n_44_54), .A (n_48_54), .B (n_54_51), .C1 (n_58_49), .C2 (n_64_46) );
AOI211_X1 g_42_55 (.ZN (n_42_55), .A (n_46_53), .B (n_52_52), .C1 (n_56_50), .C2 (n_62_47) );
AOI211_X1 g_40_56 (.ZN (n_40_56), .A (n_44_54), .B (n_50_53), .C1 (n_54_51), .C2 (n_60_48) );
AOI211_X1 g_38_57 (.ZN (n_38_57), .A (n_42_55), .B (n_48_54), .C1 (n_52_52), .C2 (n_58_49) );
AOI211_X1 g_36_58 (.ZN (n_36_58), .A (n_40_56), .B (n_46_53), .C1 (n_50_53), .C2 (n_56_50) );
AOI211_X1 g_34_59 (.ZN (n_34_59), .A (n_38_57), .B (n_44_54), .C1 (n_48_54), .C2 (n_54_51) );
AOI211_X1 g_32_60 (.ZN (n_32_60), .A (n_36_58), .B (n_42_55), .C1 (n_46_53), .C2 (n_52_52) );
AOI211_X1 g_30_61 (.ZN (n_30_61), .A (n_34_59), .B (n_40_56), .C1 (n_44_54), .C2 (n_50_53) );
AOI211_X1 g_28_62 (.ZN (n_28_62), .A (n_32_60), .B (n_38_57), .C1 (n_42_55), .C2 (n_48_54) );
AOI211_X1 g_27_64 (.ZN (n_27_64), .A (n_30_61), .B (n_36_58), .C1 (n_40_56), .C2 (n_46_53) );
AOI211_X1 g_29_63 (.ZN (n_29_63), .A (n_28_62), .B (n_34_59), .C1 (n_38_57), .C2 (n_44_54) );
AOI211_X1 g_31_62 (.ZN (n_31_62), .A (n_27_64), .B (n_32_60), .C1 (n_36_58), .C2 (n_42_55) );
AOI211_X1 g_33_61 (.ZN (n_33_61), .A (n_29_63), .B (n_30_61), .C1 (n_34_59), .C2 (n_40_56) );
AOI211_X1 g_35_60 (.ZN (n_35_60), .A (n_31_62), .B (n_28_62), .C1 (n_32_60), .C2 (n_38_57) );
AOI211_X1 g_37_59 (.ZN (n_37_59), .A (n_33_61), .B (n_27_64), .C1 (n_30_61), .C2 (n_36_58) );
AOI211_X1 g_39_58 (.ZN (n_39_58), .A (n_35_60), .B (n_29_63), .C1 (n_28_62), .C2 (n_34_59) );
AOI211_X1 g_41_57 (.ZN (n_41_57), .A (n_37_59), .B (n_31_62), .C1 (n_27_64), .C2 (n_32_60) );
AOI211_X1 g_43_56 (.ZN (n_43_56), .A (n_39_58), .B (n_33_61), .C1 (n_29_63), .C2 (n_30_61) );
AOI211_X1 g_45_55 (.ZN (n_45_55), .A (n_41_57), .B (n_35_60), .C1 (n_31_62), .C2 (n_28_62) );
AOI211_X1 g_47_54 (.ZN (n_47_54), .A (n_43_56), .B (n_37_59), .C1 (n_33_61), .C2 (n_27_64) );
AOI211_X1 g_49_53 (.ZN (n_49_53), .A (n_45_55), .B (n_39_58), .C1 (n_35_60), .C2 (n_29_63) );
AOI211_X1 g_51_52 (.ZN (n_51_52), .A (n_47_54), .B (n_41_57), .C1 (n_37_59), .C2 (n_31_62) );
AOI211_X1 g_50_54 (.ZN (n_50_54), .A (n_49_53), .B (n_43_56), .C1 (n_39_58), .C2 (n_33_61) );
AOI211_X1 g_52_53 (.ZN (n_52_53), .A (n_51_52), .B (n_45_55), .C1 (n_41_57), .C2 (n_35_60) );
AOI211_X1 g_54_52 (.ZN (n_54_52), .A (n_50_54), .B (n_47_54), .C1 (n_43_56), .C2 (n_37_59) );
AOI211_X1 g_56_51 (.ZN (n_56_51), .A (n_52_53), .B (n_49_53), .C1 (n_45_55), .C2 (n_39_58) );
AOI211_X1 g_58_50 (.ZN (n_58_50), .A (n_54_52), .B (n_51_52), .C1 (n_47_54), .C2 (n_41_57) );
AOI211_X1 g_60_49 (.ZN (n_60_49), .A (n_56_51), .B (n_50_54), .C1 (n_49_53), .C2 (n_43_56) );
AOI211_X1 g_62_48 (.ZN (n_62_48), .A (n_58_50), .B (n_52_53), .C1 (n_51_52), .C2 (n_45_55) );
AOI211_X1 g_64_47 (.ZN (n_64_47), .A (n_60_49), .B (n_54_52), .C1 (n_50_54), .C2 (n_47_54) );
AOI211_X1 g_66_46 (.ZN (n_66_46), .A (n_62_48), .B (n_56_51), .C1 (n_52_53), .C2 (n_49_53) );
AOI211_X1 g_68_45 (.ZN (n_68_45), .A (n_64_47), .B (n_58_50), .C1 (n_54_52), .C2 (n_51_52) );
AOI211_X1 g_70_44 (.ZN (n_70_44), .A (n_66_46), .B (n_60_49), .C1 (n_56_51), .C2 (n_50_54) );
AOI211_X1 g_72_43 (.ZN (n_72_43), .A (n_68_45), .B (n_62_48), .C1 (n_58_50), .C2 (n_52_53) );
AOI211_X1 g_74_42 (.ZN (n_74_42), .A (n_70_44), .B (n_64_47), .C1 (n_60_49), .C2 (n_54_52) );
AOI211_X1 g_76_41 (.ZN (n_76_41), .A (n_72_43), .B (n_66_46), .C1 (n_62_48), .C2 (n_56_51) );
AOI211_X1 g_78_40 (.ZN (n_78_40), .A (n_74_42), .B (n_68_45), .C1 (n_64_47), .C2 (n_58_50) );
AOI211_X1 g_80_39 (.ZN (n_80_39), .A (n_76_41), .B (n_70_44), .C1 (n_66_46), .C2 (n_60_49) );
AOI211_X1 g_82_38 (.ZN (n_82_38), .A (n_78_40), .B (n_72_43), .C1 (n_68_45), .C2 (n_62_48) );
AOI211_X1 g_84_37 (.ZN (n_84_37), .A (n_80_39), .B (n_74_42), .C1 (n_70_44), .C2 (n_64_47) );
AOI211_X1 g_86_36 (.ZN (n_86_36), .A (n_82_38), .B (n_76_41), .C1 (n_72_43), .C2 (n_66_46) );
AOI211_X1 g_88_35 (.ZN (n_88_35), .A (n_84_37), .B (n_78_40), .C1 (n_74_42), .C2 (n_68_45) );
AOI211_X1 g_90_34 (.ZN (n_90_34), .A (n_86_36), .B (n_80_39), .C1 (n_76_41), .C2 (n_70_44) );
AOI211_X1 g_92_33 (.ZN (n_92_33), .A (n_88_35), .B (n_82_38), .C1 (n_78_40), .C2 (n_72_43) );
AOI211_X1 g_94_32 (.ZN (n_94_32), .A (n_90_34), .B (n_84_37), .C1 (n_80_39), .C2 (n_74_42) );
AOI211_X1 g_96_31 (.ZN (n_96_31), .A (n_92_33), .B (n_86_36), .C1 (n_82_38), .C2 (n_76_41) );
AOI211_X1 g_97_33 (.ZN (n_97_33), .A (n_94_32), .B (n_88_35), .C1 (n_84_37), .C2 (n_78_40) );
AOI211_X1 g_98_31 (.ZN (n_98_31), .A (n_96_31), .B (n_90_34), .C1 (n_86_36), .C2 (n_80_39) );
AOI211_X1 g_99_29 (.ZN (n_99_29), .A (n_97_33), .B (n_92_33), .C1 (n_88_35), .C2 (n_82_38) );
AOI211_X1 g_100_31 (.ZN (n_100_31), .A (n_98_31), .B (n_94_32), .C1 (n_90_34), .C2 (n_84_37) );
AOI211_X1 g_99_33 (.ZN (n_99_33), .A (n_99_29), .B (n_96_31), .C1 (n_92_33), .C2 (n_86_36) );
AOI211_X1 g_100_35 (.ZN (n_100_35), .A (n_100_31), .B (n_97_33), .C1 (n_94_32), .C2 (n_88_35) );
AOI211_X1 g_98_34 (.ZN (n_98_34), .A (n_99_33), .B (n_98_31), .C1 (n_96_31), .C2 (n_90_34) );
AOI211_X1 g_100_33 (.ZN (n_100_33), .A (n_100_35), .B (n_99_29), .C1 (n_97_33), .C2 (n_92_33) );
AOI211_X1 g_99_31 (.ZN (n_99_31), .A (n_98_34), .B (n_100_31), .C1 (n_98_31), .C2 (n_94_32) );
AOI211_X1 g_97_30 (.ZN (n_97_30), .A (n_100_33), .B (n_99_33), .C1 (n_99_29), .C2 (n_96_31) );
AOI211_X1 g_98_32 (.ZN (n_98_32), .A (n_99_31), .B (n_100_35), .C1 (n_100_31), .C2 (n_97_33) );
AOI211_X1 g_96_33 (.ZN (n_96_33), .A (n_97_30), .B (n_98_34), .C1 (n_99_33), .C2 (n_98_31) );
AOI211_X1 g_95_31 (.ZN (n_95_31), .A (n_98_32), .B (n_100_33), .C1 (n_100_35), .C2 (n_99_29) );
AOI211_X1 g_97_32 (.ZN (n_97_32), .A (n_96_33), .B (n_99_31), .C1 (n_98_34), .C2 (n_100_31) );
AOI211_X1 g_95_33 (.ZN (n_95_33), .A (n_95_31), .B (n_97_30), .C1 (n_100_33), .C2 (n_99_33) );
AOI211_X1 g_93_32 (.ZN (n_93_32), .A (n_97_32), .B (n_98_32), .C1 (n_99_31), .C2 (n_100_35) );
AOI211_X1 g_91_33 (.ZN (n_91_33), .A (n_95_33), .B (n_96_33), .C1 (n_97_30), .C2 (n_98_34) );
AOI211_X1 g_89_34 (.ZN (n_89_34), .A (n_93_32), .B (n_95_31), .C1 (n_98_32), .C2 (n_100_33) );
AOI211_X1 g_87_35 (.ZN (n_87_35), .A (n_91_33), .B (n_97_32), .C1 (n_96_33), .C2 (n_99_31) );
AOI211_X1 g_85_36 (.ZN (n_85_36), .A (n_89_34), .B (n_95_33), .C1 (n_95_31), .C2 (n_97_30) );
AOI211_X1 g_84_38 (.ZN (n_84_38), .A (n_87_35), .B (n_93_32), .C1 (n_97_32), .C2 (n_98_32) );
AOI211_X1 g_86_37 (.ZN (n_86_37), .A (n_85_36), .B (n_91_33), .C1 (n_95_33), .C2 (n_96_33) );
AOI211_X1 g_88_36 (.ZN (n_88_36), .A (n_84_38), .B (n_89_34), .C1 (n_93_32), .C2 (n_95_31) );
AOI211_X1 g_90_35 (.ZN (n_90_35), .A (n_86_37), .B (n_87_35), .C1 (n_91_33), .C2 (n_97_32) );
AOI211_X1 g_92_34 (.ZN (n_92_34), .A (n_88_36), .B (n_85_36), .C1 (n_89_34), .C2 (n_95_33) );
AOI211_X1 g_94_33 (.ZN (n_94_33), .A (n_90_35), .B (n_84_38), .C1 (n_87_35), .C2 (n_93_32) );
AOI211_X1 g_96_32 (.ZN (n_96_32), .A (n_92_34), .B (n_86_37), .C1 (n_85_36), .C2 (n_91_33) );
AOI211_X1 g_95_34 (.ZN (n_95_34), .A (n_94_33), .B (n_88_36), .C1 (n_84_38), .C2 (n_89_34) );
AOI211_X1 g_93_35 (.ZN (n_93_35), .A (n_96_32), .B (n_90_35), .C1 (n_86_37), .C2 (n_87_35) );
AOI211_X1 g_91_36 (.ZN (n_91_36), .A (n_95_34), .B (n_92_34), .C1 (n_88_36), .C2 (n_85_36) );
AOI211_X1 g_89_37 (.ZN (n_89_37), .A (n_93_35), .B (n_94_33), .C1 (n_90_35), .C2 (n_84_38) );
AOI211_X1 g_87_38 (.ZN (n_87_38), .A (n_91_36), .B (n_96_32), .C1 (n_92_34), .C2 (n_86_37) );
AOI211_X1 g_85_39 (.ZN (n_85_39), .A (n_89_37), .B (n_95_34), .C1 (n_94_33), .C2 (n_88_36) );
AOI211_X1 g_83_40 (.ZN (n_83_40), .A (n_87_38), .B (n_93_35), .C1 (n_96_32), .C2 (n_90_35) );
AOI211_X1 g_81_41 (.ZN (n_81_41), .A (n_85_39), .B (n_91_36), .C1 (n_95_34), .C2 (n_92_34) );
AOI211_X1 g_82_39 (.ZN (n_82_39), .A (n_83_40), .B (n_89_37), .C1 (n_93_35), .C2 (n_94_33) );
AOI211_X1 g_80_40 (.ZN (n_80_40), .A (n_81_41), .B (n_87_38), .C1 (n_91_36), .C2 (n_96_32) );
AOI211_X1 g_78_41 (.ZN (n_78_41), .A (n_82_39), .B (n_85_39), .C1 (n_89_37), .C2 (n_95_34) );
AOI211_X1 g_76_42 (.ZN (n_76_42), .A (n_80_40), .B (n_83_40), .C1 (n_87_38), .C2 (n_93_35) );
AOI211_X1 g_77_40 (.ZN (n_77_40), .A (n_78_41), .B (n_81_41), .C1 (n_85_39), .C2 (n_91_36) );
AOI211_X1 g_75_41 (.ZN (n_75_41), .A (n_76_42), .B (n_82_39), .C1 (n_83_40), .C2 (n_89_37) );
AOI211_X1 g_73_42 (.ZN (n_73_42), .A (n_77_40), .B (n_80_40), .C1 (n_81_41), .C2 (n_87_38) );
AOI211_X1 g_71_43 (.ZN (n_71_43), .A (n_75_41), .B (n_78_41), .C1 (n_82_39), .C2 (n_85_39) );
AOI211_X1 g_69_44 (.ZN (n_69_44), .A (n_73_42), .B (n_76_42), .C1 (n_80_40), .C2 (n_83_40) );
AOI211_X1 g_67_45 (.ZN (n_67_45), .A (n_71_43), .B (n_77_40), .C1 (n_78_41), .C2 (n_81_41) );
AOI211_X1 g_65_46 (.ZN (n_65_46), .A (n_69_44), .B (n_75_41), .C1 (n_76_42), .C2 (n_82_39) );
AOI211_X1 g_63_47 (.ZN (n_63_47), .A (n_67_45), .B (n_73_42), .C1 (n_77_40), .C2 (n_80_40) );
AOI211_X1 g_61_48 (.ZN (n_61_48), .A (n_65_46), .B (n_71_43), .C1 (n_75_41), .C2 (n_78_41) );
AOI211_X1 g_59_49 (.ZN (n_59_49), .A (n_63_47), .B (n_69_44), .C1 (n_73_42), .C2 (n_76_42) );
AOI211_X1 g_57_50 (.ZN (n_57_50), .A (n_61_48), .B (n_67_45), .C1 (n_71_43), .C2 (n_77_40) );
AOI211_X1 g_55_51 (.ZN (n_55_51), .A (n_59_49), .B (n_65_46), .C1 (n_69_44), .C2 (n_75_41) );
AOI211_X1 g_53_52 (.ZN (n_53_52), .A (n_57_50), .B (n_63_47), .C1 (n_67_45), .C2 (n_73_42) );
AOI211_X1 g_51_53 (.ZN (n_51_53), .A (n_55_51), .B (n_61_48), .C1 (n_65_46), .C2 (n_71_43) );
AOI211_X1 g_50_55 (.ZN (n_50_55), .A (n_53_52), .B (n_59_49), .C1 (n_63_47), .C2 (n_69_44) );
AOI211_X1 g_52_54 (.ZN (n_52_54), .A (n_51_53), .B (n_57_50), .C1 (n_61_48), .C2 (n_67_45) );
AOI211_X1 g_54_53 (.ZN (n_54_53), .A (n_50_55), .B (n_55_51), .C1 (n_59_49), .C2 (n_65_46) );
AOI211_X1 g_56_52 (.ZN (n_56_52), .A (n_52_54), .B (n_53_52), .C1 (n_57_50), .C2 (n_63_47) );
AOI211_X1 g_58_51 (.ZN (n_58_51), .A (n_54_53), .B (n_51_53), .C1 (n_55_51), .C2 (n_61_48) );
AOI211_X1 g_60_50 (.ZN (n_60_50), .A (n_56_52), .B (n_50_55), .C1 (n_53_52), .C2 (n_59_49) );
AOI211_X1 g_62_49 (.ZN (n_62_49), .A (n_58_51), .B (n_52_54), .C1 (n_51_53), .C2 (n_57_50) );
AOI211_X1 g_64_48 (.ZN (n_64_48), .A (n_60_50), .B (n_54_53), .C1 (n_50_55), .C2 (n_55_51) );
AOI211_X1 g_66_47 (.ZN (n_66_47), .A (n_62_49), .B (n_56_52), .C1 (n_52_54), .C2 (n_53_52) );
AOI211_X1 g_68_46 (.ZN (n_68_46), .A (n_64_48), .B (n_58_51), .C1 (n_54_53), .C2 (n_51_53) );
AOI211_X1 g_70_45 (.ZN (n_70_45), .A (n_66_47), .B (n_60_50), .C1 (n_56_52), .C2 (n_50_55) );
AOI211_X1 g_72_44 (.ZN (n_72_44), .A (n_68_46), .B (n_62_49), .C1 (n_58_51), .C2 (n_52_54) );
AOI211_X1 g_74_43 (.ZN (n_74_43), .A (n_70_45), .B (n_64_48), .C1 (n_60_50), .C2 (n_54_53) );
AOI211_X1 g_73_45 (.ZN (n_73_45), .A (n_72_44), .B (n_66_47), .C1 (n_62_49), .C2 (n_56_52) );
AOI211_X1 g_75_44 (.ZN (n_75_44), .A (n_74_43), .B (n_68_46), .C1 (n_64_48), .C2 (n_58_51) );
AOI211_X1 g_77_43 (.ZN (n_77_43), .A (n_73_45), .B (n_70_45), .C1 (n_66_47), .C2 (n_60_50) );
AOI211_X1 g_79_42 (.ZN (n_79_42), .A (n_75_44), .B (n_72_44), .C1 (n_68_46), .C2 (n_62_49) );
AOI211_X1 g_78_44 (.ZN (n_78_44), .A (n_77_43), .B (n_74_43), .C1 (n_70_45), .C2 (n_64_48) );
AOI211_X1 g_77_42 (.ZN (n_77_42), .A (n_79_42), .B (n_73_45), .C1 (n_72_44), .C2 (n_66_47) );
AOI211_X1 g_79_41 (.ZN (n_79_41), .A (n_78_44), .B (n_75_44), .C1 (n_74_43), .C2 (n_68_46) );
AOI211_X1 g_81_40 (.ZN (n_81_40), .A (n_77_42), .B (n_77_43), .C1 (n_73_45), .C2 (n_70_45) );
AOI211_X1 g_83_39 (.ZN (n_83_39), .A (n_79_41), .B (n_79_42), .C1 (n_75_44), .C2 (n_72_44) );
AOI211_X1 g_85_38 (.ZN (n_85_38), .A (n_81_40), .B (n_78_44), .C1 (n_77_43), .C2 (n_74_43) );
AOI211_X1 g_87_37 (.ZN (n_87_37), .A (n_83_39), .B (n_77_42), .C1 (n_79_42), .C2 (n_73_45) );
AOI211_X1 g_89_36 (.ZN (n_89_36), .A (n_85_38), .B (n_79_41), .C1 (n_78_44), .C2 (n_75_44) );
AOI211_X1 g_91_35 (.ZN (n_91_35), .A (n_87_37), .B (n_81_40), .C1 (n_77_42), .C2 (n_77_43) );
AOI211_X1 g_93_34 (.ZN (n_93_34), .A (n_89_36), .B (n_83_39), .C1 (n_79_41), .C2 (n_79_42) );
AOI211_X1 g_92_36 (.ZN (n_92_36), .A (n_91_35), .B (n_85_38), .C1 (n_81_40), .C2 (n_78_44) );
AOI211_X1 g_94_35 (.ZN (n_94_35), .A (n_93_34), .B (n_87_37), .C1 (n_83_39), .C2 (n_77_42) );
AOI211_X1 g_96_34 (.ZN (n_96_34), .A (n_92_36), .B (n_89_36), .C1 (n_85_38), .C2 (n_79_41) );
AOI211_X1 g_98_33 (.ZN (n_98_33), .A (n_94_35), .B (n_91_35), .C1 (n_87_37), .C2 (n_81_40) );
AOI211_X1 g_100_32 (.ZN (n_100_32), .A (n_96_34), .B (n_93_34), .C1 (n_89_36), .C2 (n_83_39) );
AOI211_X1 g_99_34 (.ZN (n_99_34), .A (n_98_33), .B (n_92_36), .C1 (n_91_35), .C2 (n_85_38) );
AOI211_X1 g_97_35 (.ZN (n_97_35), .A (n_100_32), .B (n_94_35), .C1 (n_93_34), .C2 (n_87_37) );
AOI211_X1 g_95_36 (.ZN (n_95_36), .A (n_99_34), .B (n_96_34), .C1 (n_92_36), .C2 (n_89_36) );
AOI211_X1 g_94_34 (.ZN (n_94_34), .A (n_97_35), .B (n_98_33), .C1 (n_94_35), .C2 (n_91_35) );
AOI211_X1 g_92_35 (.ZN (n_92_35), .A (n_95_36), .B (n_100_32), .C1 (n_96_34), .C2 (n_93_34) );
AOI211_X1 g_90_36 (.ZN (n_90_36), .A (n_94_34), .B (n_99_34), .C1 (n_98_33), .C2 (n_92_36) );
AOI211_X1 g_88_37 (.ZN (n_88_37), .A (n_92_35), .B (n_97_35), .C1 (n_100_32), .C2 (n_94_35) );
AOI211_X1 g_86_38 (.ZN (n_86_38), .A (n_90_36), .B (n_95_36), .C1 (n_99_34), .C2 (n_96_34) );
AOI211_X1 g_84_39 (.ZN (n_84_39), .A (n_88_37), .B (n_94_34), .C1 (n_97_35), .C2 (n_98_33) );
AOI211_X1 g_82_40 (.ZN (n_82_40), .A (n_86_38), .B (n_92_35), .C1 (n_95_36), .C2 (n_100_32) );
AOI211_X1 g_80_41 (.ZN (n_80_41), .A (n_84_39), .B (n_90_36), .C1 (n_94_34), .C2 (n_99_34) );
AOI211_X1 g_78_42 (.ZN (n_78_42), .A (n_82_40), .B (n_88_37), .C1 (n_92_35), .C2 (n_97_35) );
AOI211_X1 g_76_43 (.ZN (n_76_43), .A (n_80_41), .B (n_86_38), .C1 (n_90_36), .C2 (n_95_36) );
AOI211_X1 g_74_44 (.ZN (n_74_44), .A (n_78_42), .B (n_84_39), .C1 (n_88_37), .C2 (n_94_34) );
AOI211_X1 g_72_45 (.ZN (n_72_45), .A (n_76_43), .B (n_82_40), .C1 (n_86_38), .C2 (n_92_35) );
AOI211_X1 g_70_46 (.ZN (n_70_46), .A (n_74_44), .B (n_80_41), .C1 (n_84_39), .C2 (n_90_36) );
AOI211_X1 g_68_47 (.ZN (n_68_47), .A (n_72_45), .B (n_78_42), .C1 (n_82_40), .C2 (n_88_37) );
AOI211_X1 g_66_48 (.ZN (n_66_48), .A (n_70_46), .B (n_76_43), .C1 (n_80_41), .C2 (n_86_38) );
AOI211_X1 g_64_49 (.ZN (n_64_49), .A (n_68_47), .B (n_74_44), .C1 (n_78_42), .C2 (n_84_39) );
AOI211_X1 g_65_47 (.ZN (n_65_47), .A (n_66_48), .B (n_72_45), .C1 (n_76_43), .C2 (n_82_40) );
AOI211_X1 g_63_48 (.ZN (n_63_48), .A (n_64_49), .B (n_70_46), .C1 (n_74_44), .C2 (n_80_41) );
AOI211_X1 g_61_49 (.ZN (n_61_49), .A (n_65_47), .B (n_68_47), .C1 (n_72_45), .C2 (n_78_42) );
AOI211_X1 g_59_50 (.ZN (n_59_50), .A (n_63_48), .B (n_66_48), .C1 (n_70_46), .C2 (n_76_43) );
AOI211_X1 g_57_51 (.ZN (n_57_51), .A (n_61_49), .B (n_64_49), .C1 (n_68_47), .C2 (n_74_44) );
AOI211_X1 g_55_52 (.ZN (n_55_52), .A (n_59_50), .B (n_65_47), .C1 (n_66_48), .C2 (n_72_45) );
AOI211_X1 g_53_53 (.ZN (n_53_53), .A (n_57_51), .B (n_63_48), .C1 (n_64_49), .C2 (n_70_46) );
AOI211_X1 g_51_54 (.ZN (n_51_54), .A (n_55_52), .B (n_61_49), .C1 (n_65_47), .C2 (n_68_47) );
AOI211_X1 g_49_55 (.ZN (n_49_55), .A (n_53_53), .B (n_59_50), .C1 (n_63_48), .C2 (n_66_48) );
AOI211_X1 g_47_56 (.ZN (n_47_56), .A (n_51_54), .B (n_57_51), .C1 (n_61_49), .C2 (n_64_49) );
AOI211_X1 g_45_57 (.ZN (n_45_57), .A (n_49_55), .B (n_55_52), .C1 (n_59_50), .C2 (n_65_47) );
AOI211_X1 g_46_55 (.ZN (n_46_55), .A (n_47_56), .B (n_53_53), .C1 (n_57_51), .C2 (n_63_48) );
AOI211_X1 g_44_56 (.ZN (n_44_56), .A (n_45_57), .B (n_51_54), .C1 (n_55_52), .C2 (n_61_49) );
AOI211_X1 g_42_57 (.ZN (n_42_57), .A (n_46_55), .B (n_49_55), .C1 (n_53_53), .C2 (n_59_50) );
AOI211_X1 g_40_58 (.ZN (n_40_58), .A (n_44_56), .B (n_47_56), .C1 (n_51_54), .C2 (n_57_51) );
AOI211_X1 g_38_59 (.ZN (n_38_59), .A (n_42_57), .B (n_45_57), .C1 (n_49_55), .C2 (n_55_52) );
AOI211_X1 g_36_60 (.ZN (n_36_60), .A (n_40_58), .B (n_46_55), .C1 (n_47_56), .C2 (n_53_53) );
AOI211_X1 g_34_61 (.ZN (n_34_61), .A (n_38_59), .B (n_44_56), .C1 (n_45_57), .C2 (n_51_54) );
AOI211_X1 g_32_62 (.ZN (n_32_62), .A (n_36_60), .B (n_42_57), .C1 (n_46_55), .C2 (n_49_55) );
AOI211_X1 g_30_63 (.ZN (n_30_63), .A (n_34_61), .B (n_40_58), .C1 (n_44_56), .C2 (n_47_56) );
AOI211_X1 g_28_64 (.ZN (n_28_64), .A (n_32_62), .B (n_38_59), .C1 (n_42_57), .C2 (n_45_57) );
AOI211_X1 g_26_65 (.ZN (n_26_65), .A (n_30_63), .B (n_36_60), .C1 (n_40_58), .C2 (n_46_55) );
AOI211_X1 g_24_66 (.ZN (n_24_66), .A (n_28_64), .B (n_34_61), .C1 (n_38_59), .C2 (n_44_56) );
AOI211_X1 g_22_67 (.ZN (n_22_67), .A (n_26_65), .B (n_32_62), .C1 (n_36_60), .C2 (n_42_57) );
AOI211_X1 g_20_68 (.ZN (n_20_68), .A (n_24_66), .B (n_30_63), .C1 (n_34_61), .C2 (n_40_58) );
AOI211_X1 g_18_69 (.ZN (n_18_69), .A (n_22_67), .B (n_28_64), .C1 (n_32_62), .C2 (n_38_59) );
AOI211_X1 g_16_70 (.ZN (n_16_70), .A (n_20_68), .B (n_26_65), .C1 (n_30_63), .C2 (n_36_60) );
AOI211_X1 g_14_71 (.ZN (n_14_71), .A (n_18_69), .B (n_24_66), .C1 (n_28_64), .C2 (n_34_61) );
AOI211_X1 g_12_72 (.ZN (n_12_72), .A (n_16_70), .B (n_22_67), .C1 (n_26_65), .C2 (n_32_62) );
AOI211_X1 g_10_73 (.ZN (n_10_73), .A (n_14_71), .B (n_20_68), .C1 (n_24_66), .C2 (n_30_63) );
AOI211_X1 g_11_71 (.ZN (n_11_71), .A (n_12_72), .B (n_18_69), .C1 (n_22_67), .C2 (n_28_64) );
AOI211_X1 g_13_72 (.ZN (n_13_72), .A (n_10_73), .B (n_16_70), .C1 (n_20_68), .C2 (n_26_65) );
AOI211_X1 g_14_70 (.ZN (n_14_70), .A (n_11_71), .B (n_14_71), .C1 (n_18_69), .C2 (n_24_66) );
AOI211_X1 g_16_69 (.ZN (n_16_69), .A (n_13_72), .B (n_12_72), .C1 (n_16_70), .C2 (n_22_67) );
AOI211_X1 g_18_68 (.ZN (n_18_68), .A (n_14_70), .B (n_10_73), .C1 (n_14_71), .C2 (n_20_68) );
AOI211_X1 g_20_67 (.ZN (n_20_67), .A (n_16_69), .B (n_11_71), .C1 (n_12_72), .C2 (n_18_69) );
AOI211_X1 g_22_66 (.ZN (n_22_66), .A (n_18_68), .B (n_13_72), .C1 (n_10_73), .C2 (n_16_70) );
AOI211_X1 g_24_65 (.ZN (n_24_65), .A (n_20_67), .B (n_14_70), .C1 (n_11_71), .C2 (n_14_71) );
AOI211_X1 g_26_64 (.ZN (n_26_64), .A (n_22_66), .B (n_16_69), .C1 (n_13_72), .C2 (n_12_72) );
AOI211_X1 g_28_63 (.ZN (n_28_63), .A (n_24_65), .B (n_18_68), .C1 (n_14_70), .C2 (n_10_73) );
AOI211_X1 g_30_62 (.ZN (n_30_62), .A (n_26_64), .B (n_20_67), .C1 (n_16_69), .C2 (n_11_71) );
AOI211_X1 g_32_61 (.ZN (n_32_61), .A (n_28_63), .B (n_22_66), .C1 (n_18_68), .C2 (n_13_72) );
AOI211_X1 g_31_63 (.ZN (n_31_63), .A (n_30_62), .B (n_24_65), .C1 (n_20_67), .C2 (n_14_70) );
AOI211_X1 g_33_62 (.ZN (n_33_62), .A (n_32_61), .B (n_26_64), .C1 (n_22_66), .C2 (n_16_69) );
AOI211_X1 g_35_61 (.ZN (n_35_61), .A (n_31_63), .B (n_28_63), .C1 (n_24_65), .C2 (n_18_68) );
AOI211_X1 g_37_60 (.ZN (n_37_60), .A (n_33_62), .B (n_30_62), .C1 (n_26_64), .C2 (n_20_67) );
AOI211_X1 g_39_59 (.ZN (n_39_59), .A (n_35_61), .B (n_32_61), .C1 (n_28_63), .C2 (n_22_66) );
AOI211_X1 g_41_58 (.ZN (n_41_58), .A (n_37_60), .B (n_31_63), .C1 (n_30_62), .C2 (n_24_65) );
AOI211_X1 g_43_57 (.ZN (n_43_57), .A (n_39_59), .B (n_33_62), .C1 (n_32_61), .C2 (n_26_64) );
AOI211_X1 g_45_56 (.ZN (n_45_56), .A (n_41_58), .B (n_35_61), .C1 (n_31_63), .C2 (n_28_63) );
AOI211_X1 g_47_55 (.ZN (n_47_55), .A (n_43_57), .B (n_37_60), .C1 (n_33_62), .C2 (n_30_62) );
AOI211_X1 g_46_57 (.ZN (n_46_57), .A (n_45_56), .B (n_39_59), .C1 (n_35_61), .C2 (n_32_61) );
AOI211_X1 g_48_56 (.ZN (n_48_56), .A (n_47_55), .B (n_41_58), .C1 (n_37_60), .C2 (n_31_63) );
AOI211_X1 g_47_58 (.ZN (n_47_58), .A (n_46_57), .B (n_43_57), .C1 (n_39_59), .C2 (n_33_62) );
AOI211_X1 g_46_56 (.ZN (n_46_56), .A (n_48_56), .B (n_45_56), .C1 (n_41_58), .C2 (n_35_61) );
AOI211_X1 g_48_55 (.ZN (n_48_55), .A (n_47_58), .B (n_47_55), .C1 (n_43_57), .C2 (n_37_60) );
AOI211_X1 g_49_57 (.ZN (n_49_57), .A (n_46_56), .B (n_46_57), .C1 (n_45_56), .C2 (n_39_59) );
AOI211_X1 g_51_56 (.ZN (n_51_56), .A (n_48_55), .B (n_48_56), .C1 (n_47_55), .C2 (n_41_58) );
AOI211_X1 g_53_55 (.ZN (n_53_55), .A (n_49_57), .B (n_47_58), .C1 (n_46_57), .C2 (n_43_57) );
AOI211_X1 g_55_54 (.ZN (n_55_54), .A (n_51_56), .B (n_46_56), .C1 (n_48_56), .C2 (n_45_56) );
AOI211_X1 g_57_53 (.ZN (n_57_53), .A (n_53_55), .B (n_48_55), .C1 (n_47_58), .C2 (n_47_55) );
AOI211_X1 g_59_52 (.ZN (n_59_52), .A (n_55_54), .B (n_49_57), .C1 (n_46_56), .C2 (n_46_57) );
AOI211_X1 g_61_51 (.ZN (n_61_51), .A (n_57_53), .B (n_51_56), .C1 (n_48_55), .C2 (n_48_56) );
AOI211_X1 g_63_50 (.ZN (n_63_50), .A (n_59_52), .B (n_53_55), .C1 (n_49_57), .C2 (n_47_58) );
AOI211_X1 g_65_49 (.ZN (n_65_49), .A (n_61_51), .B (n_55_54), .C1 (n_51_56), .C2 (n_46_56) );
AOI211_X1 g_67_48 (.ZN (n_67_48), .A (n_63_50), .B (n_57_53), .C1 (n_53_55), .C2 (n_48_55) );
AOI211_X1 g_69_47 (.ZN (n_69_47), .A (n_65_49), .B (n_59_52), .C1 (n_55_54), .C2 (n_49_57) );
AOI211_X1 g_71_46 (.ZN (n_71_46), .A (n_67_48), .B (n_61_51), .C1 (n_57_53), .C2 (n_51_56) );
AOI211_X1 g_70_48 (.ZN (n_70_48), .A (n_69_47), .B (n_63_50), .C1 (n_59_52), .C2 (n_53_55) );
AOI211_X1 g_69_46 (.ZN (n_69_46), .A (n_71_46), .B (n_65_49), .C1 (n_61_51), .C2 (n_55_54) );
AOI211_X1 g_71_45 (.ZN (n_71_45), .A (n_70_48), .B (n_67_48), .C1 (n_63_50), .C2 (n_57_53) );
AOI211_X1 g_73_44 (.ZN (n_73_44), .A (n_69_46), .B (n_69_47), .C1 (n_65_49), .C2 (n_59_52) );
AOI211_X1 g_75_43 (.ZN (n_75_43), .A (n_71_45), .B (n_71_46), .C1 (n_67_48), .C2 (n_61_51) );
AOI211_X1 g_76_45 (.ZN (n_76_45), .A (n_73_44), .B (n_70_48), .C1 (n_69_47), .C2 (n_63_50) );
AOI211_X1 g_74_46 (.ZN (n_74_46), .A (n_75_43), .B (n_69_46), .C1 (n_71_46), .C2 (n_65_49) );
AOI211_X1 g_72_47 (.ZN (n_72_47), .A (n_76_45), .B (n_71_45), .C1 (n_70_48), .C2 (n_67_48) );
AOI211_X1 g_71_49 (.ZN (n_71_49), .A (n_74_46), .B (n_73_44), .C1 (n_69_46), .C2 (n_69_47) );
AOI211_X1 g_70_47 (.ZN (n_70_47), .A (n_72_47), .B (n_75_43), .C1 (n_71_45), .C2 (n_71_46) );
AOI211_X1 g_72_46 (.ZN (n_72_46), .A (n_71_49), .B (n_76_45), .C1 (n_73_44), .C2 (n_70_48) );
AOI211_X1 g_74_45 (.ZN (n_74_45), .A (n_70_47), .B (n_74_46), .C1 (n_75_43), .C2 (n_69_46) );
AOI211_X1 g_76_44 (.ZN (n_76_44), .A (n_72_46), .B (n_72_47), .C1 (n_76_45), .C2 (n_71_45) );
AOI211_X1 g_78_43 (.ZN (n_78_43), .A (n_74_45), .B (n_71_49), .C1 (n_74_46), .C2 (n_73_44) );
AOI211_X1 g_80_42 (.ZN (n_80_42), .A (n_76_44), .B (n_70_47), .C1 (n_72_47), .C2 (n_75_43) );
AOI211_X1 g_82_41 (.ZN (n_82_41), .A (n_78_43), .B (n_72_46), .C1 (n_71_49), .C2 (n_76_45) );
AOI211_X1 g_84_40 (.ZN (n_84_40), .A (n_80_42), .B (n_74_45), .C1 (n_70_47), .C2 (n_74_46) );
AOI211_X1 g_86_39 (.ZN (n_86_39), .A (n_82_41), .B (n_76_44), .C1 (n_72_46), .C2 (n_72_47) );
AOI211_X1 g_88_38 (.ZN (n_88_38), .A (n_84_40), .B (n_78_43), .C1 (n_74_45), .C2 (n_71_49) );
AOI211_X1 g_90_37 (.ZN (n_90_37), .A (n_86_39), .B (n_80_42), .C1 (n_76_44), .C2 (n_70_47) );
AOI211_X1 g_89_39 (.ZN (n_89_39), .A (n_88_38), .B (n_82_41), .C1 (n_78_43), .C2 (n_72_46) );
AOI211_X1 g_91_38 (.ZN (n_91_38), .A (n_90_37), .B (n_84_40), .C1 (n_80_42), .C2 (n_74_45) );
AOI211_X1 g_93_37 (.ZN (n_93_37), .A (n_89_39), .B (n_86_39), .C1 (n_82_41), .C2 (n_76_44) );
AOI211_X1 g_92_39 (.ZN (n_92_39), .A (n_91_38), .B (n_88_38), .C1 (n_84_40), .C2 (n_78_43) );
AOI211_X1 g_91_37 (.ZN (n_91_37), .A (n_93_37), .B (n_90_37), .C1 (n_86_39), .C2 (n_80_42) );
AOI211_X1 g_93_36 (.ZN (n_93_36), .A (n_92_39), .B (n_89_39), .C1 (n_88_38), .C2 (n_82_41) );
AOI211_X1 g_95_35 (.ZN (n_95_35), .A (n_91_37), .B (n_91_38), .C1 (n_90_37), .C2 (n_84_40) );
AOI211_X1 g_97_34 (.ZN (n_97_34), .A (n_93_36), .B (n_93_37), .C1 (n_89_39), .C2 (n_86_39) );
AOI211_X1 g_99_35 (.ZN (n_99_35), .A (n_95_35), .B (n_92_39), .C1 (n_91_38), .C2 (n_88_38) );
AOI211_X1 g_100_37 (.ZN (n_100_37), .A (n_97_34), .B (n_91_37), .C1 (n_93_37), .C2 (n_90_37) );
AOI211_X1 g_98_36 (.ZN (n_98_36), .A (n_99_35), .B (n_93_36), .C1 (n_92_39), .C2 (n_89_39) );
AOI211_X1 g_96_35 (.ZN (n_96_35), .A (n_100_37), .B (n_95_35), .C1 (n_91_37), .C2 (n_91_38) );
AOI211_X1 g_94_36 (.ZN (n_94_36), .A (n_98_36), .B (n_97_34), .C1 (n_93_36), .C2 (n_93_37) );
AOI211_X1 g_92_37 (.ZN (n_92_37), .A (n_96_35), .B (n_99_35), .C1 (n_95_35), .C2 (n_92_39) );
AOI211_X1 g_90_38 (.ZN (n_90_38), .A (n_94_36), .B (n_100_37), .C1 (n_97_34), .C2 (n_91_37) );
AOI211_X1 g_88_39 (.ZN (n_88_39), .A (n_92_37), .B (n_98_36), .C1 (n_99_35), .C2 (n_93_36) );
AOI211_X1 g_86_40 (.ZN (n_86_40), .A (n_90_38), .B (n_96_35), .C1 (n_100_37), .C2 (n_95_35) );
AOI211_X1 g_84_41 (.ZN (n_84_41), .A (n_88_39), .B (n_94_36), .C1 (n_98_36), .C2 (n_97_34) );
AOI211_X1 g_82_42 (.ZN (n_82_42), .A (n_86_40), .B (n_92_37), .C1 (n_96_35), .C2 (n_99_35) );
AOI211_X1 g_80_43 (.ZN (n_80_43), .A (n_84_41), .B (n_90_38), .C1 (n_94_36), .C2 (n_100_37) );
AOI211_X1 g_79_45 (.ZN (n_79_45), .A (n_82_42), .B (n_88_39), .C1 (n_92_37), .C2 (n_98_36) );
AOI211_X1 g_77_44 (.ZN (n_77_44), .A (n_80_43), .B (n_86_40), .C1 (n_90_38), .C2 (n_96_35) );
AOI211_X1 g_79_43 (.ZN (n_79_43), .A (n_79_45), .B (n_84_41), .C1 (n_88_39), .C2 (n_94_36) );
AOI211_X1 g_81_42 (.ZN (n_81_42), .A (n_77_44), .B (n_82_42), .C1 (n_86_40), .C2 (n_92_37) );
AOI211_X1 g_83_41 (.ZN (n_83_41), .A (n_79_43), .B (n_80_43), .C1 (n_84_41), .C2 (n_90_38) );
AOI211_X1 g_85_40 (.ZN (n_85_40), .A (n_81_42), .B (n_79_45), .C1 (n_82_42), .C2 (n_88_39) );
AOI211_X1 g_87_39 (.ZN (n_87_39), .A (n_83_41), .B (n_77_44), .C1 (n_80_43), .C2 (n_86_40) );
AOI211_X1 g_89_38 (.ZN (n_89_38), .A (n_85_40), .B (n_79_43), .C1 (n_79_45), .C2 (n_84_41) );
AOI211_X1 g_90_40 (.ZN (n_90_40), .A (n_87_39), .B (n_81_42), .C1 (n_77_44), .C2 (n_82_42) );
AOI211_X1 g_88_41 (.ZN (n_88_41), .A (n_89_38), .B (n_83_41), .C1 (n_79_43), .C2 (n_80_43) );
AOI211_X1 g_86_42 (.ZN (n_86_42), .A (n_90_40), .B (n_85_40), .C1 (n_81_42), .C2 (n_79_45) );
AOI211_X1 g_87_40 (.ZN (n_87_40), .A (n_88_41), .B (n_87_39), .C1 (n_83_41), .C2 (n_77_44) );
AOI211_X1 g_85_41 (.ZN (n_85_41), .A (n_86_42), .B (n_89_38), .C1 (n_85_40), .C2 (n_79_43) );
AOI211_X1 g_83_42 (.ZN (n_83_42), .A (n_87_40), .B (n_90_40), .C1 (n_87_39), .C2 (n_81_42) );
AOI211_X1 g_81_43 (.ZN (n_81_43), .A (n_85_41), .B (n_88_41), .C1 (n_89_38), .C2 (n_83_41) );
AOI211_X1 g_79_44 (.ZN (n_79_44), .A (n_83_42), .B (n_86_42), .C1 (n_90_40), .C2 (n_85_40) );
AOI211_X1 g_77_45 (.ZN (n_77_45), .A (n_81_43), .B (n_87_40), .C1 (n_88_41), .C2 (n_87_39) );
AOI211_X1 g_75_46 (.ZN (n_75_46), .A (n_79_44), .B (n_85_41), .C1 (n_86_42), .C2 (n_89_38) );
AOI211_X1 g_73_47 (.ZN (n_73_47), .A (n_77_45), .B (n_83_42), .C1 (n_87_40), .C2 (n_90_40) );
AOI211_X1 g_71_48 (.ZN (n_71_48), .A (n_75_46), .B (n_81_43), .C1 (n_85_41), .C2 (n_88_41) );
AOI211_X1 g_69_49 (.ZN (n_69_49), .A (n_73_47), .B (n_79_44), .C1 (n_83_42), .C2 (n_86_42) );
AOI211_X1 g_67_50 (.ZN (n_67_50), .A (n_71_48), .B (n_77_45), .C1 (n_81_43), .C2 (n_87_40) );
AOI211_X1 g_68_48 (.ZN (n_68_48), .A (n_69_49), .B (n_75_46), .C1 (n_79_44), .C2 (n_85_41) );
AOI211_X1 g_66_49 (.ZN (n_66_49), .A (n_67_50), .B (n_73_47), .C1 (n_77_45), .C2 (n_83_42) );
AOI211_X1 g_67_47 (.ZN (n_67_47), .A (n_68_48), .B (n_71_48), .C1 (n_75_46), .C2 (n_81_43) );
AOI211_X1 g_65_48 (.ZN (n_65_48), .A (n_66_49), .B (n_69_49), .C1 (n_73_47), .C2 (n_79_44) );
AOI211_X1 g_63_49 (.ZN (n_63_49), .A (n_67_47), .B (n_67_50), .C1 (n_71_48), .C2 (n_77_45) );
AOI211_X1 g_61_50 (.ZN (n_61_50), .A (n_65_48), .B (n_68_48), .C1 (n_69_49), .C2 (n_75_46) );
AOI211_X1 g_59_51 (.ZN (n_59_51), .A (n_63_49), .B (n_66_49), .C1 (n_67_50), .C2 (n_73_47) );
AOI211_X1 g_57_52 (.ZN (n_57_52), .A (n_61_50), .B (n_67_47), .C1 (n_68_48), .C2 (n_71_48) );
AOI211_X1 g_55_53 (.ZN (n_55_53), .A (n_59_51), .B (n_65_48), .C1 (n_66_49), .C2 (n_69_49) );
AOI211_X1 g_53_54 (.ZN (n_53_54), .A (n_57_52), .B (n_63_49), .C1 (n_67_47), .C2 (n_67_50) );
AOI211_X1 g_51_55 (.ZN (n_51_55), .A (n_55_53), .B (n_61_50), .C1 (n_65_48), .C2 (n_68_48) );
AOI211_X1 g_49_56 (.ZN (n_49_56), .A (n_53_54), .B (n_59_51), .C1 (n_63_49), .C2 (n_66_49) );
AOI211_X1 g_47_57 (.ZN (n_47_57), .A (n_51_55), .B (n_57_52), .C1 (n_61_50), .C2 (n_67_47) );
AOI211_X1 g_45_58 (.ZN (n_45_58), .A (n_49_56), .B (n_55_53), .C1 (n_59_51), .C2 (n_65_48) );
AOI211_X1 g_43_59 (.ZN (n_43_59), .A (n_47_57), .B (n_53_54), .C1 (n_57_52), .C2 (n_63_49) );
AOI211_X1 g_44_57 (.ZN (n_44_57), .A (n_45_58), .B (n_51_55), .C1 (n_55_53), .C2 (n_61_50) );
AOI211_X1 g_42_58 (.ZN (n_42_58), .A (n_43_59), .B (n_49_56), .C1 (n_53_54), .C2 (n_59_51) );
AOI211_X1 g_40_59 (.ZN (n_40_59), .A (n_44_57), .B (n_47_57), .C1 (n_51_55), .C2 (n_57_52) );
AOI211_X1 g_38_60 (.ZN (n_38_60), .A (n_42_58), .B (n_45_58), .C1 (n_49_56), .C2 (n_55_53) );
AOI211_X1 g_36_61 (.ZN (n_36_61), .A (n_40_59), .B (n_43_59), .C1 (n_47_57), .C2 (n_53_54) );
AOI211_X1 g_34_62 (.ZN (n_34_62), .A (n_38_60), .B (n_44_57), .C1 (n_45_58), .C2 (n_51_55) );
AOI211_X1 g_32_63 (.ZN (n_32_63), .A (n_36_61), .B (n_42_58), .C1 (n_43_59), .C2 (n_49_56) );
AOI211_X1 g_30_64 (.ZN (n_30_64), .A (n_34_62), .B (n_40_59), .C1 (n_44_57), .C2 (n_47_57) );
AOI211_X1 g_28_65 (.ZN (n_28_65), .A (n_32_63), .B (n_38_60), .C1 (n_42_58), .C2 (n_45_58) );
AOI211_X1 g_26_66 (.ZN (n_26_66), .A (n_30_64), .B (n_36_61), .C1 (n_40_59), .C2 (n_43_59) );
AOI211_X1 g_24_67 (.ZN (n_24_67), .A (n_28_65), .B (n_34_62), .C1 (n_38_60), .C2 (n_44_57) );
AOI211_X1 g_25_65 (.ZN (n_25_65), .A (n_26_66), .B (n_32_63), .C1 (n_36_61), .C2 (n_42_58) );
AOI211_X1 g_23_66 (.ZN (n_23_66), .A (n_24_67), .B (n_30_64), .C1 (n_34_62), .C2 (n_40_59) );
AOI211_X1 g_21_67 (.ZN (n_21_67), .A (n_25_65), .B (n_28_65), .C1 (n_32_63), .C2 (n_38_60) );
AOI211_X1 g_19_68 (.ZN (n_19_68), .A (n_23_66), .B (n_26_66), .C1 (n_30_64), .C2 (n_36_61) );
AOI211_X1 g_18_70 (.ZN (n_18_70), .A (n_21_67), .B (n_24_67), .C1 (n_28_65), .C2 (n_34_62) );
AOI211_X1 g_20_69 (.ZN (n_20_69), .A (n_19_68), .B (n_25_65), .C1 (n_26_66), .C2 (n_32_63) );
AOI211_X1 g_22_68 (.ZN (n_22_68), .A (n_18_70), .B (n_23_66), .C1 (n_24_67), .C2 (n_30_64) );
AOI211_X1 g_21_70 (.ZN (n_21_70), .A (n_20_69), .B (n_21_67), .C1 (n_25_65), .C2 (n_28_65) );
AOI211_X1 g_19_69 (.ZN (n_19_69), .A (n_22_68), .B (n_19_68), .C1 (n_23_66), .C2 (n_26_66) );
AOI211_X1 g_21_68 (.ZN (n_21_68), .A (n_21_70), .B (n_18_70), .C1 (n_21_67), .C2 (n_24_67) );
AOI211_X1 g_23_67 (.ZN (n_23_67), .A (n_19_69), .B (n_20_69), .C1 (n_19_68), .C2 (n_25_65) );
AOI211_X1 g_25_66 (.ZN (n_25_66), .A (n_21_68), .B (n_22_68), .C1 (n_18_70), .C2 (n_23_66) );
AOI211_X1 g_27_65 (.ZN (n_27_65), .A (n_23_67), .B (n_21_70), .C1 (n_20_69), .C2 (n_21_67) );
AOI211_X1 g_29_64 (.ZN (n_29_64), .A (n_25_66), .B (n_19_69), .C1 (n_22_68), .C2 (n_19_68) );
AOI211_X1 g_28_66 (.ZN (n_28_66), .A (n_27_65), .B (n_21_68), .C1 (n_21_70), .C2 (n_18_70) );
AOI211_X1 g_30_65 (.ZN (n_30_65), .A (n_29_64), .B (n_23_67), .C1 (n_19_69), .C2 (n_20_69) );
AOI211_X1 g_32_64 (.ZN (n_32_64), .A (n_28_66), .B (n_25_66), .C1 (n_21_68), .C2 (n_22_68) );
AOI211_X1 g_34_63 (.ZN (n_34_63), .A (n_30_65), .B (n_27_65), .C1 (n_23_67), .C2 (n_21_70) );
AOI211_X1 g_36_62 (.ZN (n_36_62), .A (n_32_64), .B (n_29_64), .C1 (n_25_66), .C2 (n_19_69) );
AOI211_X1 g_38_61 (.ZN (n_38_61), .A (n_34_63), .B (n_28_66), .C1 (n_27_65), .C2 (n_21_68) );
AOI211_X1 g_40_60 (.ZN (n_40_60), .A (n_36_62), .B (n_30_65), .C1 (n_29_64), .C2 (n_23_67) );
AOI211_X1 g_42_59 (.ZN (n_42_59), .A (n_38_61), .B (n_32_64), .C1 (n_28_66), .C2 (n_25_66) );
AOI211_X1 g_44_58 (.ZN (n_44_58), .A (n_40_60), .B (n_34_63), .C1 (n_30_65), .C2 (n_27_65) );
AOI211_X1 g_46_59 (.ZN (n_46_59), .A (n_42_59), .B (n_36_62), .C1 (n_32_64), .C2 (n_29_64) );
AOI211_X1 g_48_58 (.ZN (n_48_58), .A (n_44_58), .B (n_38_61), .C1 (n_34_63), .C2 (n_28_66) );
AOI211_X1 g_50_57 (.ZN (n_50_57), .A (n_46_59), .B (n_40_60), .C1 (n_36_62), .C2 (n_30_65) );
AOI211_X1 g_52_56 (.ZN (n_52_56), .A (n_48_58), .B (n_42_59), .C1 (n_38_61), .C2 (n_32_64) );
AOI211_X1 g_54_55 (.ZN (n_54_55), .A (n_50_57), .B (n_44_58), .C1 (n_40_60), .C2 (n_34_63) );
AOI211_X1 g_56_54 (.ZN (n_56_54), .A (n_52_56), .B (n_46_59), .C1 (n_42_59), .C2 (n_36_62) );
AOI211_X1 g_58_53 (.ZN (n_58_53), .A (n_54_55), .B (n_48_58), .C1 (n_44_58), .C2 (n_38_61) );
AOI211_X1 g_60_52 (.ZN (n_60_52), .A (n_56_54), .B (n_50_57), .C1 (n_46_59), .C2 (n_40_60) );
AOI211_X1 g_62_51 (.ZN (n_62_51), .A (n_58_53), .B (n_52_56), .C1 (n_48_58), .C2 (n_42_59) );
AOI211_X1 g_64_50 (.ZN (n_64_50), .A (n_60_52), .B (n_54_55), .C1 (n_50_57), .C2 (n_44_58) );
AOI211_X1 g_63_52 (.ZN (n_63_52), .A (n_62_51), .B (n_56_54), .C1 (n_52_56), .C2 (n_46_59) );
AOI211_X1 g_65_51 (.ZN (n_65_51), .A (n_64_50), .B (n_58_53), .C1 (n_54_55), .C2 (n_48_58) );
AOI211_X1 g_64_53 (.ZN (n_64_53), .A (n_63_52), .B (n_60_52), .C1 (n_56_54), .C2 (n_50_57) );
AOI211_X1 g_63_51 (.ZN (n_63_51), .A (n_65_51), .B (n_62_51), .C1 (n_58_53), .C2 (n_52_56) );
AOI211_X1 g_65_50 (.ZN (n_65_50), .A (n_64_53), .B (n_64_50), .C1 (n_60_52), .C2 (n_54_55) );
AOI211_X1 g_67_49 (.ZN (n_67_49), .A (n_63_51), .B (n_63_52), .C1 (n_62_51), .C2 (n_56_54) );
AOI211_X1 g_69_48 (.ZN (n_69_48), .A (n_65_50), .B (n_65_51), .C1 (n_64_50), .C2 (n_58_53) );
AOI211_X1 g_71_47 (.ZN (n_71_47), .A (n_67_49), .B (n_64_53), .C1 (n_63_52), .C2 (n_60_52) );
AOI211_X1 g_73_46 (.ZN (n_73_46), .A (n_69_48), .B (n_63_51), .C1 (n_65_51), .C2 (n_62_51) );
AOI211_X1 g_75_45 (.ZN (n_75_45), .A (n_71_47), .B (n_65_50), .C1 (n_64_53), .C2 (n_64_50) );
AOI211_X1 g_77_46 (.ZN (n_77_46), .A (n_73_46), .B (n_67_49), .C1 (n_63_51), .C2 (n_63_52) );
AOI211_X1 g_75_47 (.ZN (n_75_47), .A (n_75_45), .B (n_69_48), .C1 (n_65_50), .C2 (n_65_51) );
AOI211_X1 g_73_48 (.ZN (n_73_48), .A (n_77_46), .B (n_71_47), .C1 (n_67_49), .C2 (n_64_53) );
AOI211_X1 g_72_50 (.ZN (n_72_50), .A (n_75_47), .B (n_73_46), .C1 (n_69_48), .C2 (n_63_51) );
AOI211_X1 g_70_49 (.ZN (n_70_49), .A (n_73_48), .B (n_75_45), .C1 (n_71_47), .C2 (n_65_50) );
AOI211_X1 g_72_48 (.ZN (n_72_48), .A (n_72_50), .B (n_77_46), .C1 (n_73_46), .C2 (n_67_49) );
AOI211_X1 g_74_47 (.ZN (n_74_47), .A (n_70_49), .B (n_75_47), .C1 (n_75_45), .C2 (n_69_48) );
AOI211_X1 g_76_46 (.ZN (n_76_46), .A (n_72_48), .B (n_73_48), .C1 (n_77_46), .C2 (n_71_47) );
AOI211_X1 g_78_45 (.ZN (n_78_45), .A (n_74_47), .B (n_72_50), .C1 (n_75_47), .C2 (n_73_46) );
AOI211_X1 g_80_44 (.ZN (n_80_44), .A (n_76_46), .B (n_70_49), .C1 (n_73_48), .C2 (n_75_45) );
AOI211_X1 g_82_43 (.ZN (n_82_43), .A (n_78_45), .B (n_72_48), .C1 (n_72_50), .C2 (n_77_46) );
AOI211_X1 g_84_42 (.ZN (n_84_42), .A (n_80_44), .B (n_74_47), .C1 (n_70_49), .C2 (n_75_47) );
AOI211_X1 g_86_41 (.ZN (n_86_41), .A (n_82_43), .B (n_76_46), .C1 (n_72_48), .C2 (n_73_48) );
AOI211_X1 g_88_40 (.ZN (n_88_40), .A (n_84_42), .B (n_78_45), .C1 (n_74_47), .C2 (n_72_50) );
AOI211_X1 g_90_39 (.ZN (n_90_39), .A (n_86_41), .B (n_80_44), .C1 (n_76_46), .C2 (n_70_49) );
AOI211_X1 g_92_38 (.ZN (n_92_38), .A (n_88_40), .B (n_82_43), .C1 (n_78_45), .C2 (n_72_48) );
AOI211_X1 g_94_37 (.ZN (n_94_37), .A (n_90_39), .B (n_84_42), .C1 (n_80_44), .C2 (n_74_47) );
AOI211_X1 g_96_36 (.ZN (n_96_36), .A (n_92_38), .B (n_86_41), .C1 (n_82_43), .C2 (n_76_46) );
AOI211_X1 g_98_35 (.ZN (n_98_35), .A (n_94_37), .B (n_88_40), .C1 (n_84_42), .C2 (n_78_45) );
AOI211_X1 g_100_36 (.ZN (n_100_36), .A (n_96_36), .B (n_90_39), .C1 (n_86_41), .C2 (n_80_44) );
AOI211_X1 g_98_37 (.ZN (n_98_37), .A (n_98_35), .B (n_92_38), .C1 (n_88_40), .C2 (n_82_43) );
AOI211_X1 g_99_39 (.ZN (n_99_39), .A (n_100_36), .B (n_94_37), .C1 (n_90_39), .C2 (n_84_42) );
AOI211_X1 g_100_41 (.ZN (n_100_41), .A (n_98_37), .B (n_96_36), .C1 (n_92_38), .C2 (n_86_41) );
AOI211_X1 g_98_42 (.ZN (n_98_42), .A (n_99_39), .B (n_98_35), .C1 (n_94_37), .C2 (n_88_40) );
AOI211_X1 g_100_43 (.ZN (n_100_43), .A (n_100_41), .B (n_100_36), .C1 (n_96_36), .C2 (n_90_39) );
AOI211_X1 g_99_41 (.ZN (n_99_41), .A (n_98_42), .B (n_98_37), .C1 (n_98_35), .C2 (n_92_38) );
AOI211_X1 g_100_39 (.ZN (n_100_39), .A (n_100_43), .B (n_99_39), .C1 (n_100_36), .C2 (n_94_37) );
AOI211_X1 g_99_37 (.ZN (n_99_37), .A (n_99_41), .B (n_100_41), .C1 (n_98_37), .C2 (n_96_36) );
AOI211_X1 g_97_36 (.ZN (n_97_36), .A (n_100_39), .B (n_98_42), .C1 (n_99_39), .C2 (n_98_35) );
AOI211_X1 g_98_38 (.ZN (n_98_38), .A (n_99_37), .B (n_100_43), .C1 (n_100_41), .C2 (n_100_36) );
AOI211_X1 g_96_37 (.ZN (n_96_37), .A (n_97_36), .B (n_99_41), .C1 (n_98_42), .C2 (n_98_37) );
AOI211_X1 g_94_38 (.ZN (n_94_38), .A (n_98_38), .B (n_100_39), .C1 (n_100_43), .C2 (n_99_39) );
AOI211_X1 g_93_40 (.ZN (n_93_40), .A (n_96_37), .B (n_99_37), .C1 (n_99_41), .C2 (n_100_41) );
AOI211_X1 g_91_39 (.ZN (n_91_39), .A (n_94_38), .B (n_97_36), .C1 (n_100_39), .C2 (n_98_42) );
AOI211_X1 g_93_38 (.ZN (n_93_38), .A (n_93_40), .B (n_98_38), .C1 (n_99_37), .C2 (n_100_43) );
AOI211_X1 g_95_37 (.ZN (n_95_37), .A (n_91_39), .B (n_96_37), .C1 (n_97_36), .C2 (n_99_41) );
AOI211_X1 g_97_38 (.ZN (n_97_38), .A (n_93_38), .B (n_94_38), .C1 (n_98_38), .C2 (n_100_39) );
AOI211_X1 g_95_39 (.ZN (n_95_39), .A (n_95_37), .B (n_93_40), .C1 (n_96_37), .C2 (n_99_37) );
AOI211_X1 g_97_40 (.ZN (n_97_40), .A (n_97_38), .B (n_91_39), .C1 (n_94_38), .C2 (n_97_36) );
AOI211_X1 g_96_38 (.ZN (n_96_38), .A (n_95_39), .B (n_93_38), .C1 (n_93_40), .C2 (n_98_38) );
AOI211_X1 g_94_39 (.ZN (n_94_39), .A (n_97_40), .B (n_95_37), .C1 (n_91_39), .C2 (n_96_37) );
AOI211_X1 g_92_40 (.ZN (n_92_40), .A (n_96_38), .B (n_97_38), .C1 (n_93_38), .C2 (n_94_38) );
AOI211_X1 g_90_41 (.ZN (n_90_41), .A (n_94_39), .B (n_95_39), .C1 (n_95_37), .C2 (n_93_40) );
AOI211_X1 g_88_42 (.ZN (n_88_42), .A (n_92_40), .B (n_97_40), .C1 (n_97_38), .C2 (n_91_39) );
AOI211_X1 g_89_40 (.ZN (n_89_40), .A (n_90_41), .B (n_96_38), .C1 (n_95_39), .C2 (n_93_38) );
AOI211_X1 g_87_41 (.ZN (n_87_41), .A (n_88_42), .B (n_94_39), .C1 (n_97_40), .C2 (n_95_37) );
AOI211_X1 g_85_42 (.ZN (n_85_42), .A (n_89_40), .B (n_92_40), .C1 (n_96_38), .C2 (n_97_38) );
AOI211_X1 g_83_43 (.ZN (n_83_43), .A (n_87_41), .B (n_90_41), .C1 (n_94_39), .C2 (n_95_39) );
AOI211_X1 g_81_44 (.ZN (n_81_44), .A (n_85_42), .B (n_88_42), .C1 (n_92_40), .C2 (n_97_40) );
AOI211_X1 g_80_46 (.ZN (n_80_46), .A (n_83_43), .B (n_89_40), .C1 (n_90_41), .C2 (n_96_38) );
AOI211_X1 g_82_45 (.ZN (n_82_45), .A (n_81_44), .B (n_87_41), .C1 (n_88_42), .C2 (n_94_39) );
AOI211_X1 g_84_44 (.ZN (n_84_44), .A (n_80_46), .B (n_85_42), .C1 (n_89_40), .C2 (n_92_40) );
AOI211_X1 g_86_43 (.ZN (n_86_43), .A (n_82_45), .B (n_83_43), .C1 (n_87_41), .C2 (n_90_41) );
AOI211_X1 g_85_45 (.ZN (n_85_45), .A (n_84_44), .B (n_81_44), .C1 (n_85_42), .C2 (n_88_42) );
AOI211_X1 g_84_43 (.ZN (n_84_43), .A (n_86_43), .B (n_80_46), .C1 (n_83_43), .C2 (n_89_40) );
AOI211_X1 g_82_44 (.ZN (n_82_44), .A (n_85_45), .B (n_82_45), .C1 (n_81_44), .C2 (n_87_41) );
AOI211_X1 g_80_45 (.ZN (n_80_45), .A (n_84_43), .B (n_84_44), .C1 (n_80_46), .C2 (n_85_42) );
AOI211_X1 g_78_46 (.ZN (n_78_46), .A (n_82_44), .B (n_86_43), .C1 (n_82_45), .C2 (n_83_43) );
AOI211_X1 g_76_47 (.ZN (n_76_47), .A (n_80_45), .B (n_85_45), .C1 (n_84_44), .C2 (n_81_44) );
AOI211_X1 g_74_48 (.ZN (n_74_48), .A (n_78_46), .B (n_84_43), .C1 (n_86_43), .C2 (n_80_46) );
AOI211_X1 g_72_49 (.ZN (n_72_49), .A (n_76_47), .B (n_82_44), .C1 (n_85_45), .C2 (n_82_45) );
AOI211_X1 g_70_50 (.ZN (n_70_50), .A (n_74_48), .B (n_80_45), .C1 (n_84_43), .C2 (n_84_44) );
AOI211_X1 g_68_49 (.ZN (n_68_49), .A (n_72_49), .B (n_78_46), .C1 (n_82_44), .C2 (n_86_43) );
AOI211_X1 g_66_50 (.ZN (n_66_50), .A (n_70_50), .B (n_76_47), .C1 (n_80_45), .C2 (n_85_45) );
AOI211_X1 g_68_51 (.ZN (n_68_51), .A (n_68_49), .B (n_74_48), .C1 (n_78_46), .C2 (n_84_43) );
AOI211_X1 g_66_52 (.ZN (n_66_52), .A (n_66_50), .B (n_72_49), .C1 (n_76_47), .C2 (n_82_44) );
AOI211_X1 g_64_51 (.ZN (n_64_51), .A (n_68_51), .B (n_70_50), .C1 (n_74_48), .C2 (n_80_45) );
AOI211_X1 g_62_50 (.ZN (n_62_50), .A (n_66_52), .B (n_68_49), .C1 (n_72_49), .C2 (n_78_46) );
AOI211_X1 g_60_51 (.ZN (n_60_51), .A (n_64_51), .B (n_66_50), .C1 (n_70_50), .C2 (n_76_47) );
AOI211_X1 g_62_52 (.ZN (n_62_52), .A (n_62_50), .B (n_68_51), .C1 (n_68_49), .C2 (n_74_48) );
AOI211_X1 g_60_53 (.ZN (n_60_53), .A (n_60_51), .B (n_66_52), .C1 (n_66_50), .C2 (n_72_49) );
AOI211_X1 g_58_52 (.ZN (n_58_52), .A (n_62_52), .B (n_64_51), .C1 (n_68_51), .C2 (n_70_50) );
AOI211_X1 g_56_53 (.ZN (n_56_53), .A (n_60_53), .B (n_62_50), .C1 (n_66_52), .C2 (n_68_49) );
AOI211_X1 g_54_54 (.ZN (n_54_54), .A (n_58_52), .B (n_60_51), .C1 (n_64_51), .C2 (n_66_50) );
AOI211_X1 g_52_55 (.ZN (n_52_55), .A (n_56_53), .B (n_62_52), .C1 (n_62_50), .C2 (n_68_51) );
AOI211_X1 g_50_56 (.ZN (n_50_56), .A (n_54_54), .B (n_60_53), .C1 (n_60_51), .C2 (n_66_52) );
AOI211_X1 g_48_57 (.ZN (n_48_57), .A (n_52_55), .B (n_58_52), .C1 (n_62_52), .C2 (n_64_51) );
AOI211_X1 g_46_58 (.ZN (n_46_58), .A (n_50_56), .B (n_56_53), .C1 (n_60_53), .C2 (n_62_50) );
AOI211_X1 g_44_59 (.ZN (n_44_59), .A (n_48_57), .B (n_54_54), .C1 (n_58_52), .C2 (n_60_51) );
AOI211_X1 g_42_60 (.ZN (n_42_60), .A (n_46_58), .B (n_52_55), .C1 (n_56_53), .C2 (n_62_52) );
AOI211_X1 g_43_58 (.ZN (n_43_58), .A (n_44_59), .B (n_50_56), .C1 (n_54_54), .C2 (n_60_53) );
AOI211_X1 g_41_59 (.ZN (n_41_59), .A (n_42_60), .B (n_48_57), .C1 (n_52_55), .C2 (n_58_52) );
AOI211_X1 g_39_60 (.ZN (n_39_60), .A (n_43_58), .B (n_46_58), .C1 (n_50_56), .C2 (n_56_53) );
AOI211_X1 g_37_61 (.ZN (n_37_61), .A (n_41_59), .B (n_44_59), .C1 (n_48_57), .C2 (n_54_54) );
AOI211_X1 g_35_62 (.ZN (n_35_62), .A (n_39_60), .B (n_42_60), .C1 (n_46_58), .C2 (n_52_55) );
AOI211_X1 g_33_63 (.ZN (n_33_63), .A (n_37_61), .B (n_43_58), .C1 (n_44_59), .C2 (n_50_56) );
AOI211_X1 g_31_64 (.ZN (n_31_64), .A (n_35_62), .B (n_41_59), .C1 (n_42_60), .C2 (n_48_57) );
AOI211_X1 g_29_65 (.ZN (n_29_65), .A (n_33_63), .B (n_39_60), .C1 (n_43_58), .C2 (n_46_58) );
AOI211_X1 g_27_66 (.ZN (n_27_66), .A (n_31_64), .B (n_37_61), .C1 (n_41_59), .C2 (n_44_59) );
AOI211_X1 g_25_67 (.ZN (n_25_67), .A (n_29_65), .B (n_35_62), .C1 (n_39_60), .C2 (n_42_60) );
AOI211_X1 g_23_68 (.ZN (n_23_68), .A (n_27_66), .B (n_33_63), .C1 (n_37_61), .C2 (n_43_58) );
AOI211_X1 g_21_69 (.ZN (n_21_69), .A (n_25_67), .B (n_31_64), .C1 (n_35_62), .C2 (n_41_59) );
AOI211_X1 g_19_70 (.ZN (n_19_70), .A (n_23_68), .B (n_29_65), .C1 (n_33_63), .C2 (n_39_60) );
AOI211_X1 g_17_71 (.ZN (n_17_71), .A (n_21_69), .B (n_27_66), .C1 (n_31_64), .C2 (n_37_61) );
AOI211_X1 g_15_70 (.ZN (n_15_70), .A (n_19_70), .B (n_25_67), .C1 (n_29_65), .C2 (n_35_62) );
AOI211_X1 g_13_71 (.ZN (n_13_71), .A (n_17_71), .B (n_23_68), .C1 (n_27_66), .C2 (n_33_63) );
AOI211_X1 g_11_72 (.ZN (n_11_72), .A (n_15_70), .B (n_21_69), .C1 (n_25_67), .C2 (n_31_64) );
AOI211_X1 g_12_74 (.ZN (n_12_74), .A (n_13_71), .B (n_19_70), .C1 (n_23_68), .C2 (n_29_65) );
AOI211_X1 g_14_73 (.ZN (n_14_73), .A (n_11_72), .B (n_17_71), .C1 (n_21_69), .C2 (n_27_66) );
AOI211_X1 g_15_71 (.ZN (n_15_71), .A (n_12_74), .B (n_15_70), .C1 (n_19_70), .C2 (n_25_67) );
AOI211_X1 g_17_70 (.ZN (n_17_70), .A (n_14_73), .B (n_13_71), .C1 (n_17_71), .C2 (n_23_68) );
AOI211_X1 g_16_72 (.ZN (n_16_72), .A (n_15_71), .B (n_11_72), .C1 (n_15_70), .C2 (n_21_69) );
AOI211_X1 g_18_71 (.ZN (n_18_71), .A (n_17_70), .B (n_12_74), .C1 (n_13_71), .C2 (n_19_70) );
AOI211_X1 g_20_70 (.ZN (n_20_70), .A (n_16_72), .B (n_14_73), .C1 (n_11_72), .C2 (n_17_71) );
AOI211_X1 g_22_69 (.ZN (n_22_69), .A (n_18_71), .B (n_15_71), .C1 (n_12_74), .C2 (n_15_70) );
AOI211_X1 g_24_68 (.ZN (n_24_68), .A (n_20_70), .B (n_17_70), .C1 (n_14_73), .C2 (n_13_71) );
AOI211_X1 g_26_67 (.ZN (n_26_67), .A (n_22_69), .B (n_16_72), .C1 (n_15_71), .C2 (n_11_72) );
AOI211_X1 g_25_69 (.ZN (n_25_69), .A (n_24_68), .B (n_18_71), .C1 (n_17_70), .C2 (n_12_74) );
AOI211_X1 g_27_68 (.ZN (n_27_68), .A (n_26_67), .B (n_20_70), .C1 (n_16_72), .C2 (n_14_73) );
AOI211_X1 g_29_67 (.ZN (n_29_67), .A (n_25_69), .B (n_22_69), .C1 (n_18_71), .C2 (n_15_71) );
AOI211_X1 g_31_66 (.ZN (n_31_66), .A (n_27_68), .B (n_24_68), .C1 (n_20_70), .C2 (n_17_70) );
AOI211_X1 g_33_65 (.ZN (n_33_65), .A (n_29_67), .B (n_26_67), .C1 (n_22_69), .C2 (n_16_72) );
AOI211_X1 g_35_64 (.ZN (n_35_64), .A (n_31_66), .B (n_25_69), .C1 (n_24_68), .C2 (n_18_71) );
AOI211_X1 g_37_63 (.ZN (n_37_63), .A (n_33_65), .B (n_27_68), .C1 (n_26_67), .C2 (n_20_70) );
AOI211_X1 g_39_62 (.ZN (n_39_62), .A (n_35_64), .B (n_29_67), .C1 (n_25_69), .C2 (n_22_69) );
AOI211_X1 g_41_61 (.ZN (n_41_61), .A (n_37_63), .B (n_31_66), .C1 (n_27_68), .C2 (n_24_68) );
AOI211_X1 g_43_60 (.ZN (n_43_60), .A (n_39_62), .B (n_33_65), .C1 (n_29_67), .C2 (n_26_67) );
AOI211_X1 g_45_59 (.ZN (n_45_59), .A (n_41_61), .B (n_35_64), .C1 (n_31_66), .C2 (n_25_69) );
AOI211_X1 g_44_61 (.ZN (n_44_61), .A (n_43_60), .B (n_37_63), .C1 (n_33_65), .C2 (n_27_68) );
AOI211_X1 g_46_60 (.ZN (n_46_60), .A (n_45_59), .B (n_39_62), .C1 (n_35_64), .C2 (n_29_67) );
AOI211_X1 g_48_59 (.ZN (n_48_59), .A (n_44_61), .B (n_41_61), .C1 (n_37_63), .C2 (n_31_66) );
AOI211_X1 g_50_58 (.ZN (n_50_58), .A (n_46_60), .B (n_43_60), .C1 (n_39_62), .C2 (n_33_65) );
AOI211_X1 g_52_57 (.ZN (n_52_57), .A (n_48_59), .B (n_45_59), .C1 (n_41_61), .C2 (n_35_64) );
AOI211_X1 g_54_56 (.ZN (n_54_56), .A (n_50_58), .B (n_44_61), .C1 (n_43_60), .C2 (n_37_63) );
AOI211_X1 g_56_55 (.ZN (n_56_55), .A (n_52_57), .B (n_46_60), .C1 (n_45_59), .C2 (n_39_62) );
AOI211_X1 g_58_54 (.ZN (n_58_54), .A (n_54_56), .B (n_48_59), .C1 (n_44_61), .C2 (n_41_61) );
AOI211_X1 g_57_56 (.ZN (n_57_56), .A (n_56_55), .B (n_50_58), .C1 (n_46_60), .C2 (n_43_60) );
AOI211_X1 g_55_55 (.ZN (n_55_55), .A (n_58_54), .B (n_52_57), .C1 (n_48_59), .C2 (n_45_59) );
AOI211_X1 g_57_54 (.ZN (n_57_54), .A (n_57_56), .B (n_54_56), .C1 (n_50_58), .C2 (n_44_61) );
AOI211_X1 g_59_53 (.ZN (n_59_53), .A (n_55_55), .B (n_56_55), .C1 (n_52_57), .C2 (n_46_60) );
AOI211_X1 g_61_52 (.ZN (n_61_52), .A (n_57_54), .B (n_58_54), .C1 (n_54_56), .C2 (n_48_59) );
AOI211_X1 g_62_54 (.ZN (n_62_54), .A (n_59_53), .B (n_57_56), .C1 (n_56_55), .C2 (n_50_58) );
AOI211_X1 g_60_55 (.ZN (n_60_55), .A (n_61_52), .B (n_55_55), .C1 (n_58_54), .C2 (n_52_57) );
AOI211_X1 g_61_53 (.ZN (n_61_53), .A (n_62_54), .B (n_57_54), .C1 (n_57_56), .C2 (n_54_56) );
AOI211_X1 g_59_54 (.ZN (n_59_54), .A (n_60_55), .B (n_59_53), .C1 (n_55_55), .C2 (n_56_55) );
AOI211_X1 g_57_55 (.ZN (n_57_55), .A (n_61_53), .B (n_61_52), .C1 (n_57_54), .C2 (n_58_54) );
AOI211_X1 g_55_56 (.ZN (n_55_56), .A (n_59_54), .B (n_62_54), .C1 (n_59_53), .C2 (n_57_56) );
AOI211_X1 g_53_57 (.ZN (n_53_57), .A (n_57_55), .B (n_60_55), .C1 (n_61_52), .C2 (n_55_55) );
AOI211_X1 g_51_58 (.ZN (n_51_58), .A (n_55_56), .B (n_61_53), .C1 (n_62_54), .C2 (n_57_54) );
AOI211_X1 g_49_59 (.ZN (n_49_59), .A (n_53_57), .B (n_59_54), .C1 (n_60_55), .C2 (n_59_53) );
AOI211_X1 g_47_60 (.ZN (n_47_60), .A (n_51_58), .B (n_57_55), .C1 (n_61_53), .C2 (n_61_52) );
AOI211_X1 g_45_61 (.ZN (n_45_61), .A (n_49_59), .B (n_55_56), .C1 (n_59_54), .C2 (n_62_54) );
AOI211_X1 g_43_62 (.ZN (n_43_62), .A (n_47_60), .B (n_53_57), .C1 (n_57_55), .C2 (n_60_55) );
AOI211_X1 g_44_60 (.ZN (n_44_60), .A (n_45_61), .B (n_51_58), .C1 (n_55_56), .C2 (n_61_53) );
AOI211_X1 g_42_61 (.ZN (n_42_61), .A (n_43_62), .B (n_49_59), .C1 (n_53_57), .C2 (n_59_54) );
AOI211_X1 g_40_62 (.ZN (n_40_62), .A (n_44_60), .B (n_47_60), .C1 (n_51_58), .C2 (n_57_55) );
AOI211_X1 g_41_60 (.ZN (n_41_60), .A (n_42_61), .B (n_45_61), .C1 (n_49_59), .C2 (n_55_56) );
AOI211_X1 g_39_61 (.ZN (n_39_61), .A (n_40_62), .B (n_43_62), .C1 (n_47_60), .C2 (n_53_57) );
AOI211_X1 g_37_62 (.ZN (n_37_62), .A (n_41_60), .B (n_44_60), .C1 (n_45_61), .C2 (n_51_58) );
AOI211_X1 g_35_63 (.ZN (n_35_63), .A (n_39_61), .B (n_42_61), .C1 (n_43_62), .C2 (n_49_59) );
AOI211_X1 g_33_64 (.ZN (n_33_64), .A (n_37_62), .B (n_40_62), .C1 (n_44_60), .C2 (n_47_60) );
AOI211_X1 g_31_65 (.ZN (n_31_65), .A (n_35_63), .B (n_41_60), .C1 (n_42_61), .C2 (n_45_61) );
AOI211_X1 g_29_66 (.ZN (n_29_66), .A (n_33_64), .B (n_39_61), .C1 (n_40_62), .C2 (n_43_62) );
AOI211_X1 g_27_67 (.ZN (n_27_67), .A (n_31_65), .B (n_37_62), .C1 (n_41_60), .C2 (n_44_60) );
AOI211_X1 g_25_68 (.ZN (n_25_68), .A (n_29_66), .B (n_35_63), .C1 (n_39_61), .C2 (n_42_61) );
AOI211_X1 g_23_69 (.ZN (n_23_69), .A (n_27_67), .B (n_33_64), .C1 (n_37_62), .C2 (n_40_62) );
AOI211_X1 g_22_71 (.ZN (n_22_71), .A (n_25_68), .B (n_31_65), .C1 (n_35_63), .C2 (n_41_60) );
AOI211_X1 g_24_70 (.ZN (n_24_70), .A (n_23_69), .B (n_29_66), .C1 (n_33_64), .C2 (n_39_61) );
AOI211_X1 g_26_69 (.ZN (n_26_69), .A (n_22_71), .B (n_27_67), .C1 (n_31_65), .C2 (n_37_62) );
AOI211_X1 g_28_68 (.ZN (n_28_68), .A (n_24_70), .B (n_25_68), .C1 (n_29_66), .C2 (n_35_63) );
AOI211_X1 g_30_67 (.ZN (n_30_67), .A (n_26_69), .B (n_23_69), .C1 (n_27_67), .C2 (n_33_64) );
AOI211_X1 g_32_66 (.ZN (n_32_66), .A (n_28_68), .B (n_22_71), .C1 (n_25_68), .C2 (n_31_65) );
AOI211_X1 g_34_65 (.ZN (n_34_65), .A (n_30_67), .B (n_24_70), .C1 (n_23_69), .C2 (n_29_66) );
AOI211_X1 g_36_64 (.ZN (n_36_64), .A (n_32_66), .B (n_26_69), .C1 (n_22_71), .C2 (n_27_67) );
AOI211_X1 g_38_63 (.ZN (n_38_63), .A (n_34_65), .B (n_28_68), .C1 (n_24_70), .C2 (n_25_68) );
AOI211_X1 g_37_65 (.ZN (n_37_65), .A (n_36_64), .B (n_30_67), .C1 (n_26_69), .C2 (n_23_69) );
AOI211_X1 g_36_63 (.ZN (n_36_63), .A (n_38_63), .B (n_32_66), .C1 (n_28_68), .C2 (n_22_71) );
AOI211_X1 g_38_62 (.ZN (n_38_62), .A (n_37_65), .B (n_34_65), .C1 (n_30_67), .C2 (n_24_70) );
AOI211_X1 g_40_61 (.ZN (n_40_61), .A (n_36_63), .B (n_36_64), .C1 (n_32_66), .C2 (n_26_69) );
AOI211_X1 g_41_63 (.ZN (n_41_63), .A (n_38_62), .B (n_38_63), .C1 (n_34_65), .C2 (n_28_68) );
AOI211_X1 g_39_64 (.ZN (n_39_64), .A (n_40_61), .B (n_37_65), .C1 (n_36_64), .C2 (n_30_67) );
AOI211_X1 g_38_66 (.ZN (n_38_66), .A (n_41_63), .B (n_36_63), .C1 (n_38_63), .C2 (n_32_66) );
AOI211_X1 g_37_64 (.ZN (n_37_64), .A (n_39_64), .B (n_38_62), .C1 (n_37_65), .C2 (n_34_65) );
AOI211_X1 g_39_63 (.ZN (n_39_63), .A (n_38_66), .B (n_40_61), .C1 (n_36_63), .C2 (n_36_64) );
AOI211_X1 g_41_62 (.ZN (n_41_62), .A (n_37_64), .B (n_41_63), .C1 (n_38_62), .C2 (n_38_63) );
AOI211_X1 g_43_61 (.ZN (n_43_61), .A (n_39_63), .B (n_39_64), .C1 (n_40_61), .C2 (n_37_65) );
AOI211_X1 g_45_60 (.ZN (n_45_60), .A (n_41_62), .B (n_38_66), .C1 (n_41_63), .C2 (n_36_63) );
AOI211_X1 g_47_59 (.ZN (n_47_59), .A (n_43_61), .B (n_37_64), .C1 (n_39_64), .C2 (n_38_62) );
AOI211_X1 g_49_58 (.ZN (n_49_58), .A (n_45_60), .B (n_39_63), .C1 (n_38_66), .C2 (n_40_61) );
AOI211_X1 g_51_57 (.ZN (n_51_57), .A (n_47_59), .B (n_41_62), .C1 (n_37_64), .C2 (n_41_63) );
AOI211_X1 g_53_56 (.ZN (n_53_56), .A (n_49_58), .B (n_43_61), .C1 (n_39_63), .C2 (n_39_64) );
AOI211_X1 g_55_57 (.ZN (n_55_57), .A (n_51_57), .B (n_45_60), .C1 (n_41_62), .C2 (n_38_66) );
AOI211_X1 g_53_58 (.ZN (n_53_58), .A (n_53_56), .B (n_47_59), .C1 (n_43_61), .C2 (n_37_64) );
AOI211_X1 g_51_59 (.ZN (n_51_59), .A (n_55_57), .B (n_49_58), .C1 (n_45_60), .C2 (n_39_63) );
AOI211_X1 g_49_60 (.ZN (n_49_60), .A (n_53_58), .B (n_51_57), .C1 (n_47_59), .C2 (n_41_62) );
AOI211_X1 g_47_61 (.ZN (n_47_61), .A (n_51_59), .B (n_53_56), .C1 (n_49_58), .C2 (n_43_61) );
AOI211_X1 g_45_62 (.ZN (n_45_62), .A (n_49_60), .B (n_55_57), .C1 (n_51_57), .C2 (n_45_60) );
AOI211_X1 g_43_63 (.ZN (n_43_63), .A (n_47_61), .B (n_53_58), .C1 (n_53_56), .C2 (n_47_59) );
AOI211_X1 g_41_64 (.ZN (n_41_64), .A (n_45_62), .B (n_51_59), .C1 (n_55_57), .C2 (n_49_58) );
AOI211_X1 g_42_62 (.ZN (n_42_62), .A (n_43_63), .B (n_49_60), .C1 (n_53_58), .C2 (n_51_57) );
AOI211_X1 g_40_63 (.ZN (n_40_63), .A (n_41_64), .B (n_47_61), .C1 (n_51_59), .C2 (n_53_56) );
AOI211_X1 g_38_64 (.ZN (n_38_64), .A (n_42_62), .B (n_45_62), .C1 (n_49_60), .C2 (n_55_57) );
AOI211_X1 g_36_65 (.ZN (n_36_65), .A (n_40_63), .B (n_43_63), .C1 (n_47_61), .C2 (n_53_58) );
AOI211_X1 g_34_64 (.ZN (n_34_64), .A (n_38_64), .B (n_41_64), .C1 (n_45_62), .C2 (n_51_59) );
AOI211_X1 g_32_65 (.ZN (n_32_65), .A (n_36_65), .B (n_42_62), .C1 (n_43_63), .C2 (n_49_60) );
AOI211_X1 g_30_66 (.ZN (n_30_66), .A (n_34_64), .B (n_40_63), .C1 (n_41_64), .C2 (n_47_61) );
AOI211_X1 g_28_67 (.ZN (n_28_67), .A (n_32_65), .B (n_38_64), .C1 (n_42_62), .C2 (n_45_62) );
AOI211_X1 g_26_68 (.ZN (n_26_68), .A (n_30_66), .B (n_36_65), .C1 (n_40_63), .C2 (n_43_63) );
AOI211_X1 g_24_69 (.ZN (n_24_69), .A (n_28_67), .B (n_34_64), .C1 (n_38_64), .C2 (n_41_64) );
AOI211_X1 g_22_70 (.ZN (n_22_70), .A (n_26_68), .B (n_32_65), .C1 (n_36_65), .C2 (n_42_62) );
AOI211_X1 g_20_71 (.ZN (n_20_71), .A (n_24_69), .B (n_30_66), .C1 (n_34_64), .C2 (n_40_63) );
AOI211_X1 g_18_72 (.ZN (n_18_72), .A (n_22_70), .B (n_28_67), .C1 (n_32_65), .C2 (n_38_64) );
AOI211_X1 g_16_71 (.ZN (n_16_71), .A (n_20_71), .B (n_26_68), .C1 (n_30_66), .C2 (n_36_65) );
AOI211_X1 g_14_72 (.ZN (n_14_72), .A (n_18_72), .B (n_24_69), .C1 (n_28_67), .C2 (n_34_64) );
AOI211_X1 g_12_71 (.ZN (n_12_71), .A (n_16_71), .B (n_22_70), .C1 (n_26_68), .C2 (n_32_65) );
AOI211_X1 g_10_72 (.ZN (n_10_72), .A (n_14_72), .B (n_20_71), .C1 (n_24_69), .C2 (n_30_66) );
AOI211_X1 g_8_73 (.ZN (n_8_73), .A (n_12_71), .B (n_18_72), .C1 (n_22_70), .C2 (n_28_67) );
AOI211_X1 g_6_74 (.ZN (n_6_74), .A (n_10_72), .B (n_16_71), .C1 (n_20_71), .C2 (n_26_68) );
AOI211_X1 g_5_76 (.ZN (n_5_76), .A (n_8_73), .B (n_14_72), .C1 (n_18_72), .C2 (n_24_69) );
AOI211_X1 g_7_75 (.ZN (n_7_75), .A (n_6_74), .B (n_12_71), .C1 (n_16_71), .C2 (n_22_70) );
AOI211_X1 g_9_74 (.ZN (n_9_74), .A (n_5_76), .B (n_10_72), .C1 (n_14_72), .C2 (n_20_71) );
AOI211_X1 g_7_73 (.ZN (n_7_73), .A (n_7_75), .B (n_8_73), .C1 (n_12_71), .C2 (n_18_72) );
AOI211_X1 g_6_75 (.ZN (n_6_75), .A (n_9_74), .B (n_6_74), .C1 (n_10_72), .C2 (n_16_71) );
AOI211_X1 g_8_74 (.ZN (n_8_74), .A (n_7_73), .B (n_5_76), .C1 (n_8_73), .C2 (n_14_72) );
AOI211_X1 g_7_76 (.ZN (n_7_76), .A (n_6_75), .B (n_7_75), .C1 (n_6_74), .C2 (n_12_71) );
AOI211_X1 g_5_77 (.ZN (n_5_77), .A (n_8_74), .B (n_9_74), .C1 (n_5_76), .C2 (n_10_72) );
AOI211_X1 g_4_79 (.ZN (n_4_79), .A (n_7_76), .B (n_7_73), .C1 (n_7_75), .C2 (n_8_73) );
AOI211_X1 g_6_78 (.ZN (n_6_78), .A (n_5_77), .B (n_6_75), .C1 (n_9_74), .C2 (n_6_74) );
AOI211_X1 g_8_77 (.ZN (n_8_77), .A (n_4_79), .B (n_8_74), .C1 (n_7_73), .C2 (n_5_76) );
AOI211_X1 g_9_75 (.ZN (n_9_75), .A (n_6_78), .B (n_7_76), .C1 (n_6_75), .C2 (n_7_75) );
AOI211_X1 g_11_74 (.ZN (n_11_74), .A (n_8_77), .B (n_5_77), .C1 (n_8_74), .C2 (n_9_74) );
AOI211_X1 g_13_73 (.ZN (n_13_73), .A (n_9_75), .B (n_4_79), .C1 (n_7_76), .C2 (n_7_73) );
AOI211_X1 g_15_72 (.ZN (n_15_72), .A (n_11_74), .B (n_6_78), .C1 (n_5_77), .C2 (n_6_75) );
AOI211_X1 g_17_73 (.ZN (n_17_73), .A (n_13_73), .B (n_8_77), .C1 (n_4_79), .C2 (n_8_74) );
AOI211_X1 g_19_72 (.ZN (n_19_72), .A (n_15_72), .B (n_9_75), .C1 (n_6_78), .C2 (n_7_76) );
AOI211_X1 g_21_71 (.ZN (n_21_71), .A (n_17_73), .B (n_11_74), .C1 (n_8_77), .C2 (n_5_77) );
AOI211_X1 g_23_70 (.ZN (n_23_70), .A (n_19_72), .B (n_13_73), .C1 (n_9_75), .C2 (n_4_79) );
AOI211_X1 g_22_72 (.ZN (n_22_72), .A (n_21_71), .B (n_15_72), .C1 (n_11_74), .C2 (n_6_78) );
AOI211_X1 g_24_71 (.ZN (n_24_71), .A (n_23_70), .B (n_17_73), .C1 (n_13_73), .C2 (n_8_77) );
AOI211_X1 g_26_70 (.ZN (n_26_70), .A (n_22_72), .B (n_19_72), .C1 (n_15_72), .C2 (n_9_75) );
AOI211_X1 g_28_69 (.ZN (n_28_69), .A (n_24_71), .B (n_21_71), .C1 (n_17_73), .C2 (n_11_74) );
AOI211_X1 g_30_68 (.ZN (n_30_68), .A (n_26_70), .B (n_23_70), .C1 (n_19_72), .C2 (n_13_73) );
AOI211_X1 g_32_67 (.ZN (n_32_67), .A (n_28_69), .B (n_22_72), .C1 (n_21_71), .C2 (n_15_72) );
AOI211_X1 g_34_66 (.ZN (n_34_66), .A (n_30_68), .B (n_24_71), .C1 (n_23_70), .C2 (n_17_73) );
AOI211_X1 g_36_67 (.ZN (n_36_67), .A (n_32_67), .B (n_26_70), .C1 (n_22_72), .C2 (n_19_72) );
AOI211_X1 g_35_65 (.ZN (n_35_65), .A (n_34_66), .B (n_28_69), .C1 (n_24_71), .C2 (n_21_71) );
AOI211_X1 g_33_66 (.ZN (n_33_66), .A (n_36_67), .B (n_30_68), .C1 (n_26_70), .C2 (n_23_70) );
AOI211_X1 g_31_67 (.ZN (n_31_67), .A (n_35_65), .B (n_32_67), .C1 (n_28_69), .C2 (n_22_72) );
AOI211_X1 g_29_68 (.ZN (n_29_68), .A (n_33_66), .B (n_34_66), .C1 (n_30_68), .C2 (n_24_71) );
AOI211_X1 g_27_69 (.ZN (n_27_69), .A (n_31_67), .B (n_36_67), .C1 (n_32_67), .C2 (n_26_70) );
AOI211_X1 g_25_70 (.ZN (n_25_70), .A (n_29_68), .B (n_35_65), .C1 (n_34_66), .C2 (n_28_69) );
AOI211_X1 g_23_71 (.ZN (n_23_71), .A (n_27_69), .B (n_33_66), .C1 (n_36_67), .C2 (n_30_68) );
AOI211_X1 g_21_72 (.ZN (n_21_72), .A (n_25_70), .B (n_31_67), .C1 (n_35_65), .C2 (n_32_67) );
AOI211_X1 g_19_71 (.ZN (n_19_71), .A (n_23_71), .B (n_29_68), .C1 (n_33_66), .C2 (n_34_66) );
AOI211_X1 g_17_72 (.ZN (n_17_72), .A (n_21_72), .B (n_27_69), .C1 (n_31_67), .C2 (n_36_67) );
AOI211_X1 g_15_73 (.ZN (n_15_73), .A (n_19_71), .B (n_25_70), .C1 (n_29_68), .C2 (n_35_65) );
AOI211_X1 g_13_74 (.ZN (n_13_74), .A (n_17_72), .B (n_23_71), .C1 (n_27_69), .C2 (n_33_66) );
AOI211_X1 g_11_73 (.ZN (n_11_73), .A (n_15_73), .B (n_21_72), .C1 (n_25_70), .C2 (n_31_67) );
AOI211_X1 g_10_75 (.ZN (n_10_75), .A (n_13_74), .B (n_19_71), .C1 (n_23_71), .C2 (n_29_68) );
AOI211_X1 g_8_76 (.ZN (n_8_76), .A (n_11_73), .B (n_17_72), .C1 (n_21_72), .C2 (n_27_69) );
AOI211_X1 g_6_77 (.ZN (n_6_77), .A (n_10_75), .B (n_15_73), .C1 (n_19_71), .C2 (n_25_70) );
AOI211_X1 g_4_78 (.ZN (n_4_78), .A (n_8_76), .B (n_13_74), .C1 (n_17_72), .C2 (n_23_71) );
AOI211_X1 g_3_80 (.ZN (n_3_80), .A (n_6_77), .B (n_11_73), .C1 (n_15_73), .C2 (n_21_72) );
AOI211_X1 g_2_82 (.ZN (n_2_82), .A (n_4_78), .B (n_10_75), .C1 (n_13_74), .C2 (n_19_71) );
AOI211_X1 g_4_81 (.ZN (n_4_81), .A (n_3_80), .B (n_8_76), .C1 (n_11_73), .C2 (n_17_72) );
AOI211_X1 g_5_79 (.ZN (n_5_79), .A (n_2_82), .B (n_6_77), .C1 (n_10_75), .C2 (n_15_73) );
AOI211_X1 g_7_78 (.ZN (n_7_78), .A (n_4_81), .B (n_4_78), .C1 (n_8_76), .C2 (n_13_74) );
AOI211_X1 g_6_80 (.ZN (n_6_80), .A (n_5_79), .B (n_3_80), .C1 (n_6_77), .C2 (n_11_73) );
AOI211_X1 g_8_79 (.ZN (n_8_79), .A (n_7_78), .B (n_2_82), .C1 (n_4_78), .C2 (n_10_75) );
AOI211_X1 g_9_77 (.ZN (n_9_77), .A (n_6_80), .B (n_4_81), .C1 (n_3_80), .C2 (n_8_76) );
AOI211_X1 g_8_75 (.ZN (n_8_75), .A (n_8_79), .B (n_5_79), .C1 (n_2_82), .C2 (n_6_77) );
AOI211_X1 g_7_77 (.ZN (n_7_77), .A (n_9_77), .B (n_7_78), .C1 (n_4_81), .C2 (n_4_78) );
AOI211_X1 g_6_79 (.ZN (n_6_79), .A (n_8_75), .B (n_6_80), .C1 (n_5_79), .C2 (n_3_80) );
AOI211_X1 g_5_81 (.ZN (n_5_81), .A (n_7_77), .B (n_8_79), .C1 (n_7_78), .C2 (n_2_82) );
AOI211_X1 g_4_83 (.ZN (n_4_83), .A (n_6_79), .B (n_9_77), .C1 (n_6_80), .C2 (n_4_81) );
AOI211_X1 g_6_84 (.ZN (n_6_84), .A (n_5_81), .B (n_8_75), .C1 (n_8_79), .C2 (n_5_79) );
AOI211_X1 g_4_85 (.ZN (n_4_85), .A (n_4_83), .B (n_7_77), .C1 (n_9_77), .C2 (n_7_78) );
AOI211_X1 g_2_86 (.ZN (n_2_86), .A (n_6_84), .B (n_6_79), .C1 (n_8_75), .C2 (n_6_80) );
AOI211_X1 g_3_84 (.ZN (n_3_84), .A (n_4_85), .B (n_5_81), .C1 (n_7_77), .C2 (n_8_79) );
AOI211_X1 g_5_83 (.ZN (n_5_83), .A (n_2_86), .B (n_4_83), .C1 (n_6_79), .C2 (n_9_77) );
AOI211_X1 g_7_82 (.ZN (n_7_82), .A (n_3_84), .B (n_6_84), .C1 (n_5_81), .C2 (n_8_75) );
AOI211_X1 g_8_80 (.ZN (n_8_80), .A (n_5_83), .B (n_4_85), .C1 (n_4_83), .C2 (n_7_77) );
AOI211_X1 g_6_81 (.ZN (n_6_81), .A (n_7_82), .B (n_2_86), .C1 (n_6_84), .C2 (n_6_79) );
AOI211_X1 g_4_82 (.ZN (n_4_82), .A (n_8_80), .B (n_3_84), .C1 (n_4_85), .C2 (n_5_81) );
AOI211_X1 g_5_80 (.ZN (n_5_80), .A (n_6_81), .B (n_5_83), .C1 (n_2_86), .C2 (n_4_83) );
AOI211_X1 g_7_79 (.ZN (n_7_79), .A (n_4_82), .B (n_7_82), .C1 (n_3_84), .C2 (n_6_84) );
AOI211_X1 g_9_78 (.ZN (n_9_78), .A (n_5_80), .B (n_8_80), .C1 (n_5_83), .C2 (n_4_85) );
AOI211_X1 g_10_76 (.ZN (n_10_76), .A (n_7_79), .B (n_6_81), .C1 (n_7_82), .C2 (n_2_86) );
AOI211_X1 g_12_75 (.ZN (n_12_75), .A (n_9_78), .B (n_4_82), .C1 (n_8_80), .C2 (n_3_84) );
AOI211_X1 g_10_74 (.ZN (n_10_74), .A (n_10_76), .B (n_5_80), .C1 (n_6_81), .C2 (n_5_83) );
AOI211_X1 g_12_73 (.ZN (n_12_73), .A (n_12_75), .B (n_7_79), .C1 (n_4_82), .C2 (n_7_82) );
AOI211_X1 g_11_75 (.ZN (n_11_75), .A (n_10_74), .B (n_9_78), .C1 (n_5_80), .C2 (n_8_80) );
AOI211_X1 g_9_76 (.ZN (n_9_76), .A (n_12_73), .B (n_10_76), .C1 (n_7_79), .C2 (n_6_81) );
AOI211_X1 g_8_78 (.ZN (n_8_78), .A (n_11_75), .B (n_12_75), .C1 (n_9_78), .C2 (n_4_82) );
AOI211_X1 g_10_77 (.ZN (n_10_77), .A (n_9_76), .B (n_10_74), .C1 (n_10_76), .C2 (n_5_80) );
AOI211_X1 g_12_76 (.ZN (n_12_76), .A (n_8_78), .B (n_12_73), .C1 (n_12_75), .C2 (n_7_79) );
AOI211_X1 g_14_75 (.ZN (n_14_75), .A (n_10_77), .B (n_11_75), .C1 (n_10_74), .C2 (n_9_78) );
AOI211_X1 g_16_74 (.ZN (n_16_74), .A (n_12_76), .B (n_9_76), .C1 (n_12_73), .C2 (n_10_76) );
AOI211_X1 g_18_73 (.ZN (n_18_73), .A (n_14_75), .B (n_8_78), .C1 (n_11_75), .C2 (n_12_75) );
AOI211_X1 g_20_72 (.ZN (n_20_72), .A (n_16_74), .B (n_10_77), .C1 (n_9_76), .C2 (n_10_74) );
AOI211_X1 g_19_74 (.ZN (n_19_74), .A (n_18_73), .B (n_12_76), .C1 (n_8_78), .C2 (n_12_73) );
AOI211_X1 g_21_73 (.ZN (n_21_73), .A (n_20_72), .B (n_14_75), .C1 (n_10_77), .C2 (n_11_75) );
AOI211_X1 g_23_72 (.ZN (n_23_72), .A (n_19_74), .B (n_16_74), .C1 (n_12_76), .C2 (n_9_76) );
AOI211_X1 g_25_71 (.ZN (n_25_71), .A (n_21_73), .B (n_18_73), .C1 (n_14_75), .C2 (n_8_78) );
AOI211_X1 g_27_70 (.ZN (n_27_70), .A (n_23_72), .B (n_20_72), .C1 (n_16_74), .C2 (n_10_77) );
AOI211_X1 g_29_69 (.ZN (n_29_69), .A (n_25_71), .B (n_19_74), .C1 (n_18_73), .C2 (n_12_76) );
AOI211_X1 g_31_68 (.ZN (n_31_68), .A (n_27_70), .B (n_21_73), .C1 (n_20_72), .C2 (n_14_75) );
AOI211_X1 g_33_67 (.ZN (n_33_67), .A (n_29_69), .B (n_23_72), .C1 (n_19_74), .C2 (n_16_74) );
AOI211_X1 g_35_66 (.ZN (n_35_66), .A (n_31_68), .B (n_25_71), .C1 (n_21_73), .C2 (n_18_73) );
AOI211_X1 g_34_68 (.ZN (n_34_68), .A (n_33_67), .B (n_27_70), .C1 (n_23_72), .C2 (n_20_72) );
AOI211_X1 g_32_69 (.ZN (n_32_69), .A (n_35_66), .B (n_29_69), .C1 (n_25_71), .C2 (n_19_74) );
AOI211_X1 g_30_70 (.ZN (n_30_70), .A (n_34_68), .B (n_31_68), .C1 (n_27_70), .C2 (n_21_73) );
AOI211_X1 g_28_71 (.ZN (n_28_71), .A (n_32_69), .B (n_33_67), .C1 (n_29_69), .C2 (n_23_72) );
AOI211_X1 g_26_72 (.ZN (n_26_72), .A (n_30_70), .B (n_35_66), .C1 (n_31_68), .C2 (n_25_71) );
AOI211_X1 g_24_73 (.ZN (n_24_73), .A (n_28_71), .B (n_34_68), .C1 (n_33_67), .C2 (n_27_70) );
AOI211_X1 g_22_74 (.ZN (n_22_74), .A (n_26_72), .B (n_32_69), .C1 (n_35_66), .C2 (n_29_69) );
AOI211_X1 g_20_73 (.ZN (n_20_73), .A (n_24_73), .B (n_30_70), .C1 (n_34_68), .C2 (n_31_68) );
AOI211_X1 g_18_74 (.ZN (n_18_74), .A (n_22_74), .B (n_28_71), .C1 (n_32_69), .C2 (n_33_67) );
AOI211_X1 g_16_73 (.ZN (n_16_73), .A (n_20_73), .B (n_26_72), .C1 (n_30_70), .C2 (n_35_66) );
AOI211_X1 g_14_74 (.ZN (n_14_74), .A (n_18_74), .B (n_24_73), .C1 (n_28_71), .C2 (n_34_68) );
AOI211_X1 g_16_75 (.ZN (n_16_75), .A (n_16_73), .B (n_22_74), .C1 (n_26_72), .C2 (n_32_69) );
AOI211_X1 g_14_76 (.ZN (n_14_76), .A (n_14_74), .B (n_20_73), .C1 (n_24_73), .C2 (n_30_70) );
AOI211_X1 g_15_74 (.ZN (n_15_74), .A (n_16_75), .B (n_18_74), .C1 (n_22_74), .C2 (n_28_71) );
AOI211_X1 g_13_75 (.ZN (n_13_75), .A (n_14_76), .B (n_16_73), .C1 (n_20_73), .C2 (n_26_72) );
AOI211_X1 g_11_76 (.ZN (n_11_76), .A (n_15_74), .B (n_14_74), .C1 (n_18_74), .C2 (n_24_73) );
AOI211_X1 g_10_78 (.ZN (n_10_78), .A (n_13_75), .B (n_16_75), .C1 (n_16_73), .C2 (n_22_74) );
AOI211_X1 g_12_77 (.ZN (n_12_77), .A (n_11_76), .B (n_14_76), .C1 (n_14_74), .C2 (n_20_73) );
AOI211_X1 g_11_79 (.ZN (n_11_79), .A (n_10_78), .B (n_15_74), .C1 (n_16_75), .C2 (n_18_74) );
AOI211_X1 g_9_80 (.ZN (n_9_80), .A (n_12_77), .B (n_13_75), .C1 (n_14_76), .C2 (n_16_73) );
AOI211_X1 g_7_81 (.ZN (n_7_81), .A (n_11_79), .B (n_11_76), .C1 (n_15_74), .C2 (n_14_74) );
AOI211_X1 g_6_83 (.ZN (n_6_83), .A (n_9_80), .B (n_10_78), .C1 (n_13_75), .C2 (n_16_75) );
AOI211_X1 g_5_85 (.ZN (n_5_85), .A (n_7_81), .B (n_12_77), .C1 (n_11_76), .C2 (n_14_76) );
AOI211_X1 g_4_87 (.ZN (n_4_87), .A (n_6_83), .B (n_11_79), .C1 (n_10_78), .C2 (n_15_74) );
AOI211_X1 g_6_88 (.ZN (n_6_88), .A (n_5_85), .B (n_9_80), .C1 (n_12_77), .C2 (n_13_75) );
AOI211_X1 g_4_89 (.ZN (n_4_89), .A (n_4_87), .B (n_7_81), .C1 (n_11_79), .C2 (n_11_76) );
AOI211_X1 g_2_90 (.ZN (n_2_90), .A (n_6_88), .B (n_6_83), .C1 (n_9_80), .C2 (n_10_78) );
AOI211_X1 g_3_88 (.ZN (n_3_88), .A (n_4_89), .B (n_5_85), .C1 (n_7_81), .C2 (n_12_77) );
AOI211_X1 g_5_87 (.ZN (n_5_87), .A (n_2_90), .B (n_4_87), .C1 (n_6_83), .C2 (n_11_79) );
AOI211_X1 g_7_86 (.ZN (n_7_86), .A (n_3_88), .B (n_6_88), .C1 (n_5_85), .C2 (n_9_80) );
AOI211_X1 g_8_84 (.ZN (n_8_84), .A (n_5_87), .B (n_4_89), .C1 (n_4_87), .C2 (n_7_81) );
AOI211_X1 g_6_85 (.ZN (n_6_85), .A (n_7_86), .B (n_2_90), .C1 (n_6_88), .C2 (n_6_83) );
AOI211_X1 g_4_86 (.ZN (n_4_86), .A (n_8_84), .B (n_3_88), .C1 (n_4_89), .C2 (n_5_85) );
AOI211_X1 g_5_84 (.ZN (n_5_84), .A (n_6_85), .B (n_5_87), .C1 (n_2_90), .C2 (n_4_87) );
AOI211_X1 g_7_83 (.ZN (n_7_83), .A (n_4_86), .B (n_7_86), .C1 (n_3_88), .C2 (n_6_88) );
AOI211_X1 g_9_82 (.ZN (n_9_82), .A (n_5_84), .B (n_8_84), .C1 (n_5_87), .C2 (n_4_89) );
AOI211_X1 g_10_80 (.ZN (n_10_80), .A (n_7_83), .B (n_6_85), .C1 (n_7_86), .C2 (n_2_90) );
AOI211_X1 g_11_78 (.ZN (n_11_78), .A (n_9_82), .B (n_4_86), .C1 (n_8_84), .C2 (n_3_88) );
AOI211_X1 g_13_77 (.ZN (n_13_77), .A (n_10_80), .B (n_5_84), .C1 (n_6_85), .C2 (n_5_87) );
AOI211_X1 g_15_76 (.ZN (n_15_76), .A (n_11_78), .B (n_7_83), .C1 (n_4_86), .C2 (n_7_86) );
AOI211_X1 g_17_75 (.ZN (n_17_75), .A (n_13_77), .B (n_9_82), .C1 (n_5_84), .C2 (n_8_84) );
AOI211_X1 g_16_77 (.ZN (n_16_77), .A (n_15_76), .B (n_10_80), .C1 (n_7_83), .C2 (n_6_85) );
AOI211_X1 g_15_75 (.ZN (n_15_75), .A (n_17_75), .B (n_11_78), .C1 (n_9_82), .C2 (n_4_86) );
AOI211_X1 g_17_74 (.ZN (n_17_74), .A (n_16_77), .B (n_13_77), .C1 (n_10_80), .C2 (n_5_84) );
AOI211_X1 g_19_73 (.ZN (n_19_73), .A (n_15_75), .B (n_15_76), .C1 (n_11_78), .C2 (n_7_83) );
AOI211_X1 g_20_75 (.ZN (n_20_75), .A (n_17_74), .B (n_17_75), .C1 (n_13_77), .C2 (n_9_82) );
AOI211_X1 g_18_76 (.ZN (n_18_76), .A (n_19_73), .B (n_16_77), .C1 (n_15_76), .C2 (n_10_80) );
AOI211_X1 g_17_78 (.ZN (n_17_78), .A (n_20_75), .B (n_15_75), .C1 (n_17_75), .C2 (n_11_78) );
AOI211_X1 g_16_76 (.ZN (n_16_76), .A (n_18_76), .B (n_17_74), .C1 (n_16_77), .C2 (n_13_77) );
AOI211_X1 g_18_75 (.ZN (n_18_75), .A (n_17_78), .B (n_19_73), .C1 (n_15_75), .C2 (n_15_76) );
AOI211_X1 g_20_74 (.ZN (n_20_74), .A (n_16_76), .B (n_20_75), .C1 (n_17_74), .C2 (n_17_75) );
AOI211_X1 g_22_73 (.ZN (n_22_73), .A (n_18_75), .B (n_18_76), .C1 (n_19_73), .C2 (n_16_77) );
AOI211_X1 g_24_72 (.ZN (n_24_72), .A (n_20_74), .B (n_17_78), .C1 (n_20_75), .C2 (n_15_75) );
AOI211_X1 g_26_71 (.ZN (n_26_71), .A (n_22_73), .B (n_16_76), .C1 (n_18_76), .C2 (n_17_74) );
AOI211_X1 g_28_70 (.ZN (n_28_70), .A (n_24_72), .B (n_18_75), .C1 (n_17_78), .C2 (n_19_73) );
AOI211_X1 g_30_69 (.ZN (n_30_69), .A (n_26_71), .B (n_20_74), .C1 (n_16_76), .C2 (n_20_75) );
AOI211_X1 g_32_68 (.ZN (n_32_68), .A (n_28_70), .B (n_22_73), .C1 (n_18_75), .C2 (n_18_76) );
AOI211_X1 g_34_67 (.ZN (n_34_67), .A (n_30_69), .B (n_24_72), .C1 (n_20_74), .C2 (n_17_78) );
AOI211_X1 g_36_66 (.ZN (n_36_66), .A (n_32_68), .B (n_26_71), .C1 (n_22_73), .C2 (n_16_76) );
AOI211_X1 g_38_65 (.ZN (n_38_65), .A (n_34_67), .B (n_28_70), .C1 (n_24_72), .C2 (n_18_75) );
AOI211_X1 g_40_64 (.ZN (n_40_64), .A (n_36_66), .B (n_30_69), .C1 (n_26_71), .C2 (n_20_74) );
AOI211_X1 g_42_63 (.ZN (n_42_63), .A (n_38_65), .B (n_32_68), .C1 (n_28_70), .C2 (n_22_73) );
AOI211_X1 g_44_62 (.ZN (n_44_62), .A (n_40_64), .B (n_34_67), .C1 (n_30_69), .C2 (n_24_72) );
AOI211_X1 g_46_61 (.ZN (n_46_61), .A (n_42_63), .B (n_36_66), .C1 (n_32_68), .C2 (n_26_71) );
AOI211_X1 g_48_60 (.ZN (n_48_60), .A (n_44_62), .B (n_38_65), .C1 (n_34_67), .C2 (n_28_70) );
AOI211_X1 g_50_59 (.ZN (n_50_59), .A (n_46_61), .B (n_40_64), .C1 (n_36_66), .C2 (n_30_69) );
AOI211_X1 g_52_58 (.ZN (n_52_58), .A (n_48_60), .B (n_42_63), .C1 (n_38_65), .C2 (n_32_68) );
AOI211_X1 g_54_57 (.ZN (n_54_57), .A (n_50_59), .B (n_44_62), .C1 (n_40_64), .C2 (n_34_67) );
AOI211_X1 g_56_56 (.ZN (n_56_56), .A (n_52_58), .B (n_46_61), .C1 (n_42_63), .C2 (n_36_66) );
AOI211_X1 g_58_55 (.ZN (n_58_55), .A (n_54_57), .B (n_48_60), .C1 (n_44_62), .C2 (n_38_65) );
AOI211_X1 g_60_54 (.ZN (n_60_54), .A (n_56_56), .B (n_50_59), .C1 (n_46_61), .C2 (n_40_64) );
AOI211_X1 g_62_53 (.ZN (n_62_53), .A (n_58_55), .B (n_52_58), .C1 (n_48_60), .C2 (n_42_63) );
AOI211_X1 g_64_52 (.ZN (n_64_52), .A (n_60_54), .B (n_54_57), .C1 (n_50_59), .C2 (n_44_62) );
AOI211_X1 g_66_51 (.ZN (n_66_51), .A (n_62_53), .B (n_56_56), .C1 (n_52_58), .C2 (n_46_61) );
AOI211_X1 g_68_50 (.ZN (n_68_50), .A (n_64_52), .B (n_58_55), .C1 (n_54_57), .C2 (n_48_60) );
AOI211_X1 g_70_51 (.ZN (n_70_51), .A (n_66_51), .B (n_60_54), .C1 (n_56_56), .C2 (n_50_59) );
AOI211_X1 g_68_52 (.ZN (n_68_52), .A (n_68_50), .B (n_62_53), .C1 (n_58_55), .C2 (n_52_58) );
AOI211_X1 g_69_50 (.ZN (n_69_50), .A (n_70_51), .B (n_64_52), .C1 (n_60_54), .C2 (n_54_57) );
AOI211_X1 g_67_51 (.ZN (n_67_51), .A (n_68_52), .B (n_66_51), .C1 (n_62_53), .C2 (n_56_56) );
AOI211_X1 g_65_52 (.ZN (n_65_52), .A (n_69_50), .B (n_68_50), .C1 (n_64_52), .C2 (n_58_55) );
AOI211_X1 g_63_53 (.ZN (n_63_53), .A (n_67_51), .B (n_70_51), .C1 (n_66_51), .C2 (n_60_54) );
AOI211_X1 g_61_54 (.ZN (n_61_54), .A (n_65_52), .B (n_68_52), .C1 (n_68_50), .C2 (n_62_53) );
AOI211_X1 g_59_55 (.ZN (n_59_55), .A (n_63_53), .B (n_69_50), .C1 (n_70_51), .C2 (n_64_52) );
AOI211_X1 g_58_57 (.ZN (n_58_57), .A (n_61_54), .B (n_67_51), .C1 (n_68_52), .C2 (n_66_51) );
AOI211_X1 g_60_56 (.ZN (n_60_56), .A (n_59_55), .B (n_65_52), .C1 (n_69_50), .C2 (n_68_50) );
AOI211_X1 g_62_55 (.ZN (n_62_55), .A (n_58_57), .B (n_63_53), .C1 (n_67_51), .C2 (n_70_51) );
AOI211_X1 g_64_54 (.ZN (n_64_54), .A (n_60_56), .B (n_61_54), .C1 (n_65_52), .C2 (n_68_52) );
AOI211_X1 g_66_53 (.ZN (n_66_53), .A (n_62_55), .B (n_59_55), .C1 (n_63_53), .C2 (n_69_50) );
AOI211_X1 g_65_55 (.ZN (n_65_55), .A (n_64_54), .B (n_58_57), .C1 (n_61_54), .C2 (n_67_51) );
AOI211_X1 g_63_54 (.ZN (n_63_54), .A (n_66_53), .B (n_60_56), .C1 (n_59_55), .C2 (n_65_52) );
AOI211_X1 g_65_53 (.ZN (n_65_53), .A (n_65_55), .B (n_62_55), .C1 (n_58_57), .C2 (n_63_53) );
AOI211_X1 g_67_52 (.ZN (n_67_52), .A (n_63_54), .B (n_64_54), .C1 (n_60_56), .C2 (n_61_54) );
AOI211_X1 g_69_51 (.ZN (n_69_51), .A (n_65_53), .B (n_66_53), .C1 (n_62_55), .C2 (n_59_55) );
AOI211_X1 g_71_50 (.ZN (n_71_50), .A (n_67_52), .B (n_65_55), .C1 (n_64_54), .C2 (n_58_57) );
AOI211_X1 g_73_49 (.ZN (n_73_49), .A (n_69_51), .B (n_63_54), .C1 (n_66_53), .C2 (n_60_56) );
AOI211_X1 g_75_48 (.ZN (n_75_48), .A (n_71_50), .B (n_65_53), .C1 (n_65_55), .C2 (n_62_55) );
AOI211_X1 g_77_47 (.ZN (n_77_47), .A (n_73_49), .B (n_67_52), .C1 (n_63_54), .C2 (n_64_54) );
AOI211_X1 g_79_46 (.ZN (n_79_46), .A (n_75_48), .B (n_69_51), .C1 (n_65_53), .C2 (n_66_53) );
AOI211_X1 g_81_45 (.ZN (n_81_45), .A (n_77_47), .B (n_71_50), .C1 (n_67_52), .C2 (n_65_55) );
AOI211_X1 g_83_44 (.ZN (n_83_44), .A (n_79_46), .B (n_73_49), .C1 (n_69_51), .C2 (n_63_54) );
AOI211_X1 g_85_43 (.ZN (n_85_43), .A (n_81_45), .B (n_75_48), .C1 (n_71_50), .C2 (n_65_53) );
AOI211_X1 g_87_42 (.ZN (n_87_42), .A (n_83_44), .B (n_77_47), .C1 (n_73_49), .C2 (n_67_52) );
AOI211_X1 g_89_41 (.ZN (n_89_41), .A (n_85_43), .B (n_79_46), .C1 (n_75_48), .C2 (n_69_51) );
AOI211_X1 g_91_40 (.ZN (n_91_40), .A (n_87_42), .B (n_81_45), .C1 (n_77_47), .C2 (n_71_50) );
AOI211_X1 g_93_39 (.ZN (n_93_39), .A (n_89_41), .B (n_83_44), .C1 (n_79_46), .C2 (n_73_49) );
AOI211_X1 g_95_38 (.ZN (n_95_38), .A (n_91_40), .B (n_85_43), .C1 (n_81_45), .C2 (n_75_48) );
AOI211_X1 g_97_37 (.ZN (n_97_37), .A (n_93_39), .B (n_87_42), .C1 (n_83_44), .C2 (n_77_47) );
AOI211_X1 g_98_39 (.ZN (n_98_39), .A (n_95_38), .B (n_89_41), .C1 (n_85_43), .C2 (n_79_46) );
AOI211_X1 g_100_40 (.ZN (n_100_40), .A (n_97_37), .B (n_91_40), .C1 (n_87_42), .C2 (n_81_45) );
AOI211_X1 g_99_38 (.ZN (n_99_38), .A (n_98_39), .B (n_93_39), .C1 (n_89_41), .C2 (n_83_44) );
AOI211_X1 g_97_39 (.ZN (n_97_39), .A (n_100_40), .B (n_95_38), .C1 (n_91_40), .C2 (n_85_43) );
AOI211_X1 g_95_40 (.ZN (n_95_40), .A (n_99_38), .B (n_97_37), .C1 (n_93_39), .C2 (n_87_42) );
AOI211_X1 g_93_41 (.ZN (n_93_41), .A (n_97_39), .B (n_98_39), .C1 (n_95_38), .C2 (n_89_41) );
AOI211_X1 g_91_42 (.ZN (n_91_42), .A (n_95_40), .B (n_100_40), .C1 (n_97_37), .C2 (n_91_40) );
AOI211_X1 g_89_43 (.ZN (n_89_43), .A (n_93_41), .B (n_99_38), .C1 (n_98_39), .C2 (n_93_39) );
AOI211_X1 g_87_44 (.ZN (n_87_44), .A (n_91_42), .B (n_97_39), .C1 (n_100_40), .C2 (n_95_38) );
AOI211_X1 g_86_46 (.ZN (n_86_46), .A (n_89_43), .B (n_95_40), .C1 (n_99_38), .C2 (n_97_37) );
AOI211_X1 g_85_44 (.ZN (n_85_44), .A (n_87_44), .B (n_93_41), .C1 (n_97_39), .C2 (n_98_39) );
AOI211_X1 g_87_43 (.ZN (n_87_43), .A (n_86_46), .B (n_91_42), .C1 (n_95_40), .C2 (n_100_40) );
AOI211_X1 g_89_42 (.ZN (n_89_42), .A (n_85_44), .B (n_89_43), .C1 (n_93_41), .C2 (n_99_38) );
AOI211_X1 g_91_41 (.ZN (n_91_41), .A (n_87_43), .B (n_87_44), .C1 (n_91_42), .C2 (n_97_39) );
AOI211_X1 g_90_43 (.ZN (n_90_43), .A (n_89_42), .B (n_86_46), .C1 (n_89_43), .C2 (n_95_40) );
AOI211_X1 g_92_42 (.ZN (n_92_42), .A (n_91_41), .B (n_85_44), .C1 (n_87_44), .C2 (n_93_41) );
AOI211_X1 g_94_41 (.ZN (n_94_41), .A (n_90_43), .B (n_87_43), .C1 (n_86_46), .C2 (n_91_42) );
AOI211_X1 g_96_40 (.ZN (n_96_40), .A (n_92_42), .B (n_89_42), .C1 (n_85_44), .C2 (n_89_43) );
AOI211_X1 g_98_41 (.ZN (n_98_41), .A (n_94_41), .B (n_91_41), .C1 (n_87_43), .C2 (n_87_44) );
AOI211_X1 g_96_42 (.ZN (n_96_42), .A (n_96_40), .B (n_90_43), .C1 (n_89_42), .C2 (n_86_46) );
AOI211_X1 g_94_43 (.ZN (n_94_43), .A (n_98_41), .B (n_92_42), .C1 (n_91_41), .C2 (n_85_44) );
AOI211_X1 g_95_41 (.ZN (n_95_41), .A (n_96_42), .B (n_94_41), .C1 (n_90_43), .C2 (n_87_43) );
AOI211_X1 g_96_39 (.ZN (n_96_39), .A (n_94_43), .B (n_96_40), .C1 (n_92_42), .C2 (n_89_42) );
AOI211_X1 g_98_40 (.ZN (n_98_40), .A (n_95_41), .B (n_98_41), .C1 (n_94_41), .C2 (n_91_41) );
AOI211_X1 g_96_41 (.ZN (n_96_41), .A (n_96_39), .B (n_96_42), .C1 (n_96_40), .C2 (n_90_43) );
AOI211_X1 g_94_40 (.ZN (n_94_40), .A (n_98_40), .B (n_94_43), .C1 (n_98_41), .C2 (n_92_42) );
AOI211_X1 g_92_41 (.ZN (n_92_41), .A (n_96_41), .B (n_95_41), .C1 (n_96_42), .C2 (n_94_41) );
AOI211_X1 g_90_42 (.ZN (n_90_42), .A (n_94_40), .B (n_96_39), .C1 (n_94_43), .C2 (n_96_40) );
AOI211_X1 g_88_43 (.ZN (n_88_43), .A (n_92_41), .B (n_98_40), .C1 (n_95_41), .C2 (n_98_41) );
AOI211_X1 g_86_44 (.ZN (n_86_44), .A (n_90_42), .B (n_96_41), .C1 (n_96_39), .C2 (n_96_42) );
AOI211_X1 g_84_45 (.ZN (n_84_45), .A (n_88_43), .B (n_94_40), .C1 (n_98_40), .C2 (n_94_43) );
AOI211_X1 g_82_46 (.ZN (n_82_46), .A (n_86_44), .B (n_92_41), .C1 (n_96_41), .C2 (n_95_41) );
AOI211_X1 g_80_47 (.ZN (n_80_47), .A (n_84_45), .B (n_90_42), .C1 (n_94_40), .C2 (n_96_39) );
AOI211_X1 g_78_48 (.ZN (n_78_48), .A (n_82_46), .B (n_88_43), .C1 (n_92_41), .C2 (n_98_40) );
AOI211_X1 g_76_49 (.ZN (n_76_49), .A (n_80_47), .B (n_86_44), .C1 (n_90_42), .C2 (n_96_41) );
AOI211_X1 g_74_50 (.ZN (n_74_50), .A (n_78_48), .B (n_84_45), .C1 (n_88_43), .C2 (n_94_40) );
AOI211_X1 g_72_51 (.ZN (n_72_51), .A (n_76_49), .B (n_82_46), .C1 (n_86_44), .C2 (n_92_41) );
AOI211_X1 g_70_52 (.ZN (n_70_52), .A (n_74_50), .B (n_80_47), .C1 (n_84_45), .C2 (n_90_42) );
AOI211_X1 g_68_53 (.ZN (n_68_53), .A (n_72_51), .B (n_78_48), .C1 (n_82_46), .C2 (n_88_43) );
AOI211_X1 g_66_54 (.ZN (n_66_54), .A (n_70_52), .B (n_76_49), .C1 (n_80_47), .C2 (n_86_44) );
AOI211_X1 g_64_55 (.ZN (n_64_55), .A (n_68_53), .B (n_74_50), .C1 (n_78_48), .C2 (n_84_45) );
AOI211_X1 g_62_56 (.ZN (n_62_56), .A (n_66_54), .B (n_72_51), .C1 (n_76_49), .C2 (n_82_46) );
AOI211_X1 g_60_57 (.ZN (n_60_57), .A (n_64_55), .B (n_70_52), .C1 (n_74_50), .C2 (n_80_47) );
AOI211_X1 g_61_55 (.ZN (n_61_55), .A (n_62_56), .B (n_68_53), .C1 (n_72_51), .C2 (n_78_48) );
AOI211_X1 g_59_56 (.ZN (n_59_56), .A (n_60_57), .B (n_66_54), .C1 (n_70_52), .C2 (n_76_49) );
AOI211_X1 g_57_57 (.ZN (n_57_57), .A (n_61_55), .B (n_64_55), .C1 (n_68_53), .C2 (n_74_50) );
AOI211_X1 g_55_58 (.ZN (n_55_58), .A (n_59_56), .B (n_62_56), .C1 (n_66_54), .C2 (n_72_51) );
AOI211_X1 g_53_59 (.ZN (n_53_59), .A (n_57_57), .B (n_60_57), .C1 (n_64_55), .C2 (n_70_52) );
AOI211_X1 g_51_60 (.ZN (n_51_60), .A (n_55_58), .B (n_61_55), .C1 (n_62_56), .C2 (n_68_53) );
AOI211_X1 g_49_61 (.ZN (n_49_61), .A (n_53_59), .B (n_59_56), .C1 (n_60_57), .C2 (n_66_54) );
AOI211_X1 g_47_62 (.ZN (n_47_62), .A (n_51_60), .B (n_57_57), .C1 (n_61_55), .C2 (n_64_55) );
AOI211_X1 g_45_63 (.ZN (n_45_63), .A (n_49_61), .B (n_55_58), .C1 (n_59_56), .C2 (n_62_56) );
AOI211_X1 g_43_64 (.ZN (n_43_64), .A (n_47_62), .B (n_53_59), .C1 (n_57_57), .C2 (n_60_57) );
AOI211_X1 g_41_65 (.ZN (n_41_65), .A (n_45_63), .B (n_51_60), .C1 (n_55_58), .C2 (n_61_55) );
AOI211_X1 g_39_66 (.ZN (n_39_66), .A (n_43_64), .B (n_49_61), .C1 (n_53_59), .C2 (n_59_56) );
AOI211_X1 g_37_67 (.ZN (n_37_67), .A (n_41_65), .B (n_47_62), .C1 (n_51_60), .C2 (n_57_57) );
AOI211_X1 g_35_68 (.ZN (n_35_68), .A (n_39_66), .B (n_45_63), .C1 (n_49_61), .C2 (n_55_58) );
AOI211_X1 g_33_69 (.ZN (n_33_69), .A (n_37_67), .B (n_43_64), .C1 (n_47_62), .C2 (n_53_59) );
AOI211_X1 g_31_70 (.ZN (n_31_70), .A (n_35_68), .B (n_41_65), .C1 (n_45_63), .C2 (n_51_60) );
AOI211_X1 g_29_71 (.ZN (n_29_71), .A (n_33_69), .B (n_39_66), .C1 (n_43_64), .C2 (n_49_61) );
AOI211_X1 g_27_72 (.ZN (n_27_72), .A (n_31_70), .B (n_37_67), .C1 (n_41_65), .C2 (n_47_62) );
AOI211_X1 g_25_73 (.ZN (n_25_73), .A (n_29_71), .B (n_35_68), .C1 (n_39_66), .C2 (n_45_63) );
AOI211_X1 g_23_74 (.ZN (n_23_74), .A (n_27_72), .B (n_33_69), .C1 (n_37_67), .C2 (n_43_64) );
AOI211_X1 g_21_75 (.ZN (n_21_75), .A (n_25_73), .B (n_31_70), .C1 (n_35_68), .C2 (n_41_65) );
AOI211_X1 g_19_76 (.ZN (n_19_76), .A (n_23_74), .B (n_29_71), .C1 (n_33_69), .C2 (n_39_66) );
AOI211_X1 g_17_77 (.ZN (n_17_77), .A (n_21_75), .B (n_27_72), .C1 (n_31_70), .C2 (n_37_67) );
AOI211_X1 g_15_78 (.ZN (n_15_78), .A (n_19_76), .B (n_25_73), .C1 (n_29_71), .C2 (n_35_68) );
AOI211_X1 g_13_79 (.ZN (n_13_79), .A (n_17_77), .B (n_23_74), .C1 (n_27_72), .C2 (n_33_69) );
AOI211_X1 g_14_77 (.ZN (n_14_77), .A (n_15_78), .B (n_21_75), .C1 (n_25_73), .C2 (n_31_70) );
AOI211_X1 g_12_78 (.ZN (n_12_78), .A (n_13_79), .B (n_19_76), .C1 (n_23_74), .C2 (n_29_71) );
AOI211_X1 g_13_76 (.ZN (n_13_76), .A (n_14_77), .B (n_17_77), .C1 (n_21_75), .C2 (n_27_72) );
AOI211_X1 g_11_77 (.ZN (n_11_77), .A (n_12_78), .B (n_15_78), .C1 (n_19_76), .C2 (n_25_73) );
AOI211_X1 g_10_79 (.ZN (n_10_79), .A (n_13_76), .B (n_13_79), .C1 (n_17_77), .C2 (n_23_74) );
AOI211_X1 g_9_81 (.ZN (n_9_81), .A (n_11_77), .B (n_14_77), .C1 (n_15_78), .C2 (n_21_75) );
AOI211_X1 g_7_80 (.ZN (n_7_80), .A (n_10_79), .B (n_12_78), .C1 (n_13_79), .C2 (n_19_76) );
AOI211_X1 g_9_79 (.ZN (n_9_79), .A (n_9_81), .B (n_13_76), .C1 (n_14_77), .C2 (n_17_77) );
AOI211_X1 g_8_81 (.ZN (n_8_81), .A (n_7_80), .B (n_11_77), .C1 (n_12_78), .C2 (n_15_78) );
AOI211_X1 g_6_82 (.ZN (n_6_82), .A (n_9_79), .B (n_10_79), .C1 (n_13_76), .C2 (n_13_79) );
AOI211_X1 g_8_83 (.ZN (n_8_83), .A (n_8_81), .B (n_9_81), .C1 (n_11_77), .C2 (n_14_77) );
AOI211_X1 g_7_85 (.ZN (n_7_85), .A (n_6_82), .B (n_7_80), .C1 (n_10_79), .C2 (n_12_78) );
AOI211_X1 g_6_87 (.ZN (n_6_87), .A (n_8_83), .B (n_9_79), .C1 (n_9_81), .C2 (n_13_76) );
AOI211_X1 g_5_89 (.ZN (n_5_89), .A (n_7_85), .B (n_8_81), .C1 (n_7_80), .C2 (n_11_77) );
AOI211_X1 g_4_91 (.ZN (n_4_91), .A (n_6_87), .B (n_6_82), .C1 (n_9_79), .C2 (n_10_79) );
AOI211_X1 g_6_92 (.ZN (n_6_92), .A (n_5_89), .B (n_8_83), .C1 (n_8_81), .C2 (n_9_81) );
AOI211_X1 g_7_90 (.ZN (n_7_90), .A (n_4_91), .B (n_7_85), .C1 (n_6_82), .C2 (n_7_80) );
AOI211_X1 g_8_88 (.ZN (n_8_88), .A (n_6_92), .B (n_6_87), .C1 (n_8_83), .C2 (n_9_79) );
AOI211_X1 g_9_86 (.ZN (n_9_86), .A (n_7_90), .B (n_5_89), .C1 (n_7_85), .C2 (n_8_81) );
AOI211_X1 g_10_84 (.ZN (n_10_84), .A (n_8_88), .B (n_4_91), .C1 (n_6_87), .C2 (n_6_82) );
AOI211_X1 g_11_82 (.ZN (n_11_82), .A (n_9_86), .B (n_6_92), .C1 (n_5_89), .C2 (n_8_83) );
AOI211_X1 g_12_80 (.ZN (n_12_80), .A (n_10_84), .B (n_7_90), .C1 (n_4_91), .C2 (n_7_85) );
AOI211_X1 g_13_78 (.ZN (n_13_78), .A (n_11_82), .B (n_8_88), .C1 (n_6_92), .C2 (n_6_87) );
AOI211_X1 g_15_77 (.ZN (n_15_77), .A (n_12_80), .B (n_9_86), .C1 (n_7_90), .C2 (n_5_89) );
AOI211_X1 g_17_76 (.ZN (n_17_76), .A (n_13_78), .B (n_10_84), .C1 (n_8_88), .C2 (n_4_91) );
AOI211_X1 g_19_75 (.ZN (n_19_75), .A (n_15_77), .B (n_11_82), .C1 (n_9_86), .C2 (n_6_92) );
AOI211_X1 g_21_74 (.ZN (n_21_74), .A (n_17_76), .B (n_12_80), .C1 (n_10_84), .C2 (n_7_90) );
AOI211_X1 g_23_73 (.ZN (n_23_73), .A (n_19_75), .B (n_13_78), .C1 (n_11_82), .C2 (n_8_88) );
AOI211_X1 g_25_72 (.ZN (n_25_72), .A (n_21_74), .B (n_15_77), .C1 (n_12_80), .C2 (n_9_86) );
AOI211_X1 g_27_71 (.ZN (n_27_71), .A (n_23_73), .B (n_17_76), .C1 (n_13_78), .C2 (n_10_84) );
AOI211_X1 g_29_70 (.ZN (n_29_70), .A (n_25_72), .B (n_19_75), .C1 (n_15_77), .C2 (n_11_82) );
AOI211_X1 g_31_69 (.ZN (n_31_69), .A (n_27_71), .B (n_21_74), .C1 (n_17_76), .C2 (n_12_80) );
AOI211_X1 g_33_68 (.ZN (n_33_68), .A (n_29_70), .B (n_23_73), .C1 (n_19_75), .C2 (n_13_78) );
AOI211_X1 g_35_67 (.ZN (n_35_67), .A (n_31_69), .B (n_25_72), .C1 (n_21_74), .C2 (n_15_77) );
AOI211_X1 g_37_66 (.ZN (n_37_66), .A (n_33_68), .B (n_27_71), .C1 (n_23_73), .C2 (n_17_76) );
AOI211_X1 g_39_65 (.ZN (n_39_65), .A (n_35_67), .B (n_29_70), .C1 (n_25_72), .C2 (n_19_75) );
AOI211_X1 g_38_67 (.ZN (n_38_67), .A (n_37_66), .B (n_31_69), .C1 (n_27_71), .C2 (n_21_74) );
AOI211_X1 g_40_66 (.ZN (n_40_66), .A (n_39_65), .B (n_33_68), .C1 (n_29_70), .C2 (n_23_73) );
AOI211_X1 g_42_65 (.ZN (n_42_65), .A (n_38_67), .B (n_35_67), .C1 (n_31_69), .C2 (n_25_72) );
AOI211_X1 g_44_64 (.ZN (n_44_64), .A (n_40_66), .B (n_37_66), .C1 (n_33_68), .C2 (n_27_71) );
AOI211_X1 g_46_63 (.ZN (n_46_63), .A (n_42_65), .B (n_39_65), .C1 (n_35_67), .C2 (n_29_70) );
AOI211_X1 g_48_62 (.ZN (n_48_62), .A (n_44_64), .B (n_38_67), .C1 (n_37_66), .C2 (n_31_69) );
AOI211_X1 g_50_61 (.ZN (n_50_61), .A (n_46_63), .B (n_40_66), .C1 (n_39_65), .C2 (n_33_68) );
AOI211_X1 g_52_60 (.ZN (n_52_60), .A (n_48_62), .B (n_42_65), .C1 (n_38_67), .C2 (n_35_67) );
AOI211_X1 g_54_59 (.ZN (n_54_59), .A (n_50_61), .B (n_44_64), .C1 (n_40_66), .C2 (n_37_66) );
AOI211_X1 g_56_58 (.ZN (n_56_58), .A (n_52_60), .B (n_46_63), .C1 (n_42_65), .C2 (n_39_65) );
AOI211_X1 g_55_60 (.ZN (n_55_60), .A (n_54_59), .B (n_48_62), .C1 (n_44_64), .C2 (n_38_67) );
AOI211_X1 g_54_58 (.ZN (n_54_58), .A (n_56_58), .B (n_50_61), .C1 (n_46_63), .C2 (n_40_66) );
AOI211_X1 g_56_57 (.ZN (n_56_57), .A (n_55_60), .B (n_52_60), .C1 (n_48_62), .C2 (n_42_65) );
AOI211_X1 g_58_56 (.ZN (n_58_56), .A (n_54_58), .B (n_54_59), .C1 (n_50_61), .C2 (n_44_64) );
AOI211_X1 g_57_58 (.ZN (n_57_58), .A (n_56_57), .B (n_56_58), .C1 (n_52_60), .C2 (n_46_63) );
AOI211_X1 g_59_57 (.ZN (n_59_57), .A (n_58_56), .B (n_55_60), .C1 (n_54_59), .C2 (n_48_62) );
AOI211_X1 g_61_56 (.ZN (n_61_56), .A (n_57_58), .B (n_54_58), .C1 (n_56_58), .C2 (n_50_61) );
AOI211_X1 g_63_55 (.ZN (n_63_55), .A (n_59_57), .B (n_56_57), .C1 (n_55_60), .C2 (n_52_60) );
AOI211_X1 g_65_54 (.ZN (n_65_54), .A (n_61_56), .B (n_58_56), .C1 (n_54_58), .C2 (n_54_59) );
AOI211_X1 g_67_53 (.ZN (n_67_53), .A (n_63_55), .B (n_57_58), .C1 (n_56_57), .C2 (n_56_58) );
AOI211_X1 g_69_52 (.ZN (n_69_52), .A (n_65_54), .B (n_59_57), .C1 (n_58_56), .C2 (n_55_60) );
AOI211_X1 g_71_51 (.ZN (n_71_51), .A (n_67_53), .B (n_61_56), .C1 (n_57_58), .C2 (n_54_58) );
AOI211_X1 g_73_50 (.ZN (n_73_50), .A (n_69_52), .B (n_63_55), .C1 (n_59_57), .C2 (n_56_57) );
AOI211_X1 g_75_49 (.ZN (n_75_49), .A (n_71_51), .B (n_65_54), .C1 (n_61_56), .C2 (n_58_56) );
AOI211_X1 g_77_48 (.ZN (n_77_48), .A (n_73_50), .B (n_67_53), .C1 (n_63_55), .C2 (n_57_58) );
AOI211_X1 g_79_47 (.ZN (n_79_47), .A (n_75_49), .B (n_69_52), .C1 (n_65_54), .C2 (n_59_57) );
AOI211_X1 g_81_46 (.ZN (n_81_46), .A (n_77_48), .B (n_71_51), .C1 (n_67_53), .C2 (n_61_56) );
AOI211_X1 g_83_45 (.ZN (n_83_45), .A (n_79_47), .B (n_73_50), .C1 (n_69_52), .C2 (n_63_55) );
AOI211_X1 g_84_47 (.ZN (n_84_47), .A (n_81_46), .B (n_75_49), .C1 (n_71_51), .C2 (n_65_54) );
AOI211_X1 g_82_48 (.ZN (n_82_48), .A (n_83_45), .B (n_77_48), .C1 (n_73_50), .C2 (n_67_53) );
AOI211_X1 g_83_46 (.ZN (n_83_46), .A (n_84_47), .B (n_79_47), .C1 (n_75_49), .C2 (n_69_52) );
AOI211_X1 g_81_47 (.ZN (n_81_47), .A (n_82_48), .B (n_81_46), .C1 (n_77_48), .C2 (n_71_51) );
AOI211_X1 g_79_48 (.ZN (n_79_48), .A (n_83_46), .B (n_83_45), .C1 (n_79_47), .C2 (n_73_50) );
AOI211_X1 g_77_49 (.ZN (n_77_49), .A (n_81_47), .B (n_84_47), .C1 (n_81_46), .C2 (n_75_49) );
AOI211_X1 g_78_47 (.ZN (n_78_47), .A (n_79_48), .B (n_82_48), .C1 (n_83_45), .C2 (n_77_48) );
AOI211_X1 g_76_48 (.ZN (n_76_48), .A (n_77_49), .B (n_83_46), .C1 (n_84_47), .C2 (n_79_47) );
AOI211_X1 g_74_49 (.ZN (n_74_49), .A (n_78_47), .B (n_81_47), .C1 (n_82_48), .C2 (n_81_46) );
AOI211_X1 g_73_51 (.ZN (n_73_51), .A (n_76_48), .B (n_79_48), .C1 (n_83_46), .C2 (n_83_45) );
AOI211_X1 g_75_50 (.ZN (n_75_50), .A (n_74_49), .B (n_77_49), .C1 (n_81_47), .C2 (n_84_47) );
AOI211_X1 g_74_52 (.ZN (n_74_52), .A (n_73_51), .B (n_78_47), .C1 (n_79_48), .C2 (n_82_48) );
AOI211_X1 g_76_51 (.ZN (n_76_51), .A (n_75_50), .B (n_76_48), .C1 (n_77_49), .C2 (n_83_46) );
AOI211_X1 g_78_50 (.ZN (n_78_50), .A (n_74_52), .B (n_74_49), .C1 (n_78_47), .C2 (n_81_47) );
AOI211_X1 g_80_49 (.ZN (n_80_49), .A (n_76_51), .B (n_73_51), .C1 (n_76_48), .C2 (n_79_48) );
AOI211_X1 g_79_51 (.ZN (n_79_51), .A (n_78_50), .B (n_75_50), .C1 (n_74_49), .C2 (n_77_49) );
AOI211_X1 g_78_49 (.ZN (n_78_49), .A (n_80_49), .B (n_74_52), .C1 (n_73_51), .C2 (n_78_47) );
AOI211_X1 g_80_48 (.ZN (n_80_48), .A (n_79_51), .B (n_76_51), .C1 (n_75_50), .C2 (n_76_48) );
AOI211_X1 g_82_47 (.ZN (n_82_47), .A (n_78_49), .B (n_78_50), .C1 (n_74_52), .C2 (n_74_49) );
AOI211_X1 g_84_46 (.ZN (n_84_46), .A (n_80_48), .B (n_80_49), .C1 (n_76_51), .C2 (n_73_51) );
AOI211_X1 g_86_45 (.ZN (n_86_45), .A (n_82_47), .B (n_79_51), .C1 (n_78_50), .C2 (n_75_50) );
AOI211_X1 g_88_44 (.ZN (n_88_44), .A (n_84_46), .B (n_78_49), .C1 (n_80_49), .C2 (n_74_52) );
AOI211_X1 g_87_46 (.ZN (n_87_46), .A (n_86_45), .B (n_80_48), .C1 (n_79_51), .C2 (n_76_51) );
AOI211_X1 g_89_45 (.ZN (n_89_45), .A (n_88_44), .B (n_82_47), .C1 (n_78_49), .C2 (n_78_50) );
AOI211_X1 g_91_44 (.ZN (n_91_44), .A (n_87_46), .B (n_84_46), .C1 (n_80_48), .C2 (n_80_49) );
AOI211_X1 g_93_43 (.ZN (n_93_43), .A (n_89_45), .B (n_86_45), .C1 (n_82_47), .C2 (n_79_51) );
AOI211_X1 g_95_42 (.ZN (n_95_42), .A (n_91_44), .B (n_88_44), .C1 (n_84_46), .C2 (n_78_49) );
AOI211_X1 g_97_41 (.ZN (n_97_41), .A (n_93_43), .B (n_87_46), .C1 (n_86_45), .C2 (n_80_48) );
AOI211_X1 g_99_42 (.ZN (n_99_42), .A (n_95_42), .B (n_89_45), .C1 (n_88_44), .C2 (n_82_47) );
AOI211_X1 g_97_43 (.ZN (n_97_43), .A (n_97_41), .B (n_91_44), .C1 (n_87_46), .C2 (n_84_46) );
AOI211_X1 g_95_44 (.ZN (n_95_44), .A (n_99_42), .B (n_93_43), .C1 (n_89_45), .C2 (n_86_45) );
AOI211_X1 g_94_42 (.ZN (n_94_42), .A (n_97_43), .B (n_95_42), .C1 (n_91_44), .C2 (n_88_44) );
AOI211_X1 g_92_43 (.ZN (n_92_43), .A (n_95_44), .B (n_97_41), .C1 (n_93_43), .C2 (n_87_46) );
AOI211_X1 g_90_44 (.ZN (n_90_44), .A (n_94_42), .B (n_99_42), .C1 (n_95_42), .C2 (n_89_45) );
AOI211_X1 g_88_45 (.ZN (n_88_45), .A (n_92_43), .B (n_97_43), .C1 (n_97_41), .C2 (n_91_44) );
AOI211_X1 g_87_47 (.ZN (n_87_47), .A (n_90_44), .B (n_95_44), .C1 (n_99_42), .C2 (n_93_43) );
AOI211_X1 g_85_46 (.ZN (n_85_46), .A (n_88_45), .B (n_94_42), .C1 (n_97_43), .C2 (n_95_42) );
AOI211_X1 g_87_45 (.ZN (n_87_45), .A (n_87_47), .B (n_92_43), .C1 (n_95_44), .C2 (n_97_41) );
AOI211_X1 g_89_44 (.ZN (n_89_44), .A (n_85_46), .B (n_90_44), .C1 (n_94_42), .C2 (n_99_42) );
AOI211_X1 g_91_43 (.ZN (n_91_43), .A (n_87_45), .B (n_88_45), .C1 (n_92_43), .C2 (n_97_43) );
AOI211_X1 g_93_42 (.ZN (n_93_42), .A (n_89_44), .B (n_87_47), .C1 (n_90_44), .C2 (n_95_44) );
AOI211_X1 g_92_44 (.ZN (n_92_44), .A (n_91_43), .B (n_85_46), .C1 (n_88_45), .C2 (n_94_42) );
AOI211_X1 g_90_45 (.ZN (n_90_45), .A (n_93_42), .B (n_87_45), .C1 (n_87_47), .C2 (n_92_43) );
AOI211_X1 g_88_46 (.ZN (n_88_46), .A (n_92_44), .B (n_89_44), .C1 (n_85_46), .C2 (n_90_44) );
AOI211_X1 g_86_47 (.ZN (n_86_47), .A (n_90_45), .B (n_91_43), .C1 (n_87_45), .C2 (n_88_45) );
AOI211_X1 g_84_48 (.ZN (n_84_48), .A (n_88_46), .B (n_93_42), .C1 (n_89_44), .C2 (n_87_47) );
AOI211_X1 g_82_49 (.ZN (n_82_49), .A (n_86_47), .B (n_92_44), .C1 (n_91_43), .C2 (n_85_46) );
AOI211_X1 g_83_47 (.ZN (n_83_47), .A (n_84_48), .B (n_90_45), .C1 (n_93_42), .C2 (n_87_45) );
AOI211_X1 g_81_48 (.ZN (n_81_48), .A (n_82_49), .B (n_88_46), .C1 (n_92_44), .C2 (n_89_44) );
AOI211_X1 g_79_49 (.ZN (n_79_49), .A (n_83_47), .B (n_86_47), .C1 (n_90_45), .C2 (n_91_43) );
AOI211_X1 g_77_50 (.ZN (n_77_50), .A (n_81_48), .B (n_84_48), .C1 (n_88_46), .C2 (n_93_42) );
AOI211_X1 g_75_51 (.ZN (n_75_51), .A (n_79_49), .B (n_82_49), .C1 (n_86_47), .C2 (n_92_44) );
AOI211_X1 g_73_52 (.ZN (n_73_52), .A (n_77_50), .B (n_83_47), .C1 (n_84_48), .C2 (n_90_45) );
AOI211_X1 g_71_53 (.ZN (n_71_53), .A (n_75_51), .B (n_81_48), .C1 (n_82_49), .C2 (n_88_46) );
AOI211_X1 g_69_54 (.ZN (n_69_54), .A (n_73_52), .B (n_79_49), .C1 (n_83_47), .C2 (n_86_47) );
AOI211_X1 g_67_55 (.ZN (n_67_55), .A (n_71_53), .B (n_77_50), .C1 (n_81_48), .C2 (n_84_48) );
AOI211_X1 g_65_56 (.ZN (n_65_56), .A (n_69_54), .B (n_75_51), .C1 (n_79_49), .C2 (n_82_49) );
AOI211_X1 g_63_57 (.ZN (n_63_57), .A (n_67_55), .B (n_73_52), .C1 (n_77_50), .C2 (n_83_47) );
AOI211_X1 g_61_58 (.ZN (n_61_58), .A (n_65_56), .B (n_71_53), .C1 (n_75_51), .C2 (n_81_48) );
AOI211_X1 g_59_59 (.ZN (n_59_59), .A (n_63_57), .B (n_69_54), .C1 (n_73_52), .C2 (n_79_49) );
AOI211_X1 g_57_60 (.ZN (n_57_60), .A (n_61_58), .B (n_67_55), .C1 (n_71_53), .C2 (n_77_50) );
AOI211_X1 g_58_58 (.ZN (n_58_58), .A (n_59_59), .B (n_65_56), .C1 (n_69_54), .C2 (n_75_51) );
AOI211_X1 g_56_59 (.ZN (n_56_59), .A (n_57_60), .B (n_63_57), .C1 (n_67_55), .C2 (n_73_52) );
AOI211_X1 g_54_60 (.ZN (n_54_60), .A (n_58_58), .B (n_61_58), .C1 (n_65_56), .C2 (n_71_53) );
AOI211_X1 g_52_59 (.ZN (n_52_59), .A (n_56_59), .B (n_59_59), .C1 (n_63_57), .C2 (n_69_54) );
AOI211_X1 g_50_60 (.ZN (n_50_60), .A (n_54_60), .B (n_57_60), .C1 (n_61_58), .C2 (n_67_55) );
AOI211_X1 g_48_61 (.ZN (n_48_61), .A (n_52_59), .B (n_58_58), .C1 (n_59_59), .C2 (n_65_56) );
AOI211_X1 g_46_62 (.ZN (n_46_62), .A (n_50_60), .B (n_56_59), .C1 (n_57_60), .C2 (n_63_57) );
AOI211_X1 g_44_63 (.ZN (n_44_63), .A (n_48_61), .B (n_54_60), .C1 (n_58_58), .C2 (n_61_58) );
AOI211_X1 g_42_64 (.ZN (n_42_64), .A (n_46_62), .B (n_52_59), .C1 (n_56_59), .C2 (n_59_59) );
AOI211_X1 g_40_65 (.ZN (n_40_65), .A (n_44_63), .B (n_50_60), .C1 (n_54_60), .C2 (n_57_60) );
AOI211_X1 g_39_67 (.ZN (n_39_67), .A (n_42_64), .B (n_48_61), .C1 (n_52_59), .C2 (n_58_58) );
AOI211_X1 g_41_66 (.ZN (n_41_66), .A (n_40_65), .B (n_46_62), .C1 (n_50_60), .C2 (n_56_59) );
AOI211_X1 g_43_65 (.ZN (n_43_65), .A (n_39_67), .B (n_44_63), .C1 (n_48_61), .C2 (n_54_60) );
AOI211_X1 g_45_64 (.ZN (n_45_64), .A (n_41_66), .B (n_42_64), .C1 (n_46_62), .C2 (n_52_59) );
AOI211_X1 g_47_63 (.ZN (n_47_63), .A (n_43_65), .B (n_40_65), .C1 (n_44_63), .C2 (n_50_60) );
AOI211_X1 g_49_62 (.ZN (n_49_62), .A (n_45_64), .B (n_39_67), .C1 (n_42_64), .C2 (n_48_61) );
AOI211_X1 g_51_61 (.ZN (n_51_61), .A (n_47_63), .B (n_41_66), .C1 (n_40_65), .C2 (n_46_62) );
AOI211_X1 g_53_60 (.ZN (n_53_60), .A (n_49_62), .B (n_43_65), .C1 (n_39_67), .C2 (n_44_63) );
AOI211_X1 g_55_59 (.ZN (n_55_59), .A (n_51_61), .B (n_45_64), .C1 (n_41_66), .C2 (n_42_64) );
AOI211_X1 g_54_61 (.ZN (n_54_61), .A (n_53_60), .B (n_47_63), .C1 (n_43_65), .C2 (n_40_65) );
AOI211_X1 g_56_60 (.ZN (n_56_60), .A (n_55_59), .B (n_49_62), .C1 (n_45_64), .C2 (n_39_67) );
AOI211_X1 g_58_59 (.ZN (n_58_59), .A (n_54_61), .B (n_51_61), .C1 (n_47_63), .C2 (n_41_66) );
AOI211_X1 g_60_58 (.ZN (n_60_58), .A (n_56_60), .B (n_53_60), .C1 (n_49_62), .C2 (n_43_65) );
AOI211_X1 g_62_57 (.ZN (n_62_57), .A (n_58_59), .B (n_55_59), .C1 (n_51_61), .C2 (n_45_64) );
AOI211_X1 g_64_56 (.ZN (n_64_56), .A (n_60_58), .B (n_54_61), .C1 (n_53_60), .C2 (n_47_63) );
AOI211_X1 g_66_55 (.ZN (n_66_55), .A (n_62_57), .B (n_56_60), .C1 (n_55_59), .C2 (n_49_62) );
AOI211_X1 g_68_54 (.ZN (n_68_54), .A (n_64_56), .B (n_58_59), .C1 (n_54_61), .C2 (n_51_61) );
AOI211_X1 g_70_53 (.ZN (n_70_53), .A (n_66_55), .B (n_60_58), .C1 (n_56_60), .C2 (n_53_60) );
AOI211_X1 g_72_52 (.ZN (n_72_52), .A (n_68_54), .B (n_62_57), .C1 (n_58_59), .C2 (n_55_59) );
AOI211_X1 g_74_51 (.ZN (n_74_51), .A (n_70_53), .B (n_64_56), .C1 (n_60_58), .C2 (n_54_61) );
AOI211_X1 g_76_50 (.ZN (n_76_50), .A (n_72_52), .B (n_66_55), .C1 (n_62_57), .C2 (n_56_60) );
AOI211_X1 g_77_52 (.ZN (n_77_52), .A (n_74_51), .B (n_68_54), .C1 (n_64_56), .C2 (n_58_59) );
AOI211_X1 g_75_53 (.ZN (n_75_53), .A (n_76_50), .B (n_70_53), .C1 (n_66_55), .C2 (n_60_58) );
AOI211_X1 g_73_54 (.ZN (n_73_54), .A (n_77_52), .B (n_72_52), .C1 (n_68_54), .C2 (n_62_57) );
AOI211_X1 g_71_55 (.ZN (n_71_55), .A (n_75_53), .B (n_74_51), .C1 (n_70_53), .C2 (n_64_56) );
AOI211_X1 g_72_53 (.ZN (n_72_53), .A (n_73_54), .B (n_76_50), .C1 (n_72_52), .C2 (n_66_55) );
AOI211_X1 g_70_54 (.ZN (n_70_54), .A (n_71_55), .B (n_77_52), .C1 (n_74_51), .C2 (n_68_54) );
AOI211_X1 g_71_52 (.ZN (n_71_52), .A (n_72_53), .B (n_75_53), .C1 (n_76_50), .C2 (n_70_53) );
AOI211_X1 g_69_53 (.ZN (n_69_53), .A (n_70_54), .B (n_73_54), .C1 (n_77_52), .C2 (n_72_52) );
AOI211_X1 g_67_54 (.ZN (n_67_54), .A (n_71_52), .B (n_71_55), .C1 (n_75_53), .C2 (n_74_51) );
AOI211_X1 g_66_56 (.ZN (n_66_56), .A (n_69_53), .B (n_72_53), .C1 (n_73_54), .C2 (n_76_50) );
AOI211_X1 g_68_55 (.ZN (n_68_55), .A (n_67_54), .B (n_70_54), .C1 (n_71_55), .C2 (n_77_52) );
AOI211_X1 g_67_57 (.ZN (n_67_57), .A (n_66_56), .B (n_71_52), .C1 (n_72_53), .C2 (n_75_53) );
AOI211_X1 g_69_56 (.ZN (n_69_56), .A (n_68_55), .B (n_69_53), .C1 (n_70_54), .C2 (n_73_54) );
AOI211_X1 g_68_58 (.ZN (n_68_58), .A (n_67_57), .B (n_67_54), .C1 (n_71_52), .C2 (n_71_55) );
AOI211_X1 g_67_56 (.ZN (n_67_56), .A (n_69_56), .B (n_66_56), .C1 (n_69_53), .C2 (n_72_53) );
AOI211_X1 g_69_55 (.ZN (n_69_55), .A (n_68_58), .B (n_68_55), .C1 (n_67_54), .C2 (n_70_54) );
AOI211_X1 g_71_54 (.ZN (n_71_54), .A (n_67_56), .B (n_67_57), .C1 (n_66_56), .C2 (n_71_52) );
AOI211_X1 g_73_53 (.ZN (n_73_53), .A (n_69_55), .B (n_69_56), .C1 (n_68_55), .C2 (n_69_53) );
AOI211_X1 g_75_52 (.ZN (n_75_52), .A (n_71_54), .B (n_68_58), .C1 (n_67_57), .C2 (n_67_54) );
AOI211_X1 g_77_51 (.ZN (n_77_51), .A (n_73_53), .B (n_67_56), .C1 (n_69_56), .C2 (n_66_56) );
AOI211_X1 g_79_50 (.ZN (n_79_50), .A (n_75_52), .B (n_69_55), .C1 (n_68_58), .C2 (n_68_55) );
AOI211_X1 g_81_49 (.ZN (n_81_49), .A (n_77_51), .B (n_71_54), .C1 (n_67_56), .C2 (n_67_57) );
AOI211_X1 g_83_48 (.ZN (n_83_48), .A (n_79_50), .B (n_73_53), .C1 (n_69_55), .C2 (n_69_56) );
AOI211_X1 g_85_47 (.ZN (n_85_47), .A (n_81_49), .B (n_75_52), .C1 (n_71_54), .C2 (n_68_58) );
AOI211_X1 g_84_49 (.ZN (n_84_49), .A (n_83_48), .B (n_77_51), .C1 (n_73_53), .C2 (n_67_56) );
AOI211_X1 g_86_48 (.ZN (n_86_48), .A (n_85_47), .B (n_79_50), .C1 (n_75_52), .C2 (n_69_55) );
AOI211_X1 g_88_47 (.ZN (n_88_47), .A (n_84_49), .B (n_81_49), .C1 (n_77_51), .C2 (n_71_54) );
AOI211_X1 g_90_46 (.ZN (n_90_46), .A (n_86_48), .B (n_83_48), .C1 (n_79_50), .C2 (n_73_53) );
AOI211_X1 g_92_45 (.ZN (n_92_45), .A (n_88_47), .B (n_85_47), .C1 (n_81_49), .C2 (n_75_52) );
AOI211_X1 g_94_44 (.ZN (n_94_44), .A (n_90_46), .B (n_84_49), .C1 (n_83_48), .C2 (n_77_51) );
AOI211_X1 g_96_43 (.ZN (n_96_43), .A (n_92_45), .B (n_86_48), .C1 (n_85_47), .C2 (n_79_50) );
AOI211_X1 g_97_45 (.ZN (n_97_45), .A (n_94_44), .B (n_88_47), .C1 (n_84_49), .C2 (n_81_49) );
AOI211_X1 g_98_43 (.ZN (n_98_43), .A (n_96_43), .B (n_90_46), .C1 (n_86_48), .C2 (n_83_48) );
AOI211_X1 g_100_44 (.ZN (n_100_44), .A (n_97_45), .B (n_92_45), .C1 (n_88_47), .C2 (n_85_47) );
AOI211_X1 g_99_46 (.ZN (n_99_46), .A (n_98_43), .B (n_94_44), .C1 (n_90_46), .C2 (n_84_49) );
AOI211_X1 g_100_48 (.ZN (n_100_48), .A (n_100_44), .B (n_96_43), .C1 (n_92_45), .C2 (n_86_48) );
AOI211_X1 g_98_47 (.ZN (n_98_47), .A (n_99_46), .B (n_97_45), .C1 (n_94_44), .C2 (n_88_47) );
AOI211_X1 g_99_45 (.ZN (n_99_45), .A (n_100_48), .B (n_98_43), .C1 (n_96_43), .C2 (n_90_46) );
AOI211_X1 g_100_47 (.ZN (n_100_47), .A (n_98_47), .B (n_100_44), .C1 (n_97_45), .C2 (n_92_45) );
AOI211_X1 g_99_49 (.ZN (n_99_49), .A (n_99_45), .B (n_99_46), .C1 (n_98_43), .C2 (n_94_44) );
AOI211_X1 g_100_51 (.ZN (n_100_51), .A (n_100_47), .B (n_100_48), .C1 (n_100_44), .C2 (n_96_43) );
AOI211_X1 g_98_50 (.ZN (n_98_50), .A (n_99_49), .B (n_98_47), .C1 (n_99_46), .C2 (n_97_45) );
AOI211_X1 g_100_49 (.ZN (n_100_49), .A (n_100_51), .B (n_99_45), .C1 (n_100_48), .C2 (n_98_43) );
AOI211_X1 g_99_47 (.ZN (n_99_47), .A (n_98_50), .B (n_100_47), .C1 (n_98_47), .C2 (n_100_44) );
AOI211_X1 g_100_45 (.ZN (n_100_45), .A (n_100_49), .B (n_99_49), .C1 (n_99_45), .C2 (n_99_46) );
AOI211_X1 g_99_43 (.ZN (n_99_43), .A (n_99_47), .B (n_100_51), .C1 (n_100_47), .C2 (n_100_48) );
AOI211_X1 g_97_42 (.ZN (n_97_42), .A (n_100_45), .B (n_98_50), .C1 (n_99_49), .C2 (n_98_47) );
AOI211_X1 g_98_44 (.ZN (n_98_44), .A (n_99_43), .B (n_100_49), .C1 (n_100_51), .C2 (n_99_45) );
AOI211_X1 g_96_45 (.ZN (n_96_45), .A (n_97_42), .B (n_99_47), .C1 (n_98_50), .C2 (n_100_47) );
AOI211_X1 g_95_43 (.ZN (n_95_43), .A (n_98_44), .B (n_100_45), .C1 (n_100_49), .C2 (n_99_49) );
AOI211_X1 g_97_44 (.ZN (n_97_44), .A (n_96_45), .B (n_99_43), .C1 (n_99_47), .C2 (n_100_51) );
AOI211_X1 g_98_46 (.ZN (n_98_46), .A (n_95_43), .B (n_97_42), .C1 (n_100_45), .C2 (n_98_50) );
AOI211_X1 g_97_48 (.ZN (n_97_48), .A (n_97_44), .B (n_98_44), .C1 (n_99_43), .C2 (n_100_49) );
AOI211_X1 g_96_46 (.ZN (n_96_46), .A (n_98_46), .B (n_96_45), .C1 (n_97_42), .C2 (n_99_47) );
AOI211_X1 g_98_45 (.ZN (n_98_45), .A (n_97_48), .B (n_95_43), .C1 (n_98_44), .C2 (n_100_45) );
AOI211_X1 g_96_44 (.ZN (n_96_44), .A (n_96_46), .B (n_97_44), .C1 (n_96_45), .C2 (n_99_43) );
AOI211_X1 g_94_45 (.ZN (n_94_45), .A (n_98_45), .B (n_98_46), .C1 (n_95_43), .C2 (n_97_42) );
AOI211_X1 g_92_46 (.ZN (n_92_46), .A (n_96_44), .B (n_97_48), .C1 (n_97_44), .C2 (n_98_44) );
AOI211_X1 g_93_44 (.ZN (n_93_44), .A (n_94_45), .B (n_96_46), .C1 (n_98_46), .C2 (n_96_45) );
AOI211_X1 g_91_45 (.ZN (n_91_45), .A (n_92_46), .B (n_98_45), .C1 (n_97_48), .C2 (n_95_43) );
AOI211_X1 g_89_46 (.ZN (n_89_46), .A (n_93_44), .B (n_96_44), .C1 (n_96_46), .C2 (n_97_44) );
AOI211_X1 g_88_48 (.ZN (n_88_48), .A (n_91_45), .B (n_94_45), .C1 (n_98_45), .C2 (n_98_46) );
AOI211_X1 g_90_47 (.ZN (n_90_47), .A (n_89_46), .B (n_92_46), .C1 (n_96_44), .C2 (n_97_48) );
AOI211_X1 g_89_49 (.ZN (n_89_49), .A (n_88_48), .B (n_93_44), .C1 (n_94_45), .C2 (n_96_46) );
AOI211_X1 g_87_48 (.ZN (n_87_48), .A (n_90_47), .B (n_91_45), .C1 (n_92_46), .C2 (n_98_45) );
AOI211_X1 g_89_47 (.ZN (n_89_47), .A (n_89_49), .B (n_89_46), .C1 (n_93_44), .C2 (n_96_44) );
AOI211_X1 g_91_46 (.ZN (n_91_46), .A (n_87_48), .B (n_88_48), .C1 (n_91_45), .C2 (n_94_45) );
AOI211_X1 g_93_45 (.ZN (n_93_45), .A (n_89_47), .B (n_90_47), .C1 (n_89_46), .C2 (n_92_46) );
AOI211_X1 g_95_46 (.ZN (n_95_46), .A (n_91_46), .B (n_89_49), .C1 (n_88_48), .C2 (n_93_44) );
AOI211_X1 g_97_47 (.ZN (n_97_47), .A (n_93_45), .B (n_87_48), .C1 (n_90_47), .C2 (n_91_45) );
AOI211_X1 g_98_49 (.ZN (n_98_49), .A (n_95_46), .B (n_89_47), .C1 (n_89_49), .C2 (n_89_46) );
AOI211_X1 g_99_51 (.ZN (n_99_51), .A (n_97_47), .B (n_91_46), .C1 (n_87_48), .C2 (n_88_48) );
AOI211_X1 g_100_53 (.ZN (n_100_53), .A (n_98_49), .B (n_93_45), .C1 (n_89_47), .C2 (n_90_47) );
AOI211_X1 g_98_54 (.ZN (n_98_54), .A (n_99_51), .B (n_95_46), .C1 (n_91_46), .C2 (n_89_49) );
AOI211_X1 g_100_55 (.ZN (n_100_55), .A (n_100_53), .B (n_97_47), .C1 (n_93_45), .C2 (n_87_48) );
AOI211_X1 g_99_53 (.ZN (n_99_53), .A (n_98_54), .B (n_98_49), .C1 (n_95_46), .C2 (n_89_47) );
AOI211_X1 g_97_52 (.ZN (n_97_52), .A (n_100_55), .B (n_99_51), .C1 (n_97_47), .C2 (n_91_46) );
AOI211_X1 g_96_50 (.ZN (n_96_50), .A (n_99_53), .B (n_100_53), .C1 (n_98_49), .C2 (n_93_45) );
AOI211_X1 g_98_51 (.ZN (n_98_51), .A (n_97_52), .B (n_98_54), .C1 (n_99_51), .C2 (n_95_46) );
AOI211_X1 g_100_52 (.ZN (n_100_52), .A (n_96_50), .B (n_100_55), .C1 (n_100_53), .C2 (n_97_47) );
AOI211_X1 g_99_50 (.ZN (n_99_50), .A (n_98_51), .B (n_99_53), .C1 (n_98_54), .C2 (n_98_49) );
AOI211_X1 g_98_48 (.ZN (n_98_48), .A (n_100_52), .B (n_97_52), .C1 (n_100_55), .C2 (n_99_51) );
AOI211_X1 g_97_46 (.ZN (n_97_46), .A (n_99_50), .B (n_96_50), .C1 (n_99_53), .C2 (n_100_53) );
AOI211_X1 g_95_45 (.ZN (n_95_45), .A (n_98_48), .B (n_98_51), .C1 (n_97_52), .C2 (n_98_54) );
AOI211_X1 g_93_46 (.ZN (n_93_46), .A (n_97_46), .B (n_100_52), .C1 (n_96_50), .C2 (n_100_55) );
AOI211_X1 g_95_47 (.ZN (n_95_47), .A (n_95_45), .B (n_99_50), .C1 (n_98_51), .C2 (n_99_53) );
AOI211_X1 g_96_49 (.ZN (n_96_49), .A (n_93_46), .B (n_98_48), .C1 (n_100_52), .C2 (n_97_52) );
AOI211_X1 g_97_51 (.ZN (n_97_51), .A (n_95_47), .B (n_97_46), .C1 (n_99_50), .C2 (n_96_50) );
AOI211_X1 g_98_53 (.ZN (n_98_53), .A (n_96_49), .B (n_95_45), .C1 (n_98_48), .C2 (n_98_51) );
AOI211_X1 g_99_55 (.ZN (n_99_55), .A (n_97_51), .B (n_93_46), .C1 (n_97_46), .C2 (n_100_52) );
AOI211_X1 g_100_57 (.ZN (n_100_57), .A (n_98_53), .B (n_95_47), .C1 (n_95_45), .C2 (n_99_50) );
AOI211_X1 g_98_58 (.ZN (n_98_58), .A (n_99_55), .B (n_96_49), .C1 (n_93_46), .C2 (n_98_48) );
AOI211_X1 g_100_59 (.ZN (n_100_59), .A (n_100_57), .B (n_97_51), .C1 (n_95_47), .C2 (n_97_46) );
AOI211_X1 g_99_57 (.ZN (n_99_57), .A (n_98_58), .B (n_98_53), .C1 (n_96_49), .C2 (n_95_45) );
AOI211_X1 g_97_56 (.ZN (n_97_56), .A (n_100_59), .B (n_99_55), .C1 (n_97_51), .C2 (n_93_46) );
AOI211_X1 g_96_54 (.ZN (n_96_54), .A (n_99_57), .B (n_100_57), .C1 (n_98_53), .C2 (n_95_47) );
AOI211_X1 g_98_55 (.ZN (n_98_55), .A (n_97_56), .B (n_98_58), .C1 (n_99_55), .C2 (n_96_49) );
AOI211_X1 g_100_56 (.ZN (n_100_56), .A (n_96_54), .B (n_100_59), .C1 (n_100_57), .C2 (n_97_51) );
AOI211_X1 g_99_54 (.ZN (n_99_54), .A (n_98_55), .B (n_99_57), .C1 (n_98_58), .C2 (n_98_53) );
AOI211_X1 g_98_52 (.ZN (n_98_52), .A (n_100_56), .B (n_97_56), .C1 (n_100_59), .C2 (n_99_55) );
AOI211_X1 g_97_50 (.ZN (n_97_50), .A (n_99_54), .B (n_96_54), .C1 (n_99_57), .C2 (n_100_57) );
AOI211_X1 g_96_48 (.ZN (n_96_48), .A (n_98_52), .B (n_98_55), .C1 (n_97_56), .C2 (n_98_58) );
AOI211_X1 g_94_47 (.ZN (n_94_47), .A (n_97_50), .B (n_100_56), .C1 (n_96_54), .C2 (n_100_59) );
AOI211_X1 g_92_48 (.ZN (n_92_48), .A (n_96_48), .B (n_99_54), .C1 (n_98_55), .C2 (n_99_57) );
AOI211_X1 g_94_49 (.ZN (n_94_49), .A (n_94_47), .B (n_98_52), .C1 (n_100_56), .C2 (n_97_56) );
AOI211_X1 g_93_47 (.ZN (n_93_47), .A (n_92_48), .B (n_97_50), .C1 (n_99_54), .C2 (n_96_54) );
AOI211_X1 g_91_48 (.ZN (n_91_48), .A (n_94_49), .B (n_96_48), .C1 (n_98_52), .C2 (n_98_55) );
AOI211_X1 g_92_50 (.ZN (n_92_50), .A (n_93_47), .B (n_94_47), .C1 (n_97_50), .C2 (n_100_56) );
AOI211_X1 g_90_49 (.ZN (n_90_49), .A (n_91_48), .B (n_92_48), .C1 (n_96_48), .C2 (n_99_54) );
AOI211_X1 g_91_47 (.ZN (n_91_47), .A (n_92_50), .B (n_94_49), .C1 (n_94_47), .C2 (n_98_52) );
AOI211_X1 g_89_48 (.ZN (n_89_48), .A (n_90_49), .B (n_93_47), .C1 (n_92_48), .C2 (n_97_50) );
AOI211_X1 g_87_49 (.ZN (n_87_49), .A (n_91_47), .B (n_91_48), .C1 (n_94_49), .C2 (n_96_48) );
AOI211_X1 g_85_48 (.ZN (n_85_48), .A (n_89_48), .B (n_92_50), .C1 (n_93_47), .C2 (n_94_47) );
AOI211_X1 g_83_49 (.ZN (n_83_49), .A (n_87_49), .B (n_90_49), .C1 (n_91_48), .C2 (n_92_48) );
AOI211_X1 g_81_50 (.ZN (n_81_50), .A (n_85_48), .B (n_91_47), .C1 (n_92_50), .C2 (n_94_49) );
AOI211_X1 g_83_51 (.ZN (n_83_51), .A (n_83_49), .B (n_89_48), .C1 (n_90_49), .C2 (n_93_47) );
AOI211_X1 g_85_50 (.ZN (n_85_50), .A (n_81_50), .B (n_87_49), .C1 (n_91_47), .C2 (n_91_48) );
AOI211_X1 g_84_52 (.ZN (n_84_52), .A (n_83_51), .B (n_85_48), .C1 (n_89_48), .C2 (n_92_50) );
AOI211_X1 g_83_50 (.ZN (n_83_50), .A (n_85_50), .B (n_83_49), .C1 (n_87_49), .C2 (n_90_49) );
AOI211_X1 g_85_49 (.ZN (n_85_49), .A (n_84_52), .B (n_81_50), .C1 (n_85_48), .C2 (n_91_47) );
AOI211_X1 g_87_50 (.ZN (n_87_50), .A (n_83_50), .B (n_83_51), .C1 (n_83_49), .C2 (n_89_48) );
AOI211_X1 g_85_51 (.ZN (n_85_51), .A (n_85_49), .B (n_85_50), .C1 (n_81_50), .C2 (n_87_49) );
AOI211_X1 g_86_49 (.ZN (n_86_49), .A (n_87_50), .B (n_84_52), .C1 (n_83_51), .C2 (n_85_48) );
AOI211_X1 g_84_50 (.ZN (n_84_50), .A (n_85_51), .B (n_83_50), .C1 (n_85_50), .C2 (n_83_49) );
AOI211_X1 g_82_51 (.ZN (n_82_51), .A (n_86_49), .B (n_85_49), .C1 (n_84_52), .C2 (n_81_50) );
AOI211_X1 g_80_50 (.ZN (n_80_50), .A (n_84_50), .B (n_87_50), .C1 (n_83_50), .C2 (n_83_51) );
AOI211_X1 g_78_51 (.ZN (n_78_51), .A (n_82_51), .B (n_85_51), .C1 (n_85_49), .C2 (n_85_50) );
AOI211_X1 g_76_52 (.ZN (n_76_52), .A (n_80_50), .B (n_86_49), .C1 (n_87_50), .C2 (n_84_52) );
AOI211_X1 g_74_53 (.ZN (n_74_53), .A (n_78_51), .B (n_84_50), .C1 (n_85_51), .C2 (n_83_50) );
AOI211_X1 g_72_54 (.ZN (n_72_54), .A (n_76_52), .B (n_82_51), .C1 (n_86_49), .C2 (n_85_49) );
AOI211_X1 g_70_55 (.ZN (n_70_55), .A (n_74_53), .B (n_80_50), .C1 (n_84_50), .C2 (n_87_50) );
AOI211_X1 g_68_56 (.ZN (n_68_56), .A (n_72_54), .B (n_78_51), .C1 (n_82_51), .C2 (n_85_51) );
AOI211_X1 g_66_57 (.ZN (n_66_57), .A (n_70_55), .B (n_76_52), .C1 (n_80_50), .C2 (n_86_49) );
AOI211_X1 g_64_58 (.ZN (n_64_58), .A (n_68_56), .B (n_74_53), .C1 (n_78_51), .C2 (n_84_50) );
AOI211_X1 g_63_56 (.ZN (n_63_56), .A (n_66_57), .B (n_72_54), .C1 (n_76_52), .C2 (n_82_51) );
AOI211_X1 g_61_57 (.ZN (n_61_57), .A (n_64_58), .B (n_70_55), .C1 (n_74_53), .C2 (n_80_50) );
AOI211_X1 g_59_58 (.ZN (n_59_58), .A (n_63_56), .B (n_68_56), .C1 (n_72_54), .C2 (n_78_51) );
AOI211_X1 g_57_59 (.ZN (n_57_59), .A (n_61_57), .B (n_66_57), .C1 (n_70_55), .C2 (n_76_52) );
AOI211_X1 g_56_61 (.ZN (n_56_61), .A (n_59_58), .B (n_64_58), .C1 (n_68_56), .C2 (n_74_53) );
AOI211_X1 g_58_60 (.ZN (n_58_60), .A (n_57_59), .B (n_63_56), .C1 (n_66_57), .C2 (n_72_54) );
AOI211_X1 g_60_59 (.ZN (n_60_59), .A (n_56_61), .B (n_61_57), .C1 (n_64_58), .C2 (n_70_55) );
AOI211_X1 g_62_58 (.ZN (n_62_58), .A (n_58_60), .B (n_59_58), .C1 (n_63_56), .C2 (n_68_56) );
AOI211_X1 g_64_57 (.ZN (n_64_57), .A (n_60_59), .B (n_57_59), .C1 (n_61_57), .C2 (n_66_57) );
AOI211_X1 g_63_59 (.ZN (n_63_59), .A (n_62_58), .B (n_56_61), .C1 (n_59_58), .C2 (n_64_58) );
AOI211_X1 g_65_58 (.ZN (n_65_58), .A (n_64_57), .B (n_58_60), .C1 (n_57_59), .C2 (n_63_56) );
AOI211_X1 g_67_59 (.ZN (n_67_59), .A (n_63_59), .B (n_60_59), .C1 (n_56_61), .C2 (n_61_57) );
AOI211_X1 g_68_57 (.ZN (n_68_57), .A (n_65_58), .B (n_62_58), .C1 (n_58_60), .C2 (n_59_58) );
AOI211_X1 g_70_56 (.ZN (n_70_56), .A (n_67_59), .B (n_64_57), .C1 (n_60_59), .C2 (n_57_59) );
AOI211_X1 g_72_55 (.ZN (n_72_55), .A (n_68_57), .B (n_63_59), .C1 (n_62_58), .C2 (n_56_61) );
AOI211_X1 g_74_54 (.ZN (n_74_54), .A (n_70_56), .B (n_65_58), .C1 (n_64_57), .C2 (n_58_60) );
AOI211_X1 g_76_53 (.ZN (n_76_53), .A (n_72_55), .B (n_67_59), .C1 (n_63_59), .C2 (n_60_59) );
AOI211_X1 g_78_52 (.ZN (n_78_52), .A (n_74_54), .B (n_68_57), .C1 (n_65_58), .C2 (n_62_58) );
AOI211_X1 g_80_51 (.ZN (n_80_51), .A (n_76_53), .B (n_70_56), .C1 (n_67_59), .C2 (n_64_57) );
AOI211_X1 g_82_50 (.ZN (n_82_50), .A (n_78_52), .B (n_72_55), .C1 (n_68_57), .C2 (n_63_59) );
AOI211_X1 g_81_52 (.ZN (n_81_52), .A (n_80_51), .B (n_74_54), .C1 (n_70_56), .C2 (n_65_58) );
AOI211_X1 g_79_53 (.ZN (n_79_53), .A (n_82_50), .B (n_76_53), .C1 (n_72_55), .C2 (n_67_59) );
AOI211_X1 g_77_54 (.ZN (n_77_54), .A (n_81_52), .B (n_78_52), .C1 (n_74_54), .C2 (n_68_57) );
AOI211_X1 g_75_55 (.ZN (n_75_55), .A (n_79_53), .B (n_80_51), .C1 (n_76_53), .C2 (n_70_56) );
AOI211_X1 g_73_56 (.ZN (n_73_56), .A (n_77_54), .B (n_82_50), .C1 (n_78_52), .C2 (n_72_55) );
AOI211_X1 g_71_57 (.ZN (n_71_57), .A (n_75_55), .B (n_81_52), .C1 (n_80_51), .C2 (n_74_54) );
AOI211_X1 g_69_58 (.ZN (n_69_58), .A (n_73_56), .B (n_79_53), .C1 (n_82_50), .C2 (n_76_53) );
AOI211_X1 g_68_60 (.ZN (n_68_60), .A (n_71_57), .B (n_77_54), .C1 (n_81_52), .C2 (n_78_52) );
AOI211_X1 g_66_59 (.ZN (n_66_59), .A (n_69_58), .B (n_75_55), .C1 (n_79_53), .C2 (n_80_51) );
AOI211_X1 g_65_57 (.ZN (n_65_57), .A (n_68_60), .B (n_73_56), .C1 (n_77_54), .C2 (n_82_50) );
AOI211_X1 g_63_58 (.ZN (n_63_58), .A (n_66_59), .B (n_71_57), .C1 (n_75_55), .C2 (n_81_52) );
AOI211_X1 g_61_59 (.ZN (n_61_59), .A (n_65_57), .B (n_69_58), .C1 (n_73_56), .C2 (n_79_53) );
AOI211_X1 g_59_60 (.ZN (n_59_60), .A (n_63_58), .B (n_68_60), .C1 (n_71_57), .C2 (n_77_54) );
AOI211_X1 g_57_61 (.ZN (n_57_61), .A (n_61_59), .B (n_66_59), .C1 (n_69_58), .C2 (n_75_55) );
AOI211_X1 g_55_62 (.ZN (n_55_62), .A (n_59_60), .B (n_65_57), .C1 (n_68_60), .C2 (n_73_56) );
AOI211_X1 g_53_61 (.ZN (n_53_61), .A (n_57_61), .B (n_63_58), .C1 (n_66_59), .C2 (n_71_57) );
AOI211_X1 g_51_62 (.ZN (n_51_62), .A (n_55_62), .B (n_61_59), .C1 (n_65_57), .C2 (n_69_58) );
AOI211_X1 g_49_63 (.ZN (n_49_63), .A (n_53_61), .B (n_59_60), .C1 (n_63_58), .C2 (n_68_60) );
AOI211_X1 g_47_64 (.ZN (n_47_64), .A (n_51_62), .B (n_57_61), .C1 (n_61_59), .C2 (n_66_59) );
AOI211_X1 g_45_65 (.ZN (n_45_65), .A (n_49_63), .B (n_55_62), .C1 (n_59_60), .C2 (n_65_57) );
AOI211_X1 g_43_66 (.ZN (n_43_66), .A (n_47_64), .B (n_53_61), .C1 (n_57_61), .C2 (n_63_58) );
AOI211_X1 g_41_67 (.ZN (n_41_67), .A (n_45_65), .B (n_51_62), .C1 (n_55_62), .C2 (n_61_59) );
AOI211_X1 g_39_68 (.ZN (n_39_68), .A (n_43_66), .B (n_49_63), .C1 (n_53_61), .C2 (n_59_60) );
AOI211_X1 g_37_69 (.ZN (n_37_69), .A (n_41_67), .B (n_47_64), .C1 (n_51_62), .C2 (n_57_61) );
AOI211_X1 g_35_70 (.ZN (n_35_70), .A (n_39_68), .B (n_45_65), .C1 (n_49_63), .C2 (n_55_62) );
AOI211_X1 g_36_68 (.ZN (n_36_68), .A (n_37_69), .B (n_43_66), .C1 (n_47_64), .C2 (n_53_61) );
AOI211_X1 g_34_69 (.ZN (n_34_69), .A (n_35_70), .B (n_41_67), .C1 (n_45_65), .C2 (n_51_62) );
AOI211_X1 g_32_70 (.ZN (n_32_70), .A (n_36_68), .B (n_39_68), .C1 (n_43_66), .C2 (n_49_63) );
AOI211_X1 g_30_71 (.ZN (n_30_71), .A (n_34_69), .B (n_37_69), .C1 (n_41_67), .C2 (n_47_64) );
AOI211_X1 g_28_72 (.ZN (n_28_72), .A (n_32_70), .B (n_35_70), .C1 (n_39_68), .C2 (n_45_65) );
AOI211_X1 g_26_73 (.ZN (n_26_73), .A (n_30_71), .B (n_36_68), .C1 (n_37_69), .C2 (n_43_66) );
AOI211_X1 g_24_74 (.ZN (n_24_74), .A (n_28_72), .B (n_34_69), .C1 (n_35_70), .C2 (n_41_67) );
AOI211_X1 g_22_75 (.ZN (n_22_75), .A (n_26_73), .B (n_32_70), .C1 (n_36_68), .C2 (n_39_68) );
AOI211_X1 g_20_76 (.ZN (n_20_76), .A (n_24_74), .B (n_30_71), .C1 (n_34_69), .C2 (n_37_69) );
AOI211_X1 g_18_77 (.ZN (n_18_77), .A (n_22_75), .B (n_28_72), .C1 (n_32_70), .C2 (n_35_70) );
AOI211_X1 g_16_78 (.ZN (n_16_78), .A (n_20_76), .B (n_26_73), .C1 (n_30_71), .C2 (n_36_68) );
AOI211_X1 g_14_79 (.ZN (n_14_79), .A (n_18_77), .B (n_24_74), .C1 (n_28_72), .C2 (n_34_69) );
AOI211_X1 g_16_80 (.ZN (n_16_80), .A (n_16_78), .B (n_22_75), .C1 (n_26_73), .C2 (n_32_70) );
AOI211_X1 g_18_79 (.ZN (n_18_79), .A (n_14_79), .B (n_20_76), .C1 (n_24_74), .C2 (n_30_71) );
AOI211_X1 g_19_77 (.ZN (n_19_77), .A (n_16_80), .B (n_18_77), .C1 (n_22_75), .C2 (n_28_72) );
AOI211_X1 g_21_76 (.ZN (n_21_76), .A (n_18_79), .B (n_16_78), .C1 (n_20_76), .C2 (n_26_73) );
AOI211_X1 g_23_75 (.ZN (n_23_75), .A (n_19_77), .B (n_14_79), .C1 (n_18_77), .C2 (n_24_74) );
AOI211_X1 g_25_74 (.ZN (n_25_74), .A (n_21_76), .B (n_16_80), .C1 (n_16_78), .C2 (n_22_75) );
AOI211_X1 g_27_73 (.ZN (n_27_73), .A (n_23_75), .B (n_18_79), .C1 (n_14_79), .C2 (n_20_76) );
AOI211_X1 g_29_72 (.ZN (n_29_72), .A (n_25_74), .B (n_19_77), .C1 (n_16_80), .C2 (n_18_77) );
AOI211_X1 g_31_71 (.ZN (n_31_71), .A (n_27_73), .B (n_21_76), .C1 (n_18_79), .C2 (n_16_78) );
AOI211_X1 g_33_70 (.ZN (n_33_70), .A (n_29_72), .B (n_23_75), .C1 (n_19_77), .C2 (n_14_79) );
AOI211_X1 g_35_69 (.ZN (n_35_69), .A (n_31_71), .B (n_25_74), .C1 (n_21_76), .C2 (n_16_80) );
AOI211_X1 g_37_68 (.ZN (n_37_68), .A (n_33_70), .B (n_27_73), .C1 (n_23_75), .C2 (n_18_79) );
AOI211_X1 g_36_70 (.ZN (n_36_70), .A (n_35_69), .B (n_29_72), .C1 (n_25_74), .C2 (n_19_77) );
AOI211_X1 g_38_69 (.ZN (n_38_69), .A (n_37_68), .B (n_31_71), .C1 (n_27_73), .C2 (n_21_76) );
AOI211_X1 g_40_68 (.ZN (n_40_68), .A (n_36_70), .B (n_33_70), .C1 (n_29_72), .C2 (n_23_75) );
AOI211_X1 g_42_67 (.ZN (n_42_67), .A (n_38_69), .B (n_35_69), .C1 (n_31_71), .C2 (n_25_74) );
AOI211_X1 g_44_66 (.ZN (n_44_66), .A (n_40_68), .B (n_37_68), .C1 (n_33_70), .C2 (n_27_73) );
AOI211_X1 g_46_65 (.ZN (n_46_65), .A (n_42_67), .B (n_36_70), .C1 (n_35_69), .C2 (n_29_72) );
AOI211_X1 g_48_64 (.ZN (n_48_64), .A (n_44_66), .B (n_38_69), .C1 (n_37_68), .C2 (n_31_71) );
AOI211_X1 g_50_63 (.ZN (n_50_63), .A (n_46_65), .B (n_40_68), .C1 (n_36_70), .C2 (n_33_70) );
AOI211_X1 g_52_62 (.ZN (n_52_62), .A (n_48_64), .B (n_42_67), .C1 (n_38_69), .C2 (n_35_69) );
AOI211_X1 g_51_64 (.ZN (n_51_64), .A (n_50_63), .B (n_44_66), .C1 (n_40_68), .C2 (n_37_68) );
AOI211_X1 g_53_63 (.ZN (n_53_63), .A (n_52_62), .B (n_46_65), .C1 (n_42_67), .C2 (n_36_70) );
AOI211_X1 g_52_61 (.ZN (n_52_61), .A (n_51_64), .B (n_48_64), .C1 (n_44_66), .C2 (n_38_69) );
AOI211_X1 g_50_62 (.ZN (n_50_62), .A (n_53_63), .B (n_50_63), .C1 (n_46_65), .C2 (n_40_68) );
AOI211_X1 g_48_63 (.ZN (n_48_63), .A (n_52_61), .B (n_52_62), .C1 (n_48_64), .C2 (n_42_67) );
AOI211_X1 g_46_64 (.ZN (n_46_64), .A (n_50_62), .B (n_51_64), .C1 (n_50_63), .C2 (n_44_66) );
AOI211_X1 g_44_65 (.ZN (n_44_65), .A (n_48_63), .B (n_53_63), .C1 (n_52_62), .C2 (n_46_65) );
AOI211_X1 g_42_66 (.ZN (n_42_66), .A (n_46_64), .B (n_52_61), .C1 (n_51_64), .C2 (n_48_64) );
AOI211_X1 g_40_67 (.ZN (n_40_67), .A (n_44_65), .B (n_50_62), .C1 (n_53_63), .C2 (n_50_63) );
AOI211_X1 g_38_68 (.ZN (n_38_68), .A (n_42_66), .B (n_48_63), .C1 (n_52_61), .C2 (n_52_62) );
AOI211_X1 g_36_69 (.ZN (n_36_69), .A (n_40_67), .B (n_46_64), .C1 (n_50_62), .C2 (n_51_64) );
AOI211_X1 g_34_70 (.ZN (n_34_70), .A (n_38_68), .B (n_44_65), .C1 (n_48_63), .C2 (n_53_63) );
AOI211_X1 g_32_71 (.ZN (n_32_71), .A (n_36_69), .B (n_42_66), .C1 (n_46_64), .C2 (n_52_61) );
AOI211_X1 g_30_72 (.ZN (n_30_72), .A (n_34_70), .B (n_40_67), .C1 (n_44_65), .C2 (n_50_62) );
AOI211_X1 g_28_73 (.ZN (n_28_73), .A (n_32_71), .B (n_38_68), .C1 (n_42_66), .C2 (n_48_63) );
AOI211_X1 g_26_74 (.ZN (n_26_74), .A (n_30_72), .B (n_36_69), .C1 (n_40_67), .C2 (n_46_64) );
AOI211_X1 g_24_75 (.ZN (n_24_75), .A (n_28_73), .B (n_34_70), .C1 (n_38_68), .C2 (n_44_65) );
AOI211_X1 g_22_76 (.ZN (n_22_76), .A (n_26_74), .B (n_32_71), .C1 (n_36_69), .C2 (n_42_66) );
AOI211_X1 g_20_77 (.ZN (n_20_77), .A (n_24_75), .B (n_30_72), .C1 (n_34_70), .C2 (n_40_67) );
AOI211_X1 g_18_78 (.ZN (n_18_78), .A (n_22_76), .B (n_28_73), .C1 (n_32_71), .C2 (n_38_68) );
AOI211_X1 g_16_79 (.ZN (n_16_79), .A (n_20_77), .B (n_26_74), .C1 (n_30_72), .C2 (n_36_69) );
AOI211_X1 g_14_78 (.ZN (n_14_78), .A (n_18_78), .B (n_24_75), .C1 (n_28_73), .C2 (n_34_70) );
AOI211_X1 g_12_79 (.ZN (n_12_79), .A (n_16_79), .B (n_22_76), .C1 (n_26_74), .C2 (n_32_71) );
AOI211_X1 g_11_81 (.ZN (n_11_81), .A (n_14_78), .B (n_20_77), .C1 (n_24_75), .C2 (n_30_72) );
AOI211_X1 g_13_80 (.ZN (n_13_80), .A (n_12_79), .B (n_18_78), .C1 (n_22_76), .C2 (n_28_73) );
AOI211_X1 g_15_79 (.ZN (n_15_79), .A (n_11_81), .B (n_16_79), .C1 (n_20_77), .C2 (n_26_74) );
AOI211_X1 g_14_81 (.ZN (n_14_81), .A (n_13_80), .B (n_14_78), .C1 (n_18_78), .C2 (n_24_75) );
AOI211_X1 g_12_82 (.ZN (n_12_82), .A (n_15_79), .B (n_12_79), .C1 (n_16_79), .C2 (n_22_76) );
AOI211_X1 g_11_80 (.ZN (n_11_80), .A (n_14_81), .B (n_11_81), .C1 (n_14_78), .C2 (n_20_77) );
AOI211_X1 g_10_82 (.ZN (n_10_82), .A (n_12_82), .B (n_13_80), .C1 (n_12_79), .C2 (n_18_78) );
AOI211_X1 g_12_81 (.ZN (n_12_81), .A (n_11_80), .B (n_15_79), .C1 (n_11_81), .C2 (n_16_79) );
AOI211_X1 g_14_80 (.ZN (n_14_80), .A (n_10_82), .B (n_14_81), .C1 (n_13_80), .C2 (n_14_78) );
AOI211_X1 g_13_82 (.ZN (n_13_82), .A (n_12_81), .B (n_12_82), .C1 (n_15_79), .C2 (n_12_79) );
AOI211_X1 g_15_81 (.ZN (n_15_81), .A (n_14_80), .B (n_11_80), .C1 (n_14_81), .C2 (n_11_81) );
AOI211_X1 g_17_80 (.ZN (n_17_80), .A (n_13_82), .B (n_10_82), .C1 (n_12_82), .C2 (n_13_80) );
AOI211_X1 g_19_79 (.ZN (n_19_79), .A (n_15_81), .B (n_12_81), .C1 (n_11_80), .C2 (n_15_79) );
AOI211_X1 g_21_78 (.ZN (n_21_78), .A (n_17_80), .B (n_14_80), .C1 (n_10_82), .C2 (n_14_81) );
AOI211_X1 g_23_77 (.ZN (n_23_77), .A (n_19_79), .B (n_13_82), .C1 (n_12_81), .C2 (n_12_82) );
AOI211_X1 g_25_76 (.ZN (n_25_76), .A (n_21_78), .B (n_15_81), .C1 (n_14_80), .C2 (n_11_80) );
AOI211_X1 g_27_75 (.ZN (n_27_75), .A (n_23_77), .B (n_17_80), .C1 (n_13_82), .C2 (n_10_82) );
AOI211_X1 g_29_74 (.ZN (n_29_74), .A (n_25_76), .B (n_19_79), .C1 (n_15_81), .C2 (n_12_81) );
AOI211_X1 g_31_73 (.ZN (n_31_73), .A (n_27_75), .B (n_21_78), .C1 (n_17_80), .C2 (n_14_80) );
AOI211_X1 g_33_72 (.ZN (n_33_72), .A (n_29_74), .B (n_23_77), .C1 (n_19_79), .C2 (n_13_82) );
AOI211_X1 g_35_71 (.ZN (n_35_71), .A (n_31_73), .B (n_25_76), .C1 (n_21_78), .C2 (n_15_81) );
AOI211_X1 g_37_70 (.ZN (n_37_70), .A (n_33_72), .B (n_27_75), .C1 (n_23_77), .C2 (n_17_80) );
AOI211_X1 g_39_69 (.ZN (n_39_69), .A (n_35_71), .B (n_29_74), .C1 (n_25_76), .C2 (n_19_79) );
AOI211_X1 g_41_68 (.ZN (n_41_68), .A (n_37_70), .B (n_31_73), .C1 (n_27_75), .C2 (n_21_78) );
AOI211_X1 g_43_67 (.ZN (n_43_67), .A (n_39_69), .B (n_33_72), .C1 (n_29_74), .C2 (n_23_77) );
AOI211_X1 g_45_66 (.ZN (n_45_66), .A (n_41_68), .B (n_35_71), .C1 (n_31_73), .C2 (n_25_76) );
AOI211_X1 g_47_65 (.ZN (n_47_65), .A (n_43_67), .B (n_37_70), .C1 (n_33_72), .C2 (n_27_75) );
AOI211_X1 g_49_64 (.ZN (n_49_64), .A (n_45_66), .B (n_39_69), .C1 (n_35_71), .C2 (n_29_74) );
AOI211_X1 g_51_63 (.ZN (n_51_63), .A (n_47_65), .B (n_41_68), .C1 (n_37_70), .C2 (n_31_73) );
AOI211_X1 g_53_62 (.ZN (n_53_62), .A (n_49_64), .B (n_43_67), .C1 (n_39_69), .C2 (n_33_72) );
AOI211_X1 g_55_61 (.ZN (n_55_61), .A (n_51_63), .B (n_45_66), .C1 (n_41_68), .C2 (n_35_71) );
AOI211_X1 g_54_63 (.ZN (n_54_63), .A (n_53_62), .B (n_47_65), .C1 (n_43_67), .C2 (n_37_70) );
AOI211_X1 g_56_62 (.ZN (n_56_62), .A (n_55_61), .B (n_49_64), .C1 (n_45_66), .C2 (n_39_69) );
AOI211_X1 g_58_61 (.ZN (n_58_61), .A (n_54_63), .B (n_51_63), .C1 (n_47_65), .C2 (n_41_68) );
AOI211_X1 g_60_60 (.ZN (n_60_60), .A (n_56_62), .B (n_53_62), .C1 (n_49_64), .C2 (n_43_67) );
AOI211_X1 g_62_59 (.ZN (n_62_59), .A (n_58_61), .B (n_55_61), .C1 (n_51_63), .C2 (n_45_66) );
AOI211_X1 g_64_60 (.ZN (n_64_60), .A (n_60_60), .B (n_54_63), .C1 (n_53_62), .C2 (n_47_65) );
AOI211_X1 g_62_61 (.ZN (n_62_61), .A (n_62_59), .B (n_56_62), .C1 (n_55_61), .C2 (n_49_64) );
AOI211_X1 g_60_62 (.ZN (n_60_62), .A (n_64_60), .B (n_58_61), .C1 (n_54_63), .C2 (n_51_63) );
AOI211_X1 g_61_60 (.ZN (n_61_60), .A (n_62_61), .B (n_60_60), .C1 (n_56_62), .C2 (n_53_62) );
AOI211_X1 g_59_61 (.ZN (n_59_61), .A (n_60_62), .B (n_62_59), .C1 (n_58_61), .C2 (n_55_61) );
AOI211_X1 g_57_62 (.ZN (n_57_62), .A (n_61_60), .B (n_64_60), .C1 (n_60_60), .C2 (n_54_63) );
AOI211_X1 g_55_63 (.ZN (n_55_63), .A (n_59_61), .B (n_62_61), .C1 (n_62_59), .C2 (n_56_62) );
AOI211_X1 g_53_64 (.ZN (n_53_64), .A (n_57_62), .B (n_60_62), .C1 (n_64_60), .C2 (n_58_61) );
AOI211_X1 g_54_62 (.ZN (n_54_62), .A (n_55_63), .B (n_61_60), .C1 (n_62_61), .C2 (n_60_60) );
AOI211_X1 g_52_63 (.ZN (n_52_63), .A (n_53_64), .B (n_59_61), .C1 (n_60_62), .C2 (n_62_59) );
AOI211_X1 g_50_64 (.ZN (n_50_64), .A (n_54_62), .B (n_57_62), .C1 (n_61_60), .C2 (n_64_60) );
AOI211_X1 g_48_65 (.ZN (n_48_65), .A (n_52_63), .B (n_55_63), .C1 (n_59_61), .C2 (n_62_61) );
AOI211_X1 g_46_66 (.ZN (n_46_66), .A (n_50_64), .B (n_53_64), .C1 (n_57_62), .C2 (n_60_62) );
AOI211_X1 g_44_67 (.ZN (n_44_67), .A (n_48_65), .B (n_54_62), .C1 (n_55_63), .C2 (n_61_60) );
AOI211_X1 g_42_68 (.ZN (n_42_68), .A (n_46_66), .B (n_52_63), .C1 (n_53_64), .C2 (n_59_61) );
AOI211_X1 g_40_69 (.ZN (n_40_69), .A (n_44_67), .B (n_50_64), .C1 (n_54_62), .C2 (n_57_62) );
AOI211_X1 g_38_70 (.ZN (n_38_70), .A (n_42_68), .B (n_48_65), .C1 (n_52_63), .C2 (n_55_63) );
AOI211_X1 g_36_71 (.ZN (n_36_71), .A (n_40_69), .B (n_46_66), .C1 (n_50_64), .C2 (n_53_64) );
AOI211_X1 g_34_72 (.ZN (n_34_72), .A (n_38_70), .B (n_44_67), .C1 (n_48_65), .C2 (n_54_62) );
AOI211_X1 g_32_73 (.ZN (n_32_73), .A (n_36_71), .B (n_42_68), .C1 (n_46_66), .C2 (n_52_63) );
AOI211_X1 g_33_71 (.ZN (n_33_71), .A (n_34_72), .B (n_40_69), .C1 (n_44_67), .C2 (n_50_64) );
AOI211_X1 g_31_72 (.ZN (n_31_72), .A (n_32_73), .B (n_38_70), .C1 (n_42_68), .C2 (n_48_65) );
AOI211_X1 g_29_73 (.ZN (n_29_73), .A (n_33_71), .B (n_36_71), .C1 (n_40_69), .C2 (n_46_66) );
AOI211_X1 g_27_74 (.ZN (n_27_74), .A (n_31_72), .B (n_34_72), .C1 (n_38_70), .C2 (n_44_67) );
AOI211_X1 g_25_75 (.ZN (n_25_75), .A (n_29_73), .B (n_32_73), .C1 (n_36_71), .C2 (n_42_68) );
AOI211_X1 g_23_76 (.ZN (n_23_76), .A (n_27_74), .B (n_33_71), .C1 (n_34_72), .C2 (n_40_69) );
AOI211_X1 g_21_77 (.ZN (n_21_77), .A (n_25_75), .B (n_31_72), .C1 (n_32_73), .C2 (n_38_70) );
AOI211_X1 g_19_78 (.ZN (n_19_78), .A (n_23_76), .B (n_29_73), .C1 (n_33_71), .C2 (n_36_71) );
AOI211_X1 g_17_79 (.ZN (n_17_79), .A (n_21_77), .B (n_27_74), .C1 (n_31_72), .C2 (n_34_72) );
AOI211_X1 g_15_80 (.ZN (n_15_80), .A (n_19_78), .B (n_25_75), .C1 (n_29_73), .C2 (n_32_73) );
AOI211_X1 g_13_81 (.ZN (n_13_81), .A (n_17_79), .B (n_23_76), .C1 (n_27_74), .C2 (n_33_71) );
AOI211_X1 g_12_83 (.ZN (n_12_83), .A (n_15_80), .B (n_21_77), .C1 (n_25_75), .C2 (n_31_72) );
AOI211_X1 g_14_82 (.ZN (n_14_82), .A (n_13_81), .B (n_19_78), .C1 (n_23_76), .C2 (n_29_73) );
AOI211_X1 g_16_81 (.ZN (n_16_81), .A (n_12_83), .B (n_17_79), .C1 (n_21_77), .C2 (n_27_74) );
AOI211_X1 g_18_80 (.ZN (n_18_80), .A (n_14_82), .B (n_15_80), .C1 (n_19_78), .C2 (n_25_75) );
AOI211_X1 g_20_79 (.ZN (n_20_79), .A (n_16_81), .B (n_13_81), .C1 (n_17_79), .C2 (n_23_76) );
AOI211_X1 g_22_78 (.ZN (n_22_78), .A (n_18_80), .B (n_12_83), .C1 (n_15_80), .C2 (n_21_77) );
AOI211_X1 g_24_77 (.ZN (n_24_77), .A (n_20_79), .B (n_14_82), .C1 (n_13_81), .C2 (n_19_78) );
AOI211_X1 g_26_76 (.ZN (n_26_76), .A (n_22_78), .B (n_16_81), .C1 (n_12_83), .C2 (n_17_79) );
AOI211_X1 g_28_75 (.ZN (n_28_75), .A (n_24_77), .B (n_18_80), .C1 (n_14_82), .C2 (n_15_80) );
AOI211_X1 g_30_74 (.ZN (n_30_74), .A (n_26_76), .B (n_20_79), .C1 (n_16_81), .C2 (n_13_81) );
AOI211_X1 g_29_76 (.ZN (n_29_76), .A (n_28_75), .B (n_22_78), .C1 (n_18_80), .C2 (n_12_83) );
AOI211_X1 g_28_74 (.ZN (n_28_74), .A (n_30_74), .B (n_24_77), .C1 (n_20_79), .C2 (n_14_82) );
AOI211_X1 g_30_73 (.ZN (n_30_73), .A (n_29_76), .B (n_26_76), .C1 (n_22_78), .C2 (n_16_81) );
AOI211_X1 g_32_72 (.ZN (n_32_72), .A (n_28_74), .B (n_28_75), .C1 (n_24_77), .C2 (n_18_80) );
AOI211_X1 g_34_71 (.ZN (n_34_71), .A (n_30_73), .B (n_30_74), .C1 (n_26_76), .C2 (n_20_79) );
AOI211_X1 g_33_73 (.ZN (n_33_73), .A (n_32_72), .B (n_29_76), .C1 (n_28_75), .C2 (n_22_78) );
AOI211_X1 g_35_72 (.ZN (n_35_72), .A (n_34_71), .B (n_28_74), .C1 (n_30_74), .C2 (n_24_77) );
AOI211_X1 g_37_71 (.ZN (n_37_71), .A (n_33_73), .B (n_30_73), .C1 (n_29_76), .C2 (n_26_76) );
AOI211_X1 g_39_70 (.ZN (n_39_70), .A (n_35_72), .B (n_32_72), .C1 (n_28_74), .C2 (n_28_75) );
AOI211_X1 g_41_69 (.ZN (n_41_69), .A (n_37_71), .B (n_34_71), .C1 (n_30_73), .C2 (n_30_74) );
AOI211_X1 g_43_68 (.ZN (n_43_68), .A (n_39_70), .B (n_33_73), .C1 (n_32_72), .C2 (n_29_76) );
AOI211_X1 g_45_67 (.ZN (n_45_67), .A (n_41_69), .B (n_35_72), .C1 (n_34_71), .C2 (n_28_74) );
AOI211_X1 g_47_66 (.ZN (n_47_66), .A (n_43_68), .B (n_37_71), .C1 (n_33_73), .C2 (n_30_73) );
AOI211_X1 g_49_65 (.ZN (n_49_65), .A (n_45_67), .B (n_39_70), .C1 (n_35_72), .C2 (n_32_72) );
AOI211_X1 g_48_67 (.ZN (n_48_67), .A (n_47_66), .B (n_41_69), .C1 (n_37_71), .C2 (n_34_71) );
AOI211_X1 g_50_66 (.ZN (n_50_66), .A (n_49_65), .B (n_43_68), .C1 (n_39_70), .C2 (n_33_73) );
AOI211_X1 g_52_65 (.ZN (n_52_65), .A (n_48_67), .B (n_45_67), .C1 (n_41_69), .C2 (n_35_72) );
AOI211_X1 g_54_64 (.ZN (n_54_64), .A (n_50_66), .B (n_47_66), .C1 (n_43_68), .C2 (n_37_71) );
AOI211_X1 g_56_63 (.ZN (n_56_63), .A (n_52_65), .B (n_49_65), .C1 (n_45_67), .C2 (n_39_70) );
AOI211_X1 g_58_62 (.ZN (n_58_62), .A (n_54_64), .B (n_48_67), .C1 (n_47_66), .C2 (n_41_69) );
AOI211_X1 g_60_61 (.ZN (n_60_61), .A (n_56_63), .B (n_50_66), .C1 (n_49_65), .C2 (n_43_68) );
AOI211_X1 g_62_60 (.ZN (n_62_60), .A (n_58_62), .B (n_52_65), .C1 (n_48_67), .C2 (n_45_67) );
AOI211_X1 g_64_59 (.ZN (n_64_59), .A (n_60_61), .B (n_54_64), .C1 (n_50_66), .C2 (n_47_66) );
AOI211_X1 g_66_58 (.ZN (n_66_58), .A (n_62_60), .B (n_56_63), .C1 (n_52_65), .C2 (n_49_65) );
AOI211_X1 g_65_60 (.ZN (n_65_60), .A (n_64_59), .B (n_58_62), .C1 (n_54_64), .C2 (n_48_67) );
AOI211_X1 g_63_61 (.ZN (n_63_61), .A (n_66_58), .B (n_60_61), .C1 (n_56_63), .C2 (n_50_66) );
AOI211_X1 g_61_62 (.ZN (n_61_62), .A (n_65_60), .B (n_62_60), .C1 (n_58_62), .C2 (n_52_65) );
AOI211_X1 g_59_63 (.ZN (n_59_63), .A (n_63_61), .B (n_64_59), .C1 (n_60_61), .C2 (n_54_64) );
AOI211_X1 g_57_64 (.ZN (n_57_64), .A (n_61_62), .B (n_66_58), .C1 (n_62_60), .C2 (n_56_63) );
AOI211_X1 g_55_65 (.ZN (n_55_65), .A (n_59_63), .B (n_65_60), .C1 (n_64_59), .C2 (n_58_62) );
AOI211_X1 g_53_66 (.ZN (n_53_66), .A (n_57_64), .B (n_63_61), .C1 (n_66_58), .C2 (n_60_61) );
AOI211_X1 g_52_64 (.ZN (n_52_64), .A (n_55_65), .B (n_61_62), .C1 (n_65_60), .C2 (n_62_60) );
AOI211_X1 g_50_65 (.ZN (n_50_65), .A (n_53_66), .B (n_59_63), .C1 (n_63_61), .C2 (n_64_59) );
AOI211_X1 g_48_66 (.ZN (n_48_66), .A (n_52_64), .B (n_57_64), .C1 (n_61_62), .C2 (n_66_58) );
AOI211_X1 g_46_67 (.ZN (n_46_67), .A (n_50_65), .B (n_55_65), .C1 (n_59_63), .C2 (n_65_60) );
AOI211_X1 g_44_68 (.ZN (n_44_68), .A (n_48_66), .B (n_53_66), .C1 (n_57_64), .C2 (n_63_61) );
AOI211_X1 g_42_69 (.ZN (n_42_69), .A (n_46_67), .B (n_52_64), .C1 (n_55_65), .C2 (n_61_62) );
AOI211_X1 g_40_70 (.ZN (n_40_70), .A (n_44_68), .B (n_50_65), .C1 (n_53_66), .C2 (n_59_63) );
AOI211_X1 g_38_71 (.ZN (n_38_71), .A (n_42_69), .B (n_48_66), .C1 (n_52_64), .C2 (n_57_64) );
AOI211_X1 g_36_72 (.ZN (n_36_72), .A (n_40_70), .B (n_46_67), .C1 (n_50_65), .C2 (n_55_65) );
AOI211_X1 g_34_73 (.ZN (n_34_73), .A (n_38_71), .B (n_44_68), .C1 (n_48_66), .C2 (n_53_66) );
AOI211_X1 g_32_74 (.ZN (n_32_74), .A (n_36_72), .B (n_42_69), .C1 (n_46_67), .C2 (n_52_64) );
AOI211_X1 g_30_75 (.ZN (n_30_75), .A (n_34_73), .B (n_40_70), .C1 (n_44_68), .C2 (n_50_65) );
AOI211_X1 g_28_76 (.ZN (n_28_76), .A (n_32_74), .B (n_38_71), .C1 (n_42_69), .C2 (n_48_66) );
AOI211_X1 g_26_75 (.ZN (n_26_75), .A (n_30_75), .B (n_36_72), .C1 (n_40_70), .C2 (n_46_67) );
AOI211_X1 g_24_76 (.ZN (n_24_76), .A (n_28_76), .B (n_34_73), .C1 (n_38_71), .C2 (n_44_68) );
AOI211_X1 g_22_77 (.ZN (n_22_77), .A (n_26_75), .B (n_32_74), .C1 (n_36_72), .C2 (n_42_69) );
AOI211_X1 g_20_78 (.ZN (n_20_78), .A (n_24_76), .B (n_30_75), .C1 (n_34_73), .C2 (n_40_70) );
AOI211_X1 g_19_80 (.ZN (n_19_80), .A (n_22_77), .B (n_28_76), .C1 (n_32_74), .C2 (n_38_71) );
AOI211_X1 g_21_79 (.ZN (n_21_79), .A (n_20_78), .B (n_26_75), .C1 (n_30_75), .C2 (n_36_72) );
AOI211_X1 g_23_78 (.ZN (n_23_78), .A (n_19_80), .B (n_24_76), .C1 (n_28_76), .C2 (n_34_73) );
AOI211_X1 g_25_77 (.ZN (n_25_77), .A (n_21_79), .B (n_22_77), .C1 (n_26_75), .C2 (n_32_74) );
AOI211_X1 g_27_76 (.ZN (n_27_76), .A (n_23_78), .B (n_20_78), .C1 (n_24_76), .C2 (n_30_75) );
AOI211_X1 g_29_75 (.ZN (n_29_75), .A (n_25_77), .B (n_19_80), .C1 (n_22_77), .C2 (n_28_76) );
AOI211_X1 g_31_74 (.ZN (n_31_74), .A (n_27_76), .B (n_21_79), .C1 (n_20_78), .C2 (n_26_75) );
AOI211_X1 g_30_76 (.ZN (n_30_76), .A (n_29_75), .B (n_23_78), .C1 (n_19_80), .C2 (n_24_76) );
AOI211_X1 g_32_75 (.ZN (n_32_75), .A (n_31_74), .B (n_25_77), .C1 (n_21_79), .C2 (n_22_77) );
AOI211_X1 g_34_74 (.ZN (n_34_74), .A (n_30_76), .B (n_27_76), .C1 (n_23_78), .C2 (n_20_78) );
AOI211_X1 g_36_73 (.ZN (n_36_73), .A (n_32_75), .B (n_29_75), .C1 (n_25_77), .C2 (n_19_80) );
AOI211_X1 g_38_72 (.ZN (n_38_72), .A (n_34_74), .B (n_31_74), .C1 (n_27_76), .C2 (n_21_79) );
AOI211_X1 g_40_71 (.ZN (n_40_71), .A (n_36_73), .B (n_30_76), .C1 (n_29_75), .C2 (n_23_78) );
AOI211_X1 g_42_70 (.ZN (n_42_70), .A (n_38_72), .B (n_32_75), .C1 (n_31_74), .C2 (n_25_77) );
AOI211_X1 g_44_69 (.ZN (n_44_69), .A (n_40_71), .B (n_34_74), .C1 (n_30_76), .C2 (n_27_76) );
AOI211_X1 g_46_68 (.ZN (n_46_68), .A (n_42_70), .B (n_36_73), .C1 (n_32_75), .C2 (n_29_75) );
AOI211_X1 g_45_70 (.ZN (n_45_70), .A (n_44_69), .B (n_38_72), .C1 (n_34_74), .C2 (n_31_74) );
AOI211_X1 g_43_69 (.ZN (n_43_69), .A (n_46_68), .B (n_40_71), .C1 (n_36_73), .C2 (n_30_76) );
AOI211_X1 g_45_68 (.ZN (n_45_68), .A (n_45_70), .B (n_42_70), .C1 (n_38_72), .C2 (n_32_75) );
AOI211_X1 g_47_67 (.ZN (n_47_67), .A (n_43_69), .B (n_44_69), .C1 (n_40_71), .C2 (n_34_74) );
AOI211_X1 g_49_66 (.ZN (n_49_66), .A (n_45_68), .B (n_46_68), .C1 (n_42_70), .C2 (n_36_73) );
AOI211_X1 g_51_65 (.ZN (n_51_65), .A (n_47_67), .B (n_45_70), .C1 (n_44_69), .C2 (n_38_72) );
AOI211_X1 g_50_67 (.ZN (n_50_67), .A (n_49_66), .B (n_43_69), .C1 (n_46_68), .C2 (n_40_71) );
AOI211_X1 g_52_66 (.ZN (n_52_66), .A (n_51_65), .B (n_45_68), .C1 (n_45_70), .C2 (n_42_70) );
AOI211_X1 g_54_65 (.ZN (n_54_65), .A (n_50_67), .B (n_47_67), .C1 (n_43_69), .C2 (n_44_69) );
AOI211_X1 g_56_64 (.ZN (n_56_64), .A (n_52_66), .B (n_49_66), .C1 (n_45_68), .C2 (n_46_68) );
AOI211_X1 g_58_63 (.ZN (n_58_63), .A (n_54_65), .B (n_51_65), .C1 (n_47_67), .C2 (n_45_70) );
AOI211_X1 g_57_65 (.ZN (n_57_65), .A (n_56_64), .B (n_50_67), .C1 (n_49_66), .C2 (n_43_69) );
AOI211_X1 g_55_64 (.ZN (n_55_64), .A (n_58_63), .B (n_52_66), .C1 (n_51_65), .C2 (n_45_68) );
AOI211_X1 g_57_63 (.ZN (n_57_63), .A (n_57_65), .B (n_54_65), .C1 (n_50_67), .C2 (n_47_67) );
AOI211_X1 g_59_62 (.ZN (n_59_62), .A (n_55_64), .B (n_56_64), .C1 (n_52_66), .C2 (n_49_66) );
AOI211_X1 g_61_61 (.ZN (n_61_61), .A (n_57_63), .B (n_58_63), .C1 (n_54_65), .C2 (n_51_65) );
AOI211_X1 g_63_60 (.ZN (n_63_60), .A (n_59_62), .B (n_57_65), .C1 (n_56_64), .C2 (n_50_67) );
AOI211_X1 g_65_59 (.ZN (n_65_59), .A (n_61_61), .B (n_55_64), .C1 (n_58_63), .C2 (n_52_66) );
AOI211_X1 g_67_58 (.ZN (n_67_58), .A (n_63_60), .B (n_57_63), .C1 (n_57_65), .C2 (n_54_65) );
AOI211_X1 g_69_57 (.ZN (n_69_57), .A (n_65_59), .B (n_59_62), .C1 (n_55_64), .C2 (n_56_64) );
AOI211_X1 g_71_56 (.ZN (n_71_56), .A (n_67_58), .B (n_61_61), .C1 (n_57_63), .C2 (n_58_63) );
AOI211_X1 g_73_55 (.ZN (n_73_55), .A (n_69_57), .B (n_63_60), .C1 (n_59_62), .C2 (n_57_65) );
AOI211_X1 g_75_54 (.ZN (n_75_54), .A (n_71_56), .B (n_65_59), .C1 (n_61_61), .C2 (n_55_64) );
AOI211_X1 g_77_53 (.ZN (n_77_53), .A (n_73_55), .B (n_67_58), .C1 (n_63_60), .C2 (n_57_63) );
AOI211_X1 g_79_52 (.ZN (n_79_52), .A (n_75_54), .B (n_69_57), .C1 (n_65_59), .C2 (n_59_62) );
AOI211_X1 g_81_51 (.ZN (n_81_51), .A (n_77_53), .B (n_71_56), .C1 (n_67_58), .C2 (n_61_61) );
AOI211_X1 g_83_52 (.ZN (n_83_52), .A (n_79_52), .B (n_73_55), .C1 (n_69_57), .C2 (n_63_60) );
AOI211_X1 g_81_53 (.ZN (n_81_53), .A (n_81_51), .B (n_75_54), .C1 (n_71_56), .C2 (n_65_59) );
AOI211_X1 g_79_54 (.ZN (n_79_54), .A (n_83_52), .B (n_77_53), .C1 (n_73_55), .C2 (n_67_58) );
AOI211_X1 g_80_52 (.ZN (n_80_52), .A (n_81_53), .B (n_79_52), .C1 (n_75_54), .C2 (n_69_57) );
AOI211_X1 g_78_53 (.ZN (n_78_53), .A (n_79_54), .B (n_81_51), .C1 (n_77_53), .C2 (n_71_56) );
AOI211_X1 g_76_54 (.ZN (n_76_54), .A (n_80_52), .B (n_83_52), .C1 (n_79_52), .C2 (n_73_55) );
AOI211_X1 g_74_55 (.ZN (n_74_55), .A (n_78_53), .B (n_81_53), .C1 (n_81_51), .C2 (n_75_54) );
AOI211_X1 g_72_56 (.ZN (n_72_56), .A (n_76_54), .B (n_79_54), .C1 (n_83_52), .C2 (n_77_53) );
AOI211_X1 g_70_57 (.ZN (n_70_57), .A (n_74_55), .B (n_80_52), .C1 (n_81_53), .C2 (n_79_52) );
AOI211_X1 g_69_59 (.ZN (n_69_59), .A (n_72_56), .B (n_78_53), .C1 (n_79_54), .C2 (n_81_51) );
AOI211_X1 g_71_58 (.ZN (n_71_58), .A (n_70_57), .B (n_76_54), .C1 (n_80_52), .C2 (n_83_52) );
AOI211_X1 g_73_57 (.ZN (n_73_57), .A (n_69_59), .B (n_74_55), .C1 (n_78_53), .C2 (n_81_53) );
AOI211_X1 g_75_56 (.ZN (n_75_56), .A (n_71_58), .B (n_72_56), .C1 (n_76_54), .C2 (n_79_54) );
AOI211_X1 g_77_55 (.ZN (n_77_55), .A (n_73_57), .B (n_70_57), .C1 (n_74_55), .C2 (n_80_52) );
AOI211_X1 g_76_57 (.ZN (n_76_57), .A (n_75_56), .B (n_69_59), .C1 (n_72_56), .C2 (n_78_53) );
AOI211_X1 g_74_56 (.ZN (n_74_56), .A (n_77_55), .B (n_71_58), .C1 (n_70_57), .C2 (n_76_54) );
AOI211_X1 g_76_55 (.ZN (n_76_55), .A (n_76_57), .B (n_73_57), .C1 (n_69_59), .C2 (n_74_55) );
AOI211_X1 g_78_54 (.ZN (n_78_54), .A (n_74_56), .B (n_75_56), .C1 (n_71_58), .C2 (n_72_56) );
AOI211_X1 g_80_53 (.ZN (n_80_53), .A (n_76_55), .B (n_77_55), .C1 (n_73_57), .C2 (n_70_57) );
AOI211_X1 g_82_52 (.ZN (n_82_52), .A (n_78_54), .B (n_76_57), .C1 (n_75_56), .C2 (n_69_59) );
AOI211_X1 g_84_51 (.ZN (n_84_51), .A (n_80_53), .B (n_74_56), .C1 (n_77_55), .C2 (n_71_58) );
AOI211_X1 g_86_50 (.ZN (n_86_50), .A (n_82_52), .B (n_76_55), .C1 (n_76_57), .C2 (n_73_57) );
AOI211_X1 g_88_49 (.ZN (n_88_49), .A (n_84_51), .B (n_78_54), .C1 (n_74_56), .C2 (n_75_56) );
AOI211_X1 g_90_48 (.ZN (n_90_48), .A (n_86_50), .B (n_80_53), .C1 (n_76_55), .C2 (n_77_55) );
AOI211_X1 g_92_47 (.ZN (n_92_47), .A (n_88_49), .B (n_82_52), .C1 (n_78_54), .C2 (n_76_57) );
AOI211_X1 g_94_46 (.ZN (n_94_46), .A (n_90_48), .B (n_84_51), .C1 (n_80_53), .C2 (n_74_56) );
AOI211_X1 g_93_48 (.ZN (n_93_48), .A (n_92_47), .B (n_86_50), .C1 (n_82_52), .C2 (n_76_55) );
AOI211_X1 g_91_49 (.ZN (n_91_49), .A (n_94_46), .B (n_88_49), .C1 (n_84_51), .C2 (n_78_54) );
AOI211_X1 g_89_50 (.ZN (n_89_50), .A (n_93_48), .B (n_90_48), .C1 (n_86_50), .C2 (n_80_53) );
AOI211_X1 g_87_51 (.ZN (n_87_51), .A (n_91_49), .B (n_92_47), .C1 (n_88_49), .C2 (n_82_52) );
AOI211_X1 g_85_52 (.ZN (n_85_52), .A (n_89_50), .B (n_94_46), .C1 (n_90_48), .C2 (n_84_51) );
AOI211_X1 g_83_53 (.ZN (n_83_53), .A (n_87_51), .B (n_93_48), .C1 (n_92_47), .C2 (n_86_50) );
AOI211_X1 g_81_54 (.ZN (n_81_54), .A (n_85_52), .B (n_91_49), .C1 (n_94_46), .C2 (n_88_49) );
AOI211_X1 g_79_55 (.ZN (n_79_55), .A (n_83_53), .B (n_89_50), .C1 (n_93_48), .C2 (n_90_48) );
AOI211_X1 g_77_56 (.ZN (n_77_56), .A (n_81_54), .B (n_87_51), .C1 (n_91_49), .C2 (n_92_47) );
AOI211_X1 g_75_57 (.ZN (n_75_57), .A (n_79_55), .B (n_85_52), .C1 (n_89_50), .C2 (n_94_46) );
AOI211_X1 g_73_58 (.ZN (n_73_58), .A (n_77_56), .B (n_83_53), .C1 (n_87_51), .C2 (n_93_48) );
AOI211_X1 g_71_59 (.ZN (n_71_59), .A (n_75_57), .B (n_81_54), .C1 (n_85_52), .C2 (n_91_49) );
AOI211_X1 g_72_57 (.ZN (n_72_57), .A (n_73_58), .B (n_79_55), .C1 (n_83_53), .C2 (n_89_50) );
AOI211_X1 g_70_58 (.ZN (n_70_58), .A (n_71_59), .B (n_77_56), .C1 (n_81_54), .C2 (n_87_51) );
AOI211_X1 g_68_59 (.ZN (n_68_59), .A (n_72_57), .B (n_75_57), .C1 (n_79_55), .C2 (n_85_52) );
AOI211_X1 g_66_60 (.ZN (n_66_60), .A (n_70_58), .B (n_73_58), .C1 (n_77_56), .C2 (n_83_53) );
AOI211_X1 g_64_61 (.ZN (n_64_61), .A (n_68_59), .B (n_71_59), .C1 (n_75_57), .C2 (n_81_54) );
AOI211_X1 g_62_62 (.ZN (n_62_62), .A (n_66_60), .B (n_72_57), .C1 (n_73_58), .C2 (n_79_55) );
AOI211_X1 g_60_63 (.ZN (n_60_63), .A (n_64_61), .B (n_70_58), .C1 (n_71_59), .C2 (n_77_56) );
AOI211_X1 g_58_64 (.ZN (n_58_64), .A (n_62_62), .B (n_68_59), .C1 (n_72_57), .C2 (n_75_57) );
AOI211_X1 g_56_65 (.ZN (n_56_65), .A (n_60_63), .B (n_66_60), .C1 (n_70_58), .C2 (n_73_58) );
AOI211_X1 g_54_66 (.ZN (n_54_66), .A (n_58_64), .B (n_64_61), .C1 (n_68_59), .C2 (n_71_59) );
AOI211_X1 g_52_67 (.ZN (n_52_67), .A (n_56_65), .B (n_62_62), .C1 (n_66_60), .C2 (n_72_57) );
AOI211_X1 g_53_65 (.ZN (n_53_65), .A (n_54_66), .B (n_60_63), .C1 (n_64_61), .C2 (n_70_58) );
AOI211_X1 g_51_66 (.ZN (n_51_66), .A (n_52_67), .B (n_58_64), .C1 (n_62_62), .C2 (n_68_59) );
AOI211_X1 g_49_67 (.ZN (n_49_67), .A (n_53_65), .B (n_56_65), .C1 (n_60_63), .C2 (n_66_60) );
AOI211_X1 g_47_68 (.ZN (n_47_68), .A (n_51_66), .B (n_54_66), .C1 (n_58_64), .C2 (n_64_61) );
AOI211_X1 g_45_69 (.ZN (n_45_69), .A (n_49_67), .B (n_52_67), .C1 (n_56_65), .C2 (n_62_62) );
AOI211_X1 g_43_70 (.ZN (n_43_70), .A (n_47_68), .B (n_53_65), .C1 (n_54_66), .C2 (n_60_63) );
AOI211_X1 g_41_71 (.ZN (n_41_71), .A (n_45_69), .B (n_51_66), .C1 (n_52_67), .C2 (n_58_64) );
AOI211_X1 g_39_72 (.ZN (n_39_72), .A (n_43_70), .B (n_49_67), .C1 (n_53_65), .C2 (n_56_65) );
AOI211_X1 g_37_73 (.ZN (n_37_73), .A (n_41_71), .B (n_47_68), .C1 (n_51_66), .C2 (n_54_66) );
AOI211_X1 g_35_74 (.ZN (n_35_74), .A (n_39_72), .B (n_45_69), .C1 (n_49_67), .C2 (n_52_67) );
AOI211_X1 g_33_75 (.ZN (n_33_75), .A (n_37_73), .B (n_43_70), .C1 (n_47_68), .C2 (n_53_65) );
AOI211_X1 g_31_76 (.ZN (n_31_76), .A (n_35_74), .B (n_41_71), .C1 (n_45_69), .C2 (n_51_66) );
AOI211_X1 g_29_77 (.ZN (n_29_77), .A (n_33_75), .B (n_39_72), .C1 (n_43_70), .C2 (n_49_67) );
AOI211_X1 g_27_78 (.ZN (n_27_78), .A (n_31_76), .B (n_37_73), .C1 (n_41_71), .C2 (n_47_68) );
AOI211_X1 g_25_79 (.ZN (n_25_79), .A (n_29_77), .B (n_35_74), .C1 (n_39_72), .C2 (n_45_69) );
AOI211_X1 g_26_77 (.ZN (n_26_77), .A (n_27_78), .B (n_33_75), .C1 (n_37_73), .C2 (n_43_70) );
AOI211_X1 g_24_78 (.ZN (n_24_78), .A (n_25_79), .B (n_31_76), .C1 (n_35_74), .C2 (n_41_71) );
AOI211_X1 g_22_79 (.ZN (n_22_79), .A (n_26_77), .B (n_29_77), .C1 (n_33_75), .C2 (n_39_72) );
AOI211_X1 g_20_80 (.ZN (n_20_80), .A (n_24_78), .B (n_27_78), .C1 (n_31_76), .C2 (n_37_73) );
AOI211_X1 g_18_81 (.ZN (n_18_81), .A (n_22_79), .B (n_25_79), .C1 (n_29_77), .C2 (n_35_74) );
AOI211_X1 g_16_82 (.ZN (n_16_82), .A (n_20_80), .B (n_26_77), .C1 (n_27_78), .C2 (n_33_75) );
AOI211_X1 g_14_83 (.ZN (n_14_83), .A (n_18_81), .B (n_24_78), .C1 (n_25_79), .C2 (n_31_76) );
AOI211_X1 g_12_84 (.ZN (n_12_84), .A (n_16_82), .B (n_22_79), .C1 (n_26_77), .C2 (n_29_77) );
AOI211_X1 g_10_83 (.ZN (n_10_83), .A (n_14_83), .B (n_20_80), .C1 (n_24_78), .C2 (n_27_78) );
AOI211_X1 g_8_82 (.ZN (n_8_82), .A (n_12_84), .B (n_18_81), .C1 (n_22_79), .C2 (n_25_79) );
AOI211_X1 g_10_81 (.ZN (n_10_81), .A (n_10_83), .B (n_16_82), .C1 (n_20_80), .C2 (n_26_77) );
AOI211_X1 g_9_83 (.ZN (n_9_83), .A (n_8_82), .B (n_14_83), .C1 (n_18_81), .C2 (n_24_78) );
AOI211_X1 g_7_84 (.ZN (n_7_84), .A (n_10_81), .B (n_12_84), .C1 (n_16_82), .C2 (n_22_79) );
AOI211_X1 g_6_86 (.ZN (n_6_86), .A (n_9_83), .B (n_10_83), .C1 (n_14_83), .C2 (n_20_80) );
AOI211_X1 g_8_85 (.ZN (n_8_85), .A (n_7_84), .B (n_8_82), .C1 (n_12_84), .C2 (n_18_81) );
AOI211_X1 g_7_87 (.ZN (n_7_87), .A (n_6_86), .B (n_10_81), .C1 (n_10_83), .C2 (n_16_82) );
AOI211_X1 g_5_88 (.ZN (n_5_88), .A (n_8_85), .B (n_9_83), .C1 (n_8_82), .C2 (n_14_83) );
AOI211_X1 g_4_90 (.ZN (n_4_90), .A (n_7_87), .B (n_7_84), .C1 (n_10_81), .C2 (n_12_84) );
AOI211_X1 g_6_89 (.ZN (n_6_89), .A (n_5_88), .B (n_6_86), .C1 (n_9_83), .C2 (n_10_83) );
AOI211_X1 g_5_91 (.ZN (n_5_91), .A (n_4_90), .B (n_8_85), .C1 (n_7_84), .C2 (n_8_82) );
AOI211_X1 g_3_92 (.ZN (n_3_92), .A (n_6_89), .B (n_7_87), .C1 (n_6_86), .C2 (n_10_81) );
AOI211_X1 g_2_94 (.ZN (n_2_94), .A (n_5_91), .B (n_5_88), .C1 (n_8_85), .C2 (n_9_83) );
AOI211_X1 g_4_93 (.ZN (n_4_93), .A (n_3_92), .B (n_4_90), .C1 (n_7_87), .C2 (n_7_84) );
AOI211_X1 g_3_95 (.ZN (n_3_95), .A (n_2_94), .B (n_6_89), .C1 (n_5_88), .C2 (n_6_86) );
AOI211_X1 g_1_96 (.ZN (n_1_96), .A (n_4_93), .B (n_5_91), .C1 (n_4_90), .C2 (n_8_85) );
AOI211_X1 g_2_98 (.ZN (n_2_98), .A (n_3_95), .B (n_3_92), .C1 (n_6_89), .C2 (n_7_87) );
AOI211_X1 g_1_100 (.ZN (n_1_100), .A (n_1_96), .B (n_2_94), .C1 (n_5_91), .C2 (n_5_88) );
AOI211_X1 g_3_99 (.ZN (n_3_99), .A (n_2_98), .B (n_4_93), .C1 (n_3_92), .C2 (n_4_90) );
AOI211_X1 g_4_97 (.ZN (n_4_97), .A (n_1_100), .B (n_3_95), .C1 (n_2_94), .C2 (n_6_89) );
AOI211_X1 g_5_95 (.ZN (n_5_95), .A (n_3_99), .B (n_1_96), .C1 (n_4_93), .C2 (n_5_91) );
AOI211_X1 g_3_96 (.ZN (n_3_96), .A (n_4_97), .B (n_2_98), .C1 (n_3_95), .C2 (n_3_92) );
AOI211_X1 g_4_94 (.ZN (n_4_94), .A (n_5_95), .B (n_1_100), .C1 (n_1_96), .C2 (n_2_94) );
AOI211_X1 g_6_93 (.ZN (n_6_93), .A (n_3_96), .B (n_3_99), .C1 (n_2_98), .C2 (n_4_93) );
AOI211_X1 g_7_91 (.ZN (n_7_91), .A (n_4_94), .B (n_4_97), .C1 (n_1_100), .C2 (n_3_95) );
AOI211_X1 g_5_92 (.ZN (n_5_92), .A (n_6_93), .B (n_5_95), .C1 (n_3_99), .C2 (n_1_96) );
AOI211_X1 g_6_90 (.ZN (n_6_90), .A (n_7_91), .B (n_3_96), .C1 (n_4_97), .C2 (n_2_98) );
AOI211_X1 g_8_89 (.ZN (n_8_89), .A (n_5_92), .B (n_4_94), .C1 (n_5_95), .C2 (n_1_100) );
AOI211_X1 g_9_87 (.ZN (n_9_87), .A (n_6_90), .B (n_6_93), .C1 (n_3_96), .C2 (n_3_99) );
AOI211_X1 g_7_88 (.ZN (n_7_88), .A (n_8_89), .B (n_7_91), .C1 (n_4_94), .C2 (n_4_97) );
AOI211_X1 g_8_86 (.ZN (n_8_86), .A (n_9_87), .B (n_5_92), .C1 (n_6_93), .C2 (n_5_95) );
AOI211_X1 g_10_85 (.ZN (n_10_85), .A (n_7_88), .B (n_6_90), .C1 (n_7_91), .C2 (n_3_96) );
AOI211_X1 g_11_83 (.ZN (n_11_83), .A (n_8_86), .B (n_8_89), .C1 (n_5_92), .C2 (n_4_94) );
AOI211_X1 g_9_84 (.ZN (n_9_84), .A (n_10_85), .B (n_9_87), .C1 (n_6_90), .C2 (n_6_93) );
AOI211_X1 g_11_85 (.ZN (n_11_85), .A (n_11_83), .B (n_7_88), .C1 (n_8_89), .C2 (n_7_91) );
AOI211_X1 g_13_84 (.ZN (n_13_84), .A (n_9_84), .B (n_8_86), .C1 (n_9_87), .C2 (n_5_92) );
AOI211_X1 g_15_83 (.ZN (n_15_83), .A (n_11_85), .B (n_10_85), .C1 (n_7_88), .C2 (n_6_90) );
AOI211_X1 g_17_82 (.ZN (n_17_82), .A (n_13_84), .B (n_11_83), .C1 (n_8_86), .C2 (n_8_89) );
AOI211_X1 g_19_81 (.ZN (n_19_81), .A (n_15_83), .B (n_9_84), .C1 (n_10_85), .C2 (n_9_87) );
AOI211_X1 g_21_80 (.ZN (n_21_80), .A (n_17_82), .B (n_11_85), .C1 (n_11_83), .C2 (n_7_88) );
AOI211_X1 g_23_79 (.ZN (n_23_79), .A (n_19_81), .B (n_13_84), .C1 (n_9_84), .C2 (n_8_86) );
AOI211_X1 g_25_78 (.ZN (n_25_78), .A (n_21_80), .B (n_15_83), .C1 (n_11_85), .C2 (n_10_85) );
AOI211_X1 g_27_77 (.ZN (n_27_77), .A (n_23_79), .B (n_17_82), .C1 (n_13_84), .C2 (n_11_83) );
AOI211_X1 g_26_79 (.ZN (n_26_79), .A (n_25_78), .B (n_19_81), .C1 (n_15_83), .C2 (n_9_84) );
AOI211_X1 g_28_78 (.ZN (n_28_78), .A (n_27_77), .B (n_21_80), .C1 (n_17_82), .C2 (n_11_85) );
AOI211_X1 g_30_77 (.ZN (n_30_77), .A (n_26_79), .B (n_23_79), .C1 (n_19_81), .C2 (n_13_84) );
AOI211_X1 g_31_75 (.ZN (n_31_75), .A (n_28_78), .B (n_25_78), .C1 (n_21_80), .C2 (n_15_83) );
AOI211_X1 g_33_74 (.ZN (n_33_74), .A (n_30_77), .B (n_27_77), .C1 (n_23_79), .C2 (n_17_82) );
AOI211_X1 g_35_73 (.ZN (n_35_73), .A (n_31_75), .B (n_26_79), .C1 (n_25_78), .C2 (n_19_81) );
AOI211_X1 g_37_72 (.ZN (n_37_72), .A (n_33_74), .B (n_28_78), .C1 (n_27_77), .C2 (n_21_80) );
AOI211_X1 g_39_71 (.ZN (n_39_71), .A (n_35_73), .B (n_30_77), .C1 (n_26_79), .C2 (n_23_79) );
AOI211_X1 g_41_70 (.ZN (n_41_70), .A (n_37_72), .B (n_31_75), .C1 (n_28_78), .C2 (n_25_78) );
AOI211_X1 g_43_71 (.ZN (n_43_71), .A (n_39_71), .B (n_33_74), .C1 (n_30_77), .C2 (n_27_77) );
AOI211_X1 g_41_72 (.ZN (n_41_72), .A (n_41_70), .B (n_35_73), .C1 (n_31_75), .C2 (n_26_79) );
AOI211_X1 g_39_73 (.ZN (n_39_73), .A (n_43_71), .B (n_37_72), .C1 (n_33_74), .C2 (n_28_78) );
AOI211_X1 g_37_74 (.ZN (n_37_74), .A (n_41_72), .B (n_39_71), .C1 (n_35_73), .C2 (n_30_77) );
AOI211_X1 g_35_75 (.ZN (n_35_75), .A (n_39_73), .B (n_41_70), .C1 (n_37_72), .C2 (n_31_75) );
AOI211_X1 g_33_76 (.ZN (n_33_76), .A (n_37_74), .B (n_43_71), .C1 (n_39_71), .C2 (n_33_74) );
AOI211_X1 g_31_77 (.ZN (n_31_77), .A (n_35_75), .B (n_41_72), .C1 (n_41_70), .C2 (n_35_73) );
AOI211_X1 g_29_78 (.ZN (n_29_78), .A (n_33_76), .B (n_39_73), .C1 (n_43_71), .C2 (n_37_72) );
AOI211_X1 g_27_79 (.ZN (n_27_79), .A (n_31_77), .B (n_37_74), .C1 (n_41_72), .C2 (n_39_71) );
AOI211_X1 g_28_77 (.ZN (n_28_77), .A (n_29_78), .B (n_35_75), .C1 (n_39_73), .C2 (n_41_70) );
AOI211_X1 g_26_78 (.ZN (n_26_78), .A (n_27_79), .B (n_33_76), .C1 (n_37_74), .C2 (n_43_71) );
AOI211_X1 g_24_79 (.ZN (n_24_79), .A (n_28_77), .B (n_31_77), .C1 (n_35_75), .C2 (n_41_72) );
AOI211_X1 g_22_80 (.ZN (n_22_80), .A (n_26_78), .B (n_29_78), .C1 (n_33_76), .C2 (n_39_73) );
AOI211_X1 g_20_81 (.ZN (n_20_81), .A (n_24_79), .B (n_27_79), .C1 (n_31_77), .C2 (n_37_74) );
AOI211_X1 g_18_82 (.ZN (n_18_82), .A (n_22_80), .B (n_28_77), .C1 (n_29_78), .C2 (n_35_75) );
AOI211_X1 g_16_83 (.ZN (n_16_83), .A (n_20_81), .B (n_26_78), .C1 (n_27_79), .C2 (n_33_76) );
AOI211_X1 g_17_81 (.ZN (n_17_81), .A (n_18_82), .B (n_24_79), .C1 (n_28_77), .C2 (n_31_77) );
AOI211_X1 g_15_82 (.ZN (n_15_82), .A (n_16_83), .B (n_22_80), .C1 (n_26_78), .C2 (n_29_78) );
AOI211_X1 g_13_83 (.ZN (n_13_83), .A (n_17_81), .B (n_20_81), .C1 (n_24_79), .C2 (n_27_79) );
AOI211_X1 g_11_84 (.ZN (n_11_84), .A (n_15_82), .B (n_18_82), .C1 (n_22_80), .C2 (n_28_77) );
AOI211_X1 g_9_85 (.ZN (n_9_85), .A (n_13_83), .B (n_16_83), .C1 (n_20_81), .C2 (n_26_78) );
AOI211_X1 g_8_87 (.ZN (n_8_87), .A (n_11_84), .B (n_17_81), .C1 (n_18_82), .C2 (n_24_79) );
AOI211_X1 g_10_86 (.ZN (n_10_86), .A (n_9_85), .B (n_15_82), .C1 (n_16_83), .C2 (n_22_80) );
AOI211_X1 g_12_85 (.ZN (n_12_85), .A (n_8_87), .B (n_13_83), .C1 (n_17_81), .C2 (n_20_81) );
AOI211_X1 g_14_84 (.ZN (n_14_84), .A (n_10_86), .B (n_11_84), .C1 (n_15_82), .C2 (n_18_82) );
AOI211_X1 g_13_86 (.ZN (n_13_86), .A (n_12_85), .B (n_9_85), .C1 (n_13_83), .C2 (n_16_83) );
AOI211_X1 g_15_85 (.ZN (n_15_85), .A (n_14_84), .B (n_8_87), .C1 (n_11_84), .C2 (n_17_81) );
AOI211_X1 g_17_84 (.ZN (n_17_84), .A (n_13_86), .B (n_10_86), .C1 (n_9_85), .C2 (n_15_82) );
AOI211_X1 g_19_83 (.ZN (n_19_83), .A (n_15_85), .B (n_12_85), .C1 (n_8_87), .C2 (n_13_83) );
AOI211_X1 g_21_82 (.ZN (n_21_82), .A (n_17_84), .B (n_14_84), .C1 (n_10_86), .C2 (n_11_84) );
AOI211_X1 g_23_81 (.ZN (n_23_81), .A (n_19_83), .B (n_13_86), .C1 (n_12_85), .C2 (n_9_85) );
AOI211_X1 g_25_80 (.ZN (n_25_80), .A (n_21_82), .B (n_15_85), .C1 (n_14_84), .C2 (n_8_87) );
AOI211_X1 g_27_81 (.ZN (n_27_81), .A (n_23_81), .B (n_17_84), .C1 (n_13_86), .C2 (n_10_86) );
AOI211_X1 g_28_79 (.ZN (n_28_79), .A (n_25_80), .B (n_19_83), .C1 (n_15_85), .C2 (n_12_85) );
AOI211_X1 g_30_78 (.ZN (n_30_78), .A (n_27_81), .B (n_21_82), .C1 (n_17_84), .C2 (n_14_84) );
AOI211_X1 g_32_77 (.ZN (n_32_77), .A (n_28_79), .B (n_23_81), .C1 (n_19_83), .C2 (n_13_86) );
AOI211_X1 g_34_76 (.ZN (n_34_76), .A (n_30_78), .B (n_25_80), .C1 (n_21_82), .C2 (n_15_85) );
AOI211_X1 g_36_75 (.ZN (n_36_75), .A (n_32_77), .B (n_27_81), .C1 (n_23_81), .C2 (n_17_84) );
AOI211_X1 g_38_74 (.ZN (n_38_74), .A (n_34_76), .B (n_28_79), .C1 (n_25_80), .C2 (n_19_83) );
AOI211_X1 g_40_73 (.ZN (n_40_73), .A (n_36_75), .B (n_30_78), .C1 (n_27_81), .C2 (n_21_82) );
AOI211_X1 g_42_72 (.ZN (n_42_72), .A (n_38_74), .B (n_32_77), .C1 (n_28_79), .C2 (n_23_81) );
AOI211_X1 g_44_71 (.ZN (n_44_71), .A (n_40_73), .B (n_34_76), .C1 (n_30_78), .C2 (n_25_80) );
AOI211_X1 g_46_70 (.ZN (n_46_70), .A (n_42_72), .B (n_36_75), .C1 (n_32_77), .C2 (n_27_81) );
AOI211_X1 g_48_69 (.ZN (n_48_69), .A (n_44_71), .B (n_38_74), .C1 (n_34_76), .C2 (n_28_79) );
AOI211_X1 g_50_68 (.ZN (n_50_68), .A (n_46_70), .B (n_40_73), .C1 (n_36_75), .C2 (n_30_78) );
AOI211_X1 g_49_70 (.ZN (n_49_70), .A (n_48_69), .B (n_42_72), .C1 (n_38_74), .C2 (n_32_77) );
AOI211_X1 g_48_68 (.ZN (n_48_68), .A (n_50_68), .B (n_44_71), .C1 (n_40_73), .C2 (n_34_76) );
AOI211_X1 g_46_69 (.ZN (n_46_69), .A (n_49_70), .B (n_46_70), .C1 (n_42_72), .C2 (n_36_75) );
AOI211_X1 g_44_70 (.ZN (n_44_70), .A (n_48_68), .B (n_48_69), .C1 (n_44_71), .C2 (n_38_74) );
AOI211_X1 g_42_71 (.ZN (n_42_71), .A (n_46_69), .B (n_50_68), .C1 (n_46_70), .C2 (n_40_73) );
AOI211_X1 g_40_72 (.ZN (n_40_72), .A (n_44_70), .B (n_49_70), .C1 (n_48_69), .C2 (n_42_72) );
AOI211_X1 g_38_73 (.ZN (n_38_73), .A (n_42_71), .B (n_48_68), .C1 (n_50_68), .C2 (n_44_71) );
AOI211_X1 g_36_74 (.ZN (n_36_74), .A (n_40_72), .B (n_46_69), .C1 (n_49_70), .C2 (n_46_70) );
AOI211_X1 g_34_75 (.ZN (n_34_75), .A (n_38_73), .B (n_44_70), .C1 (n_48_68), .C2 (n_48_69) );
AOI211_X1 g_32_76 (.ZN (n_32_76), .A (n_36_74), .B (n_42_71), .C1 (n_46_69), .C2 (n_50_68) );
AOI211_X1 g_31_78 (.ZN (n_31_78), .A (n_34_75), .B (n_40_72), .C1 (n_44_70), .C2 (n_49_70) );
AOI211_X1 g_33_77 (.ZN (n_33_77), .A (n_32_76), .B (n_38_73), .C1 (n_42_71), .C2 (n_48_68) );
AOI211_X1 g_35_76 (.ZN (n_35_76), .A (n_31_78), .B (n_36_74), .C1 (n_40_72), .C2 (n_46_69) );
AOI211_X1 g_37_75 (.ZN (n_37_75), .A (n_33_77), .B (n_34_75), .C1 (n_38_73), .C2 (n_44_70) );
AOI211_X1 g_39_74 (.ZN (n_39_74), .A (n_35_76), .B (n_32_76), .C1 (n_36_74), .C2 (n_42_71) );
AOI211_X1 g_41_73 (.ZN (n_41_73), .A (n_37_75), .B (n_31_78), .C1 (n_34_75), .C2 (n_40_72) );
AOI211_X1 g_43_72 (.ZN (n_43_72), .A (n_39_74), .B (n_33_77), .C1 (n_32_76), .C2 (n_38_73) );
AOI211_X1 g_45_71 (.ZN (n_45_71), .A (n_41_73), .B (n_35_76), .C1 (n_31_78), .C2 (n_36_74) );
AOI211_X1 g_47_70 (.ZN (n_47_70), .A (n_43_72), .B (n_37_75), .C1 (n_33_77), .C2 (n_34_75) );
AOI211_X1 g_49_69 (.ZN (n_49_69), .A (n_45_71), .B (n_39_74), .C1 (n_35_76), .C2 (n_32_76) );
AOI211_X1 g_51_68 (.ZN (n_51_68), .A (n_47_70), .B (n_41_73), .C1 (n_37_75), .C2 (n_31_78) );
AOI211_X1 g_53_67 (.ZN (n_53_67), .A (n_49_69), .B (n_43_72), .C1 (n_39_74), .C2 (n_33_77) );
AOI211_X1 g_55_66 (.ZN (n_55_66), .A (n_51_68), .B (n_45_71), .C1 (n_41_73), .C2 (n_35_76) );
AOI211_X1 g_54_68 (.ZN (n_54_68), .A (n_53_67), .B (n_47_70), .C1 (n_43_72), .C2 (n_37_75) );
AOI211_X1 g_56_67 (.ZN (n_56_67), .A (n_55_66), .B (n_49_69), .C1 (n_45_71), .C2 (n_39_74) );
AOI211_X1 g_58_66 (.ZN (n_58_66), .A (n_54_68), .B (n_51_68), .C1 (n_47_70), .C2 (n_41_73) );
AOI211_X1 g_59_64 (.ZN (n_59_64), .A (n_56_67), .B (n_53_67), .C1 (n_49_69), .C2 (n_43_72) );
AOI211_X1 g_61_63 (.ZN (n_61_63), .A (n_58_66), .B (n_55_66), .C1 (n_51_68), .C2 (n_45_71) );
AOI211_X1 g_63_62 (.ZN (n_63_62), .A (n_59_64), .B (n_54_68), .C1 (n_53_67), .C2 (n_47_70) );
AOI211_X1 g_65_61 (.ZN (n_65_61), .A (n_61_63), .B (n_56_67), .C1 (n_55_66), .C2 (n_49_69) );
AOI211_X1 g_67_60 (.ZN (n_67_60), .A (n_63_62), .B (n_58_66), .C1 (n_54_68), .C2 (n_51_68) );
AOI211_X1 g_66_62 (.ZN (n_66_62), .A (n_65_61), .B (n_59_64), .C1 (n_56_67), .C2 (n_53_67) );
AOI211_X1 g_68_61 (.ZN (n_68_61), .A (n_67_60), .B (n_61_63), .C1 (n_58_66), .C2 (n_55_66) );
AOI211_X1 g_70_60 (.ZN (n_70_60), .A (n_66_62), .B (n_63_62), .C1 (n_59_64), .C2 (n_54_68) );
AOI211_X1 g_72_59 (.ZN (n_72_59), .A (n_68_61), .B (n_65_61), .C1 (n_61_63), .C2 (n_56_67) );
AOI211_X1 g_74_58 (.ZN (n_74_58), .A (n_70_60), .B (n_67_60), .C1 (n_63_62), .C2 (n_58_66) );
AOI211_X1 g_73_60 (.ZN (n_73_60), .A (n_72_59), .B (n_66_62), .C1 (n_65_61), .C2 (n_59_64) );
AOI211_X1 g_72_58 (.ZN (n_72_58), .A (n_74_58), .B (n_68_61), .C1 (n_67_60), .C2 (n_61_63) );
AOI211_X1 g_70_59 (.ZN (n_70_59), .A (n_73_60), .B (n_70_60), .C1 (n_66_62), .C2 (n_63_62) );
AOI211_X1 g_69_61 (.ZN (n_69_61), .A (n_72_58), .B (n_72_59), .C1 (n_68_61), .C2 (n_65_61) );
AOI211_X1 g_71_60 (.ZN (n_71_60), .A (n_70_59), .B (n_74_58), .C1 (n_70_60), .C2 (n_67_60) );
AOI211_X1 g_73_59 (.ZN (n_73_59), .A (n_69_61), .B (n_73_60), .C1 (n_72_59), .C2 (n_66_62) );
AOI211_X1 g_74_57 (.ZN (n_74_57), .A (n_71_60), .B (n_72_58), .C1 (n_74_58), .C2 (n_68_61) );
AOI211_X1 g_76_56 (.ZN (n_76_56), .A (n_73_59), .B (n_70_59), .C1 (n_73_60), .C2 (n_70_60) );
AOI211_X1 g_78_55 (.ZN (n_78_55), .A (n_74_57), .B (n_69_61), .C1 (n_72_58), .C2 (n_72_59) );
AOI211_X1 g_80_54 (.ZN (n_80_54), .A (n_76_56), .B (n_71_60), .C1 (n_70_59), .C2 (n_74_58) );
AOI211_X1 g_82_53 (.ZN (n_82_53), .A (n_78_55), .B (n_73_59), .C1 (n_69_61), .C2 (n_73_60) );
AOI211_X1 g_81_55 (.ZN (n_81_55), .A (n_80_54), .B (n_74_57), .C1 (n_71_60), .C2 (n_72_58) );
AOI211_X1 g_83_54 (.ZN (n_83_54), .A (n_82_53), .B (n_76_56), .C1 (n_73_59), .C2 (n_70_59) );
AOI211_X1 g_85_53 (.ZN (n_85_53), .A (n_81_55), .B (n_78_55), .C1 (n_74_57), .C2 (n_69_61) );
AOI211_X1 g_86_51 (.ZN (n_86_51), .A (n_83_54), .B (n_80_54), .C1 (n_76_56), .C2 (n_71_60) );
AOI211_X1 g_88_50 (.ZN (n_88_50), .A (n_85_53), .B (n_82_53), .C1 (n_78_55), .C2 (n_73_59) );
AOI211_X1 g_87_52 (.ZN (n_87_52), .A (n_86_51), .B (n_81_55), .C1 (n_80_54), .C2 (n_74_57) );
AOI211_X1 g_89_51 (.ZN (n_89_51), .A (n_88_50), .B (n_83_54), .C1 (n_82_53), .C2 (n_76_56) );
AOI211_X1 g_91_50 (.ZN (n_91_50), .A (n_87_52), .B (n_85_53), .C1 (n_81_55), .C2 (n_78_55) );
AOI211_X1 g_93_49 (.ZN (n_93_49), .A (n_89_51), .B (n_86_51), .C1 (n_83_54), .C2 (n_80_54) );
AOI211_X1 g_95_48 (.ZN (n_95_48), .A (n_91_50), .B (n_88_50), .C1 (n_85_53), .C2 (n_82_53) );
AOI211_X1 g_97_49 (.ZN (n_97_49), .A (n_93_49), .B (n_87_52), .C1 (n_86_51), .C2 (n_81_55) );
AOI211_X1 g_96_47 (.ZN (n_96_47), .A (n_95_48), .B (n_89_51), .C1 (n_88_50), .C2 (n_83_54) );
AOI211_X1 g_94_48 (.ZN (n_94_48), .A (n_97_49), .B (n_91_50), .C1 (n_87_52), .C2 (n_85_53) );
AOI211_X1 g_95_50 (.ZN (n_95_50), .A (n_96_47), .B (n_93_49), .C1 (n_89_51), .C2 (n_86_51) );
AOI211_X1 g_96_52 (.ZN (n_96_52), .A (n_94_48), .B (n_95_48), .C1 (n_91_50), .C2 (n_88_50) );
AOI211_X1 g_94_51 (.ZN (n_94_51), .A (n_95_50), .B (n_97_49), .C1 (n_93_49), .C2 (n_87_52) );
AOI211_X1 g_95_49 (.ZN (n_95_49), .A (n_96_52), .B (n_96_47), .C1 (n_95_48), .C2 (n_89_51) );
AOI211_X1 g_93_50 (.ZN (n_93_50), .A (n_94_51), .B (n_94_48), .C1 (n_97_49), .C2 (n_91_50) );
AOI211_X1 g_95_51 (.ZN (n_95_51), .A (n_95_49), .B (n_95_50), .C1 (n_96_47), .C2 (n_93_49) );
AOI211_X1 g_96_53 (.ZN (n_96_53), .A (n_93_50), .B (n_96_52), .C1 (n_94_48), .C2 (n_95_48) );
AOI211_X1 g_97_55 (.ZN (n_97_55), .A (n_95_51), .B (n_94_51), .C1 (n_95_50), .C2 (n_97_49) );
AOI211_X1 g_98_57 (.ZN (n_98_57), .A (n_96_53), .B (n_95_49), .C1 (n_96_52), .C2 (n_96_47) );
AOI211_X1 g_99_59 (.ZN (n_99_59), .A (n_97_55), .B (n_93_50), .C1 (n_94_51), .C2 (n_94_48) );
AOI211_X1 g_100_61 (.ZN (n_100_61), .A (n_98_57), .B (n_95_51), .C1 (n_95_49), .C2 (n_95_50) );
AOI211_X1 g_98_62 (.ZN (n_98_62), .A (n_99_59), .B (n_96_53), .C1 (n_93_50), .C2 (n_96_52) );
AOI211_X1 g_100_63 (.ZN (n_100_63), .A (n_100_61), .B (n_97_55), .C1 (n_95_51), .C2 (n_94_51) );
AOI211_X1 g_99_61 (.ZN (n_99_61), .A (n_98_62), .B (n_98_57), .C1 (n_96_53), .C2 (n_95_49) );
AOI211_X1 g_97_60 (.ZN (n_97_60), .A (n_100_63), .B (n_99_59), .C1 (n_97_55), .C2 (n_93_50) );
AOI211_X1 g_96_58 (.ZN (n_96_58), .A (n_99_61), .B (n_100_61), .C1 (n_98_57), .C2 (n_95_51) );
AOI211_X1 g_98_59 (.ZN (n_98_59), .A (n_97_60), .B (n_98_62), .C1 (n_99_59), .C2 (n_96_53) );
AOI211_X1 g_100_60 (.ZN (n_100_60), .A (n_96_58), .B (n_100_63), .C1 (n_100_61), .C2 (n_97_55) );
AOI211_X1 g_99_58 (.ZN (n_99_58), .A (n_98_59), .B (n_99_61), .C1 (n_98_62), .C2 (n_98_57) );
AOI211_X1 g_98_56 (.ZN (n_98_56), .A (n_100_60), .B (n_97_60), .C1 (n_100_63), .C2 (n_99_59) );
AOI211_X1 g_97_54 (.ZN (n_97_54), .A (n_99_58), .B (n_96_58), .C1 (n_99_61), .C2 (n_100_61) );
AOI211_X1 g_95_53 (.ZN (n_95_53), .A (n_98_56), .B (n_98_59), .C1 (n_97_60), .C2 (n_98_62) );
AOI211_X1 g_96_51 (.ZN (n_96_51), .A (n_97_54), .B (n_100_60), .C1 (n_96_58), .C2 (n_100_63) );
AOI211_X1 g_97_53 (.ZN (n_97_53), .A (n_95_53), .B (n_99_58), .C1 (n_98_59), .C2 (n_99_61) );
AOI211_X1 g_95_52 (.ZN (n_95_52), .A (n_96_51), .B (n_98_56), .C1 (n_100_60), .C2 (n_97_60) );
AOI211_X1 g_94_50 (.ZN (n_94_50), .A (n_97_53), .B (n_97_54), .C1 (n_99_58), .C2 (n_96_58) );
AOI211_X1 g_92_49 (.ZN (n_92_49), .A (n_95_52), .B (n_95_53), .C1 (n_98_56), .C2 (n_98_59) );
AOI211_X1 g_93_51 (.ZN (n_93_51), .A (n_94_50), .B (n_96_51), .C1 (n_97_54), .C2 (n_100_60) );
AOI211_X1 g_94_53 (.ZN (n_94_53), .A (n_92_49), .B (n_97_53), .C1 (n_95_53), .C2 (n_99_58) );
AOI211_X1 g_92_52 (.ZN (n_92_52), .A (n_93_51), .B (n_95_52), .C1 (n_96_51), .C2 (n_98_56) );
AOI211_X1 g_90_51 (.ZN (n_90_51), .A (n_94_53), .B (n_94_50), .C1 (n_97_53), .C2 (n_97_54) );
AOI211_X1 g_88_52 (.ZN (n_88_52), .A (n_92_52), .B (n_92_49), .C1 (n_95_52), .C2 (n_95_53) );
AOI211_X1 g_86_53 (.ZN (n_86_53), .A (n_90_51), .B (n_93_51), .C1 (n_94_50), .C2 (n_96_51) );
AOI211_X1 g_84_54 (.ZN (n_84_54), .A (n_88_52), .B (n_94_53), .C1 (n_92_49), .C2 (n_97_53) );
AOI211_X1 g_82_55 (.ZN (n_82_55), .A (n_86_53), .B (n_92_52), .C1 (n_93_51), .C2 (n_95_52) );
AOI211_X1 g_80_56 (.ZN (n_80_56), .A (n_84_54), .B (n_90_51), .C1 (n_94_53), .C2 (n_94_50) );
AOI211_X1 g_78_57 (.ZN (n_78_57), .A (n_82_55), .B (n_88_52), .C1 (n_92_52), .C2 (n_92_49) );
AOI211_X1 g_76_58 (.ZN (n_76_58), .A (n_80_56), .B (n_86_53), .C1 (n_90_51), .C2 (n_93_51) );
AOI211_X1 g_74_59 (.ZN (n_74_59), .A (n_78_57), .B (n_84_54), .C1 (n_88_52), .C2 (n_94_53) );
AOI211_X1 g_72_60 (.ZN (n_72_60), .A (n_76_58), .B (n_82_55), .C1 (n_86_53), .C2 (n_92_52) );
AOI211_X1 g_70_61 (.ZN (n_70_61), .A (n_74_59), .B (n_80_56), .C1 (n_84_54), .C2 (n_90_51) );
AOI211_X1 g_72_62 (.ZN (n_72_62), .A (n_72_60), .B (n_78_57), .C1 (n_82_55), .C2 (n_88_52) );
AOI211_X1 g_74_61 (.ZN (n_74_61), .A (n_70_61), .B (n_76_58), .C1 (n_80_56), .C2 (n_86_53) );
AOI211_X1 g_75_59 (.ZN (n_75_59), .A (n_72_62), .B (n_74_59), .C1 (n_78_57), .C2 (n_84_54) );
AOI211_X1 g_77_58 (.ZN (n_77_58), .A (n_74_61), .B (n_72_60), .C1 (n_76_58), .C2 (n_82_55) );
AOI211_X1 g_78_56 (.ZN (n_78_56), .A (n_75_59), .B (n_70_61), .C1 (n_74_59), .C2 (n_80_56) );
AOI211_X1 g_80_55 (.ZN (n_80_55), .A (n_77_58), .B (n_72_62), .C1 (n_72_60), .C2 (n_78_57) );
AOI211_X1 g_82_54 (.ZN (n_82_54), .A (n_78_56), .B (n_74_61), .C1 (n_70_61), .C2 (n_76_58) );
AOI211_X1 g_84_53 (.ZN (n_84_53), .A (n_80_55), .B (n_75_59), .C1 (n_72_62), .C2 (n_74_59) );
AOI211_X1 g_86_52 (.ZN (n_86_52), .A (n_82_54), .B (n_77_58), .C1 (n_74_61), .C2 (n_72_60) );
AOI211_X1 g_88_51 (.ZN (n_88_51), .A (n_84_53), .B (n_78_56), .C1 (n_75_59), .C2 (n_70_61) );
AOI211_X1 g_90_50 (.ZN (n_90_50), .A (n_86_52), .B (n_80_55), .C1 (n_77_58), .C2 (n_72_62) );
AOI211_X1 g_91_52 (.ZN (n_91_52), .A (n_88_51), .B (n_82_54), .C1 (n_78_56), .C2 (n_74_61) );
AOI211_X1 g_89_53 (.ZN (n_89_53), .A (n_90_50), .B (n_84_53), .C1 (n_80_55), .C2 (n_75_59) );
AOI211_X1 g_87_54 (.ZN (n_87_54), .A (n_91_52), .B (n_86_52), .C1 (n_82_54), .C2 (n_77_58) );
AOI211_X1 g_85_55 (.ZN (n_85_55), .A (n_89_53), .B (n_88_51), .C1 (n_84_53), .C2 (n_78_56) );
AOI211_X1 g_83_56 (.ZN (n_83_56), .A (n_87_54), .B (n_90_50), .C1 (n_86_52), .C2 (n_80_55) );
AOI211_X1 g_81_57 (.ZN (n_81_57), .A (n_85_55), .B (n_91_52), .C1 (n_88_51), .C2 (n_82_54) );
AOI211_X1 g_79_56 (.ZN (n_79_56), .A (n_83_56), .B (n_89_53), .C1 (n_90_50), .C2 (n_84_53) );
AOI211_X1 g_77_57 (.ZN (n_77_57), .A (n_81_57), .B (n_87_54), .C1 (n_91_52), .C2 (n_86_52) );
AOI211_X1 g_75_58 (.ZN (n_75_58), .A (n_79_56), .B (n_85_55), .C1 (n_89_53), .C2 (n_88_51) );
AOI211_X1 g_76_60 (.ZN (n_76_60), .A (n_77_57), .B (n_83_56), .C1 (n_87_54), .C2 (n_90_50) );
AOI211_X1 g_78_59 (.ZN (n_78_59), .A (n_75_58), .B (n_81_57), .C1 (n_85_55), .C2 (n_91_52) );
AOI211_X1 g_79_57 (.ZN (n_79_57), .A (n_76_60), .B (n_79_56), .C1 (n_83_56), .C2 (n_89_53) );
AOI211_X1 g_81_56 (.ZN (n_81_56), .A (n_78_59), .B (n_77_57), .C1 (n_81_57), .C2 (n_87_54) );
AOI211_X1 g_83_55 (.ZN (n_83_55), .A (n_79_57), .B (n_75_58), .C1 (n_79_56), .C2 (n_85_55) );
AOI211_X1 g_85_54 (.ZN (n_85_54), .A (n_81_56), .B (n_76_60), .C1 (n_77_57), .C2 (n_83_56) );
AOI211_X1 g_87_53 (.ZN (n_87_53), .A (n_83_55), .B (n_78_59), .C1 (n_75_58), .C2 (n_81_57) );
AOI211_X1 g_89_52 (.ZN (n_89_52), .A (n_85_54), .B (n_79_57), .C1 (n_76_60), .C2 (n_79_56) );
AOI211_X1 g_91_51 (.ZN (n_91_51), .A (n_87_53), .B (n_81_56), .C1 (n_78_59), .C2 (n_77_57) );
AOI211_X1 g_93_52 (.ZN (n_93_52), .A (n_89_52), .B (n_83_55), .C1 (n_79_57), .C2 (n_75_58) );
AOI211_X1 g_91_53 (.ZN (n_91_53), .A (n_91_51), .B (n_85_54), .C1 (n_81_56), .C2 (n_76_60) );
AOI211_X1 g_92_51 (.ZN (n_92_51), .A (n_93_52), .B (n_87_53), .C1 (n_83_55), .C2 (n_78_59) );
AOI211_X1 g_94_52 (.ZN (n_94_52), .A (n_91_53), .B (n_89_52), .C1 (n_85_54), .C2 (n_79_57) );
AOI211_X1 g_93_54 (.ZN (n_93_54), .A (n_92_51), .B (n_91_51), .C1 (n_87_53), .C2 (n_81_56) );
AOI211_X1 g_95_55 (.ZN (n_95_55), .A (n_94_52), .B (n_93_52), .C1 (n_89_52), .C2 (n_83_55) );
AOI211_X1 g_96_57 (.ZN (n_96_57), .A (n_93_54), .B (n_91_53), .C1 (n_91_51), .C2 (n_85_54) );
AOI211_X1 g_97_59 (.ZN (n_97_59), .A (n_95_55), .B (n_92_51), .C1 (n_93_52), .C2 (n_87_53) );
AOI211_X1 g_98_61 (.ZN (n_98_61), .A (n_96_57), .B (n_94_52), .C1 (n_91_53), .C2 (n_89_52) );
AOI211_X1 g_99_63 (.ZN (n_99_63), .A (n_97_59), .B (n_93_54), .C1 (n_92_51), .C2 (n_91_51) );
AOI211_X1 g_100_65 (.ZN (n_100_65), .A (n_98_61), .B (n_95_55), .C1 (n_94_52), .C2 (n_93_52) );
AOI211_X1 g_98_66 (.ZN (n_98_66), .A (n_99_63), .B (n_96_57), .C1 (n_93_54), .C2 (n_91_53) );
AOI211_X1 g_100_67 (.ZN (n_100_67), .A (n_100_65), .B (n_97_59), .C1 (n_95_55), .C2 (n_92_51) );
AOI211_X1 g_99_65 (.ZN (n_99_65), .A (n_98_66), .B (n_98_61), .C1 (n_96_57), .C2 (n_94_52) );
AOI211_X1 g_97_64 (.ZN (n_97_64), .A (n_100_67), .B (n_99_63), .C1 (n_97_59), .C2 (n_93_54) );
AOI211_X1 g_96_62 (.ZN (n_96_62), .A (n_99_65), .B (n_100_65), .C1 (n_98_61), .C2 (n_95_55) );
AOI211_X1 g_98_63 (.ZN (n_98_63), .A (n_97_64), .B (n_98_66), .C1 (n_99_63), .C2 (n_96_57) );
AOI211_X1 g_100_64 (.ZN (n_100_64), .A (n_96_62), .B (n_100_67), .C1 (n_100_65), .C2 (n_97_59) );
AOI211_X1 g_99_62 (.ZN (n_99_62), .A (n_98_63), .B (n_99_65), .C1 (n_98_66), .C2 (n_98_61) );
AOI211_X1 g_98_60 (.ZN (n_98_60), .A (n_100_64), .B (n_97_64), .C1 (n_100_67), .C2 (n_99_63) );
AOI211_X1 g_97_58 (.ZN (n_97_58), .A (n_99_62), .B (n_96_62), .C1 (n_99_65), .C2 (n_100_65) );
AOI211_X1 g_96_56 (.ZN (n_96_56), .A (n_98_60), .B (n_98_63), .C1 (n_97_64), .C2 (n_98_66) );
AOI211_X1 g_95_54 (.ZN (n_95_54), .A (n_97_58), .B (n_100_64), .C1 (n_96_62), .C2 (n_100_67) );
AOI211_X1 g_93_53 (.ZN (n_93_53), .A (n_96_56), .B (n_99_62), .C1 (n_98_63), .C2 (n_99_65) );
AOI211_X1 g_94_55 (.ZN (n_94_55), .A (n_95_54), .B (n_98_60), .C1 (n_100_64), .C2 (n_97_64) );
AOI211_X1 g_92_54 (.ZN (n_92_54), .A (n_93_53), .B (n_97_58), .C1 (n_99_62), .C2 (n_96_62) );
AOI211_X1 g_90_53 (.ZN (n_90_53), .A (n_94_55), .B (n_96_56), .C1 (n_98_60), .C2 (n_98_63) );
AOI211_X1 g_88_54 (.ZN (n_88_54), .A (n_92_54), .B (n_95_54), .C1 (n_97_58), .C2 (n_100_64) );
AOI211_X1 g_86_55 (.ZN (n_86_55), .A (n_90_53), .B (n_93_53), .C1 (n_96_56), .C2 (n_99_62) );
AOI211_X1 g_84_56 (.ZN (n_84_56), .A (n_88_54), .B (n_94_55), .C1 (n_95_54), .C2 (n_98_60) );
AOI211_X1 g_82_57 (.ZN (n_82_57), .A (n_86_55), .B (n_92_54), .C1 (n_93_53), .C2 (n_97_58) );
AOI211_X1 g_80_58 (.ZN (n_80_58), .A (n_84_56), .B (n_90_53), .C1 (n_94_55), .C2 (n_96_56) );
AOI211_X1 g_82_59 (.ZN (n_82_59), .A (n_82_57), .B (n_88_54), .C1 (n_92_54), .C2 (n_95_54) );
AOI211_X1 g_84_58 (.ZN (n_84_58), .A (n_80_58), .B (n_86_55), .C1 (n_90_53), .C2 (n_93_53) );
AOI211_X1 g_86_57 (.ZN (n_86_57), .A (n_82_59), .B (n_84_56), .C1 (n_88_54), .C2 (n_94_55) );
AOI211_X1 g_88_56 (.ZN (n_88_56), .A (n_84_58), .B (n_82_57), .C1 (n_86_55), .C2 (n_92_54) );
AOI211_X1 g_90_55 (.ZN (n_90_55), .A (n_86_57), .B (n_80_58), .C1 (n_84_56), .C2 (n_90_53) );
AOI211_X1 g_92_56 (.ZN (n_92_56), .A (n_88_56), .B (n_82_59), .C1 (n_82_57), .C2 (n_88_54) );
AOI211_X1 g_91_54 (.ZN (n_91_54), .A (n_90_55), .B (n_84_58), .C1 (n_80_58), .C2 (n_86_55) );
AOI211_X1 g_90_52 (.ZN (n_90_52), .A (n_92_56), .B (n_86_57), .C1 (n_82_59), .C2 (n_84_56) );
AOI211_X1 g_89_54 (.ZN (n_89_54), .A (n_91_54), .B (n_88_56), .C1 (n_84_58), .C2 (n_82_57) );
AOI211_X1 g_87_55 (.ZN (n_87_55), .A (n_90_52), .B (n_90_55), .C1 (n_86_57), .C2 (n_80_58) );
AOI211_X1 g_88_53 (.ZN (n_88_53), .A (n_89_54), .B (n_92_56), .C1 (n_88_56), .C2 (n_82_59) );
AOI211_X1 g_86_54 (.ZN (n_86_54), .A (n_87_55), .B (n_91_54), .C1 (n_90_55), .C2 (n_84_58) );
AOI211_X1 g_85_56 (.ZN (n_85_56), .A (n_88_53), .B (n_90_52), .C1 (n_92_56), .C2 (n_86_57) );
AOI211_X1 g_83_57 (.ZN (n_83_57), .A (n_86_54), .B (n_89_54), .C1 (n_91_54), .C2 (n_88_56) );
AOI211_X1 g_84_55 (.ZN (n_84_55), .A (n_85_56), .B (n_87_55), .C1 (n_90_52), .C2 (n_90_55) );
AOI211_X1 g_82_56 (.ZN (n_82_56), .A (n_83_57), .B (n_88_53), .C1 (n_89_54), .C2 (n_92_56) );
AOI211_X1 g_80_57 (.ZN (n_80_57), .A (n_84_55), .B (n_86_54), .C1 (n_87_55), .C2 (n_91_54) );
AOI211_X1 g_78_58 (.ZN (n_78_58), .A (n_82_56), .B (n_85_56), .C1 (n_88_53), .C2 (n_90_52) );
AOI211_X1 g_76_59 (.ZN (n_76_59), .A (n_80_57), .B (n_83_57), .C1 (n_86_54), .C2 (n_89_54) );
AOI211_X1 g_74_60 (.ZN (n_74_60), .A (n_78_58), .B (n_84_55), .C1 (n_85_56), .C2 (n_87_55) );
AOI211_X1 g_72_61 (.ZN (n_72_61), .A (n_76_59), .B (n_82_56), .C1 (n_83_57), .C2 (n_88_53) );
AOI211_X1 g_70_62 (.ZN (n_70_62), .A (n_74_60), .B (n_80_57), .C1 (n_84_55), .C2 (n_86_54) );
AOI211_X1 g_69_60 (.ZN (n_69_60), .A (n_72_61), .B (n_78_58), .C1 (n_82_56), .C2 (n_85_56) );
AOI211_X1 g_67_61 (.ZN (n_67_61), .A (n_70_62), .B (n_76_59), .C1 (n_80_57), .C2 (n_83_57) );
AOI211_X1 g_65_62 (.ZN (n_65_62), .A (n_69_60), .B (n_74_60), .C1 (n_78_58), .C2 (n_84_55) );
AOI211_X1 g_63_63 (.ZN (n_63_63), .A (n_67_61), .B (n_72_61), .C1 (n_76_59), .C2 (n_82_56) );
AOI211_X1 g_61_64 (.ZN (n_61_64), .A (n_65_62), .B (n_70_62), .C1 (n_74_60), .C2 (n_80_57) );
AOI211_X1 g_59_65 (.ZN (n_59_65), .A (n_63_63), .B (n_69_60), .C1 (n_72_61), .C2 (n_78_58) );
AOI211_X1 g_57_66 (.ZN (n_57_66), .A (n_61_64), .B (n_67_61), .C1 (n_70_62), .C2 (n_76_59) );
AOI211_X1 g_55_67 (.ZN (n_55_67), .A (n_59_65), .B (n_65_62), .C1 (n_69_60), .C2 (n_74_60) );
AOI211_X1 g_53_68 (.ZN (n_53_68), .A (n_57_66), .B (n_63_63), .C1 (n_67_61), .C2 (n_72_61) );
AOI211_X1 g_51_67 (.ZN (n_51_67), .A (n_55_67), .B (n_61_64), .C1 (n_65_62), .C2 (n_70_62) );
AOI211_X1 g_49_68 (.ZN (n_49_68), .A (n_53_68), .B (n_59_65), .C1 (n_63_63), .C2 (n_69_60) );
AOI211_X1 g_47_69 (.ZN (n_47_69), .A (n_51_67), .B (n_57_66), .C1 (n_61_64), .C2 (n_67_61) );
AOI211_X1 g_46_71 (.ZN (n_46_71), .A (n_49_68), .B (n_55_67), .C1 (n_59_65), .C2 (n_65_62) );
AOI211_X1 g_48_70 (.ZN (n_48_70), .A (n_47_69), .B (n_53_68), .C1 (n_57_66), .C2 (n_63_63) );
AOI211_X1 g_50_69 (.ZN (n_50_69), .A (n_46_71), .B (n_51_67), .C1 (n_55_67), .C2 (n_61_64) );
AOI211_X1 g_52_68 (.ZN (n_52_68), .A (n_48_70), .B (n_49_68), .C1 (n_53_68), .C2 (n_59_65) );
AOI211_X1 g_54_67 (.ZN (n_54_67), .A (n_50_69), .B (n_47_69), .C1 (n_51_67), .C2 (n_57_66) );
AOI211_X1 g_56_66 (.ZN (n_56_66), .A (n_52_68), .B (n_46_71), .C1 (n_49_68), .C2 (n_55_67) );
AOI211_X1 g_58_65 (.ZN (n_58_65), .A (n_54_67), .B (n_48_70), .C1 (n_47_69), .C2 (n_53_68) );
AOI211_X1 g_60_64 (.ZN (n_60_64), .A (n_56_66), .B (n_50_69), .C1 (n_46_71), .C2 (n_51_67) );
AOI211_X1 g_62_63 (.ZN (n_62_63), .A (n_58_65), .B (n_52_68), .C1 (n_48_70), .C2 (n_49_68) );
AOI211_X1 g_64_62 (.ZN (n_64_62), .A (n_60_64), .B (n_54_67), .C1 (n_50_69), .C2 (n_47_69) );
AOI211_X1 g_66_61 (.ZN (n_66_61), .A (n_62_63), .B (n_56_66), .C1 (n_52_68), .C2 (n_46_71) );
AOI211_X1 g_68_62 (.ZN (n_68_62), .A (n_64_62), .B (n_58_65), .C1 (n_54_67), .C2 (n_48_70) );
AOI211_X1 g_66_63 (.ZN (n_66_63), .A (n_66_61), .B (n_60_64), .C1 (n_56_66), .C2 (n_50_69) );
AOI211_X1 g_64_64 (.ZN (n_64_64), .A (n_68_62), .B (n_62_63), .C1 (n_58_65), .C2 (n_52_68) );
AOI211_X1 g_62_65 (.ZN (n_62_65), .A (n_66_63), .B (n_64_62), .C1 (n_60_64), .C2 (n_54_67) );
AOI211_X1 g_60_66 (.ZN (n_60_66), .A (n_64_64), .B (n_66_61), .C1 (n_62_63), .C2 (n_56_66) );
AOI211_X1 g_58_67 (.ZN (n_58_67), .A (n_62_65), .B (n_68_62), .C1 (n_64_62), .C2 (n_58_65) );
AOI211_X1 g_56_68 (.ZN (n_56_68), .A (n_60_66), .B (n_66_63), .C1 (n_66_61), .C2 (n_60_64) );
AOI211_X1 g_54_69 (.ZN (n_54_69), .A (n_58_67), .B (n_64_64), .C1 (n_68_62), .C2 (n_62_63) );
AOI211_X1 g_52_70 (.ZN (n_52_70), .A (n_56_68), .B (n_62_65), .C1 (n_66_63), .C2 (n_64_62) );
AOI211_X1 g_50_71 (.ZN (n_50_71), .A (n_54_69), .B (n_60_66), .C1 (n_64_64), .C2 (n_66_61) );
AOI211_X1 g_51_69 (.ZN (n_51_69), .A (n_52_70), .B (n_58_67), .C1 (n_62_65), .C2 (n_68_62) );
AOI211_X1 g_53_70 (.ZN (n_53_70), .A (n_50_71), .B (n_56_68), .C1 (n_60_66), .C2 (n_66_63) );
AOI211_X1 g_55_69 (.ZN (n_55_69), .A (n_51_69), .B (n_54_69), .C1 (n_58_67), .C2 (n_64_64) );
AOI211_X1 g_57_68 (.ZN (n_57_68), .A (n_53_70), .B (n_52_70), .C1 (n_56_68), .C2 (n_62_65) );
AOI211_X1 g_59_67 (.ZN (n_59_67), .A (n_55_69), .B (n_50_71), .C1 (n_54_69), .C2 (n_60_66) );
AOI211_X1 g_60_65 (.ZN (n_60_65), .A (n_57_68), .B (n_51_69), .C1 (n_52_70), .C2 (n_58_67) );
AOI211_X1 g_62_64 (.ZN (n_62_64), .A (n_59_67), .B (n_53_70), .C1 (n_50_71), .C2 (n_56_68) );
AOI211_X1 g_64_63 (.ZN (n_64_63), .A (n_60_65), .B (n_55_69), .C1 (n_51_69), .C2 (n_54_69) );
AOI211_X1 g_63_65 (.ZN (n_63_65), .A (n_62_64), .B (n_57_68), .C1 (n_53_70), .C2 (n_52_70) );
AOI211_X1 g_61_66 (.ZN (n_61_66), .A (n_64_63), .B (n_59_67), .C1 (n_55_69), .C2 (n_50_71) );
AOI211_X1 g_60_68 (.ZN (n_60_68), .A (n_63_65), .B (n_60_65), .C1 (n_57_68), .C2 (n_51_69) );
AOI211_X1 g_59_66 (.ZN (n_59_66), .A (n_61_66), .B (n_62_64), .C1 (n_59_67), .C2 (n_53_70) );
AOI211_X1 g_61_65 (.ZN (n_61_65), .A (n_60_68), .B (n_64_63), .C1 (n_60_65), .C2 (n_55_69) );
AOI211_X1 g_63_64 (.ZN (n_63_64), .A (n_59_66), .B (n_63_65), .C1 (n_62_64), .C2 (n_57_68) );
AOI211_X1 g_65_63 (.ZN (n_65_63), .A (n_61_65), .B (n_61_66), .C1 (n_64_63), .C2 (n_59_67) );
AOI211_X1 g_67_62 (.ZN (n_67_62), .A (n_63_64), .B (n_60_68), .C1 (n_63_65), .C2 (n_60_65) );
AOI211_X1 g_66_64 (.ZN (n_66_64), .A (n_65_63), .B (n_59_66), .C1 (n_61_66), .C2 (n_62_64) );
AOI211_X1 g_68_63 (.ZN (n_68_63), .A (n_67_62), .B (n_61_65), .C1 (n_60_68), .C2 (n_64_63) );
AOI211_X1 g_67_65 (.ZN (n_67_65), .A (n_66_64), .B (n_63_64), .C1 (n_59_66), .C2 (n_63_65) );
AOI211_X1 g_65_64 (.ZN (n_65_64), .A (n_68_63), .B (n_65_63), .C1 (n_61_65), .C2 (n_61_66) );
AOI211_X1 g_67_63 (.ZN (n_67_63), .A (n_67_65), .B (n_67_62), .C1 (n_63_64), .C2 (n_60_68) );
AOI211_X1 g_69_62 (.ZN (n_69_62), .A (n_65_64), .B (n_66_64), .C1 (n_65_63), .C2 (n_59_66) );
AOI211_X1 g_71_61 (.ZN (n_71_61), .A (n_67_63), .B (n_68_63), .C1 (n_67_62), .C2 (n_61_65) );
AOI211_X1 g_70_63 (.ZN (n_70_63), .A (n_69_62), .B (n_67_65), .C1 (n_66_64), .C2 (n_63_64) );
AOI211_X1 g_68_64 (.ZN (n_68_64), .A (n_71_61), .B (n_65_64), .C1 (n_68_63), .C2 (n_65_63) );
AOI211_X1 g_66_65 (.ZN (n_66_65), .A (n_70_63), .B (n_67_63), .C1 (n_67_65), .C2 (n_67_62) );
AOI211_X1 g_64_66 (.ZN (n_64_66), .A (n_68_64), .B (n_69_62), .C1 (n_65_64), .C2 (n_66_64) );
AOI211_X1 g_62_67 (.ZN (n_62_67), .A (n_66_65), .B (n_71_61), .C1 (n_67_63), .C2 (n_68_63) );
AOI211_X1 g_61_69 (.ZN (n_61_69), .A (n_64_66), .B (n_70_63), .C1 (n_69_62), .C2 (n_67_65) );
AOI211_X1 g_60_67 (.ZN (n_60_67), .A (n_62_67), .B (n_68_64), .C1 (n_71_61), .C2 (n_65_64) );
AOI211_X1 g_62_66 (.ZN (n_62_66), .A (n_61_69), .B (n_66_65), .C1 (n_70_63), .C2 (n_67_63) );
AOI211_X1 g_64_65 (.ZN (n_64_65), .A (n_60_67), .B (n_64_66), .C1 (n_68_64), .C2 (n_69_62) );
AOI211_X1 g_63_67 (.ZN (n_63_67), .A (n_62_66), .B (n_62_67), .C1 (n_66_65), .C2 (n_71_61) );
AOI211_X1 g_65_66 (.ZN (n_65_66), .A (n_64_65), .B (n_61_69), .C1 (n_64_66), .C2 (n_70_63) );
AOI211_X1 g_64_68 (.ZN (n_64_68), .A (n_63_67), .B (n_60_67), .C1 (n_62_67), .C2 (n_68_64) );
AOI211_X1 g_63_66 (.ZN (n_63_66), .A (n_65_66), .B (n_62_66), .C1 (n_61_69), .C2 (n_66_65) );
AOI211_X1 g_65_65 (.ZN (n_65_65), .A (n_64_68), .B (n_64_65), .C1 (n_60_67), .C2 (n_64_66) );
AOI211_X1 g_67_64 (.ZN (n_67_64), .A (n_63_66), .B (n_63_67), .C1 (n_62_66), .C2 (n_62_67) );
AOI211_X1 g_69_63 (.ZN (n_69_63), .A (n_65_65), .B (n_65_66), .C1 (n_64_65), .C2 (n_61_69) );
AOI211_X1 g_71_62 (.ZN (n_71_62), .A (n_67_64), .B (n_64_68), .C1 (n_63_67), .C2 (n_60_67) );
AOI211_X1 g_73_61 (.ZN (n_73_61), .A (n_69_63), .B (n_63_66), .C1 (n_65_66), .C2 (n_62_66) );
AOI211_X1 g_75_60 (.ZN (n_75_60), .A (n_71_62), .B (n_65_65), .C1 (n_64_68), .C2 (n_64_65) );
AOI211_X1 g_77_59 (.ZN (n_77_59), .A (n_73_61), .B (n_67_64), .C1 (n_63_66), .C2 (n_63_67) );
AOI211_X1 g_79_58 (.ZN (n_79_58), .A (n_75_60), .B (n_69_63), .C1 (n_65_65), .C2 (n_65_66) );
AOI211_X1 g_78_60 (.ZN (n_78_60), .A (n_77_59), .B (n_71_62), .C1 (n_67_64), .C2 (n_64_68) );
AOI211_X1 g_80_59 (.ZN (n_80_59), .A (n_79_58), .B (n_73_61), .C1 (n_69_63), .C2 (n_63_66) );
AOI211_X1 g_82_58 (.ZN (n_82_58), .A (n_78_60), .B (n_75_60), .C1 (n_71_62), .C2 (n_65_65) );
AOI211_X1 g_84_57 (.ZN (n_84_57), .A (n_80_59), .B (n_77_59), .C1 (n_73_61), .C2 (n_67_64) );
AOI211_X1 g_86_56 (.ZN (n_86_56), .A (n_82_58), .B (n_79_58), .C1 (n_75_60), .C2 (n_69_63) );
AOI211_X1 g_88_55 (.ZN (n_88_55), .A (n_84_57), .B (n_78_60), .C1 (n_77_59), .C2 (n_71_62) );
AOI211_X1 g_90_54 (.ZN (n_90_54), .A (n_86_56), .B (n_80_59), .C1 (n_79_58), .C2 (n_73_61) );
AOI211_X1 g_92_53 (.ZN (n_92_53), .A (n_88_55), .B (n_82_58), .C1 (n_78_60), .C2 (n_75_60) );
AOI211_X1 g_91_55 (.ZN (n_91_55), .A (n_90_54), .B (n_84_57), .C1 (n_80_59), .C2 (n_77_59) );
AOI211_X1 g_89_56 (.ZN (n_89_56), .A (n_92_53), .B (n_86_56), .C1 (n_82_58), .C2 (n_79_58) );
AOI211_X1 g_87_57 (.ZN (n_87_57), .A (n_91_55), .B (n_88_55), .C1 (n_84_57), .C2 (n_78_60) );
AOI211_X1 g_85_58 (.ZN (n_85_58), .A (n_89_56), .B (n_90_54), .C1 (n_86_56), .C2 (n_80_59) );
AOI211_X1 g_83_59 (.ZN (n_83_59), .A (n_87_57), .B (n_92_53), .C1 (n_88_55), .C2 (n_82_58) );
AOI211_X1 g_81_58 (.ZN (n_81_58), .A (n_85_58), .B (n_91_55), .C1 (n_90_54), .C2 (n_84_57) );
AOI211_X1 g_79_59 (.ZN (n_79_59), .A (n_83_59), .B (n_89_56), .C1 (n_92_53), .C2 (n_86_56) );
AOI211_X1 g_77_60 (.ZN (n_77_60), .A (n_81_58), .B (n_87_57), .C1 (n_91_55), .C2 (n_88_55) );
AOI211_X1 g_75_61 (.ZN (n_75_61), .A (n_79_59), .B (n_85_58), .C1 (n_89_56), .C2 (n_90_54) );
AOI211_X1 g_73_62 (.ZN (n_73_62), .A (n_77_60), .B (n_83_59), .C1 (n_87_57), .C2 (n_92_53) );
AOI211_X1 g_71_63 (.ZN (n_71_63), .A (n_75_61), .B (n_81_58), .C1 (n_85_58), .C2 (n_91_55) );
AOI211_X1 g_69_64 (.ZN (n_69_64), .A (n_73_62), .B (n_79_59), .C1 (n_83_59), .C2 (n_89_56) );
AOI211_X1 g_68_66 (.ZN (n_68_66), .A (n_71_63), .B (n_77_60), .C1 (n_81_58), .C2 (n_87_57) );
AOI211_X1 g_66_67 (.ZN (n_66_67), .A (n_69_64), .B (n_75_61), .C1 (n_79_59), .C2 (n_85_58) );
AOI211_X1 g_65_69 (.ZN (n_65_69), .A (n_68_66), .B (n_73_62), .C1 (n_77_60), .C2 (n_83_59) );
AOI211_X1 g_64_67 (.ZN (n_64_67), .A (n_66_67), .B (n_71_63), .C1 (n_75_61), .C2 (n_81_58) );
AOI211_X1 g_66_66 (.ZN (n_66_66), .A (n_65_69), .B (n_69_64), .C1 (n_73_62), .C2 (n_79_59) );
AOI211_X1 g_68_65 (.ZN (n_68_65), .A (n_64_67), .B (n_68_66), .C1 (n_71_63), .C2 (n_77_60) );
AOI211_X1 g_70_64 (.ZN (n_70_64), .A (n_66_66), .B (n_66_67), .C1 (n_69_64), .C2 (n_75_61) );
AOI211_X1 g_72_63 (.ZN (n_72_63), .A (n_68_65), .B (n_65_69), .C1 (n_68_66), .C2 (n_73_62) );
AOI211_X1 g_74_62 (.ZN (n_74_62), .A (n_70_64), .B (n_64_67), .C1 (n_66_67), .C2 (n_71_63) );
AOI211_X1 g_76_61 (.ZN (n_76_61), .A (n_72_63), .B (n_66_66), .C1 (n_65_69), .C2 (n_69_64) );
AOI211_X1 g_75_63 (.ZN (n_75_63), .A (n_74_62), .B (n_68_65), .C1 (n_64_67), .C2 (n_68_66) );
AOI211_X1 g_77_62 (.ZN (n_77_62), .A (n_76_61), .B (n_70_64), .C1 (n_66_66), .C2 (n_66_67) );
AOI211_X1 g_79_61 (.ZN (n_79_61), .A (n_75_63), .B (n_72_63), .C1 (n_68_65), .C2 (n_65_69) );
AOI211_X1 g_81_60 (.ZN (n_81_60), .A (n_77_62), .B (n_74_62), .C1 (n_70_64), .C2 (n_64_67) );
AOI211_X1 g_83_61 (.ZN (n_83_61), .A (n_79_61), .B (n_76_61), .C1 (n_72_63), .C2 (n_66_66) );
AOI211_X1 g_85_60 (.ZN (n_85_60), .A (n_81_60), .B (n_75_63), .C1 (n_74_62), .C2 (n_68_65) );
AOI211_X1 g_87_59 (.ZN (n_87_59), .A (n_83_61), .B (n_77_62), .C1 (n_76_61), .C2 (n_70_64) );
AOI211_X1 g_89_58 (.ZN (n_89_58), .A (n_85_60), .B (n_79_61), .C1 (n_75_63), .C2 (n_72_63) );
AOI211_X1 g_90_56 (.ZN (n_90_56), .A (n_87_59), .B (n_81_60), .C1 (n_77_62), .C2 (n_74_62) );
AOI211_X1 g_92_55 (.ZN (n_92_55), .A (n_89_58), .B (n_83_61), .C1 (n_79_61), .C2 (n_76_61) );
AOI211_X1 g_94_54 (.ZN (n_94_54), .A (n_90_56), .B (n_85_60), .C1 (n_81_60), .C2 (n_75_63) );
AOI211_X1 g_96_55 (.ZN (n_96_55), .A (n_92_55), .B (n_87_59), .C1 (n_83_61), .C2 (n_77_62) );
AOI211_X1 g_94_56 (.ZN (n_94_56), .A (n_94_54), .B (n_89_58), .C1 (n_85_60), .C2 (n_79_61) );
AOI211_X1 g_92_57 (.ZN (n_92_57), .A (n_96_55), .B (n_90_56), .C1 (n_87_59), .C2 (n_81_60) );
AOI211_X1 g_93_55 (.ZN (n_93_55), .A (n_94_56), .B (n_92_55), .C1 (n_89_58), .C2 (n_83_61) );
AOI211_X1 g_94_57 (.ZN (n_94_57), .A (n_92_57), .B (n_94_54), .C1 (n_90_56), .C2 (n_85_60) );
AOI211_X1 g_95_59 (.ZN (n_95_59), .A (n_93_55), .B (n_96_55), .C1 (n_92_55), .C2 (n_87_59) );
AOI211_X1 g_96_61 (.ZN (n_96_61), .A (n_94_57), .B (n_94_56), .C1 (n_94_54), .C2 (n_89_58) );
AOI211_X1 g_97_63 (.ZN (n_97_63), .A (n_95_59), .B (n_92_57), .C1 (n_96_55), .C2 (n_90_56) );
AOI211_X1 g_98_65 (.ZN (n_98_65), .A (n_96_61), .B (n_93_55), .C1 (n_94_56), .C2 (n_92_55) );
AOI211_X1 g_99_67 (.ZN (n_99_67), .A (n_97_63), .B (n_94_57), .C1 (n_92_57), .C2 (n_94_54) );
AOI211_X1 g_100_69 (.ZN (n_100_69), .A (n_98_65), .B (n_95_59), .C1 (n_93_55), .C2 (n_96_55) );
AOI211_X1 g_98_70 (.ZN (n_98_70), .A (n_99_67), .B (n_96_61), .C1 (n_94_57), .C2 (n_94_56) );
AOI211_X1 g_100_71 (.ZN (n_100_71), .A (n_100_69), .B (n_97_63), .C1 (n_95_59), .C2 (n_92_57) );
AOI211_X1 g_99_69 (.ZN (n_99_69), .A (n_98_70), .B (n_98_65), .C1 (n_96_61), .C2 (n_93_55) );
AOI211_X1 g_97_68 (.ZN (n_97_68), .A (n_100_71), .B (n_99_67), .C1 (n_97_63), .C2 (n_94_57) );
AOI211_X1 g_96_66 (.ZN (n_96_66), .A (n_99_69), .B (n_100_69), .C1 (n_98_65), .C2 (n_95_59) );
AOI211_X1 g_98_67 (.ZN (n_98_67), .A (n_97_68), .B (n_98_70), .C1 (n_99_67), .C2 (n_96_61) );
AOI211_X1 g_100_68 (.ZN (n_100_68), .A (n_96_66), .B (n_100_71), .C1 (n_100_69), .C2 (n_97_63) );
AOI211_X1 g_99_66 (.ZN (n_99_66), .A (n_98_67), .B (n_99_69), .C1 (n_98_70), .C2 (n_98_65) );
AOI211_X1 g_98_64 (.ZN (n_98_64), .A (n_100_68), .B (n_97_68), .C1 (n_100_71), .C2 (n_99_67) );
AOI211_X1 g_97_62 (.ZN (n_97_62), .A (n_99_66), .B (n_96_66), .C1 (n_99_69), .C2 (n_100_69) );
AOI211_X1 g_96_60 (.ZN (n_96_60), .A (n_98_64), .B (n_98_67), .C1 (n_97_68), .C2 (n_98_70) );
AOI211_X1 g_95_58 (.ZN (n_95_58), .A (n_97_62), .B (n_100_68), .C1 (n_96_66), .C2 (n_100_71) );
AOI211_X1 g_97_57 (.ZN (n_97_57), .A (n_96_60), .B (n_99_66), .C1 (n_98_67), .C2 (n_99_69) );
AOI211_X1 g_95_56 (.ZN (n_95_56), .A (n_95_58), .B (n_98_64), .C1 (n_100_68), .C2 (n_97_68) );
AOI211_X1 g_93_57 (.ZN (n_93_57), .A (n_97_57), .B (n_97_62), .C1 (n_99_66), .C2 (n_96_66) );
AOI211_X1 g_91_56 (.ZN (n_91_56), .A (n_95_56), .B (n_96_60), .C1 (n_98_64), .C2 (n_98_67) );
AOI211_X1 g_89_55 (.ZN (n_89_55), .A (n_93_57), .B (n_95_58), .C1 (n_97_62), .C2 (n_100_68) );
AOI211_X1 g_88_57 (.ZN (n_88_57), .A (n_91_56), .B (n_97_57), .C1 (n_96_60), .C2 (n_99_66) );
AOI211_X1 g_86_58 (.ZN (n_86_58), .A (n_89_55), .B (n_95_56), .C1 (n_95_58), .C2 (n_98_64) );
AOI211_X1 g_87_56 (.ZN (n_87_56), .A (n_88_57), .B (n_93_57), .C1 (n_97_57), .C2 (n_97_62) );
AOI211_X1 g_85_57 (.ZN (n_85_57), .A (n_86_58), .B (n_91_56), .C1 (n_95_56), .C2 (n_96_60) );
AOI211_X1 g_84_59 (.ZN (n_84_59), .A (n_87_56), .B (n_89_55), .C1 (n_93_57), .C2 (n_95_58) );
AOI211_X1 g_82_60 (.ZN (n_82_60), .A (n_85_57), .B (n_88_57), .C1 (n_91_56), .C2 (n_97_57) );
AOI211_X1 g_83_58 (.ZN (n_83_58), .A (n_84_59), .B (n_86_58), .C1 (n_89_55), .C2 (n_95_56) );
AOI211_X1 g_81_59 (.ZN (n_81_59), .A (n_82_60), .B (n_87_56), .C1 (n_88_57), .C2 (n_93_57) );
AOI211_X1 g_79_60 (.ZN (n_79_60), .A (n_83_58), .B (n_85_57), .C1 (n_86_58), .C2 (n_91_56) );
AOI211_X1 g_77_61 (.ZN (n_77_61), .A (n_81_59), .B (n_84_59), .C1 (n_87_56), .C2 (n_89_55) );
AOI211_X1 g_75_62 (.ZN (n_75_62), .A (n_79_60), .B (n_82_60), .C1 (n_85_57), .C2 (n_88_57) );
AOI211_X1 g_73_63 (.ZN (n_73_63), .A (n_77_61), .B (n_83_58), .C1 (n_84_59), .C2 (n_86_58) );
AOI211_X1 g_71_64 (.ZN (n_71_64), .A (n_75_62), .B (n_81_59), .C1 (n_82_60), .C2 (n_87_56) );
AOI211_X1 g_69_65 (.ZN (n_69_65), .A (n_73_63), .B (n_79_60), .C1 (n_83_58), .C2 (n_85_57) );
AOI211_X1 g_67_66 (.ZN (n_67_66), .A (n_71_64), .B (n_77_61), .C1 (n_81_59), .C2 (n_84_59) );
AOI211_X1 g_65_67 (.ZN (n_65_67), .A (n_69_65), .B (n_75_62), .C1 (n_79_60), .C2 (n_82_60) );
AOI211_X1 g_63_68 (.ZN (n_63_68), .A (n_67_66), .B (n_73_63), .C1 (n_77_61), .C2 (n_83_58) );
AOI211_X1 g_61_67 (.ZN (n_61_67), .A (n_65_67), .B (n_71_64), .C1 (n_75_62), .C2 (n_81_59) );
AOI211_X1 g_59_68 (.ZN (n_59_68), .A (n_63_68), .B (n_69_65), .C1 (n_73_63), .C2 (n_79_60) );
AOI211_X1 g_57_67 (.ZN (n_57_67), .A (n_61_67), .B (n_67_66), .C1 (n_71_64), .C2 (n_77_61) );
AOI211_X1 g_55_68 (.ZN (n_55_68), .A (n_59_68), .B (n_65_67), .C1 (n_69_65), .C2 (n_75_62) );
AOI211_X1 g_53_69 (.ZN (n_53_69), .A (n_57_67), .B (n_63_68), .C1 (n_67_66), .C2 (n_73_63) );
AOI211_X1 g_51_70 (.ZN (n_51_70), .A (n_55_68), .B (n_61_67), .C1 (n_65_67), .C2 (n_71_64) );
AOI211_X1 g_49_71 (.ZN (n_49_71), .A (n_53_69), .B (n_59_68), .C1 (n_63_68), .C2 (n_69_65) );
AOI211_X1 g_47_72 (.ZN (n_47_72), .A (n_51_70), .B (n_57_67), .C1 (n_61_67), .C2 (n_67_66) );
AOI211_X1 g_45_73 (.ZN (n_45_73), .A (n_49_71), .B (n_55_68), .C1 (n_59_68), .C2 (n_65_67) );
AOI211_X1 g_43_74 (.ZN (n_43_74), .A (n_47_72), .B (n_53_69), .C1 (n_57_67), .C2 (n_63_68) );
AOI211_X1 g_44_72 (.ZN (n_44_72), .A (n_45_73), .B (n_51_70), .C1 (n_55_68), .C2 (n_61_67) );
AOI211_X1 g_42_73 (.ZN (n_42_73), .A (n_43_74), .B (n_49_71), .C1 (n_53_69), .C2 (n_59_68) );
AOI211_X1 g_40_74 (.ZN (n_40_74), .A (n_44_72), .B (n_47_72), .C1 (n_51_70), .C2 (n_57_67) );
AOI211_X1 g_38_75 (.ZN (n_38_75), .A (n_42_73), .B (n_45_73), .C1 (n_49_71), .C2 (n_55_68) );
AOI211_X1 g_36_76 (.ZN (n_36_76), .A (n_40_74), .B (n_43_74), .C1 (n_47_72), .C2 (n_53_69) );
AOI211_X1 g_34_77 (.ZN (n_34_77), .A (n_38_75), .B (n_44_72), .C1 (n_45_73), .C2 (n_51_70) );
AOI211_X1 g_32_78 (.ZN (n_32_78), .A (n_36_76), .B (n_42_73), .C1 (n_43_74), .C2 (n_49_71) );
AOI211_X1 g_30_79 (.ZN (n_30_79), .A (n_34_77), .B (n_40_74), .C1 (n_44_72), .C2 (n_47_72) );
AOI211_X1 g_28_80 (.ZN (n_28_80), .A (n_32_78), .B (n_38_75), .C1 (n_42_73), .C2 (n_45_73) );
AOI211_X1 g_26_81 (.ZN (n_26_81), .A (n_30_79), .B (n_36_76), .C1 (n_40_74), .C2 (n_43_74) );
AOI211_X1 g_24_80 (.ZN (n_24_80), .A (n_28_80), .B (n_34_77), .C1 (n_38_75), .C2 (n_44_72) );
AOI211_X1 g_22_81 (.ZN (n_22_81), .A (n_26_81), .B (n_32_78), .C1 (n_36_76), .C2 (n_42_73) );
AOI211_X1 g_20_82 (.ZN (n_20_82), .A (n_24_80), .B (n_30_79), .C1 (n_34_77), .C2 (n_40_74) );
AOI211_X1 g_18_83 (.ZN (n_18_83), .A (n_22_81), .B (n_28_80), .C1 (n_32_78), .C2 (n_38_75) );
AOI211_X1 g_16_84 (.ZN (n_16_84), .A (n_20_82), .B (n_26_81), .C1 (n_30_79), .C2 (n_36_76) );
AOI211_X1 g_14_85 (.ZN (n_14_85), .A (n_18_83), .B (n_24_80), .C1 (n_28_80), .C2 (n_34_77) );
AOI211_X1 g_12_86 (.ZN (n_12_86), .A (n_16_84), .B (n_22_81), .C1 (n_26_81), .C2 (n_32_78) );
AOI211_X1 g_10_87 (.ZN (n_10_87), .A (n_14_85), .B (n_20_82), .C1 (n_24_80), .C2 (n_30_79) );
AOI211_X1 g_9_89 (.ZN (n_9_89), .A (n_12_86), .B (n_18_83), .C1 (n_22_81), .C2 (n_28_80) );
AOI211_X1 g_11_88 (.ZN (n_11_88), .A (n_10_87), .B (n_16_84), .C1 (n_20_82), .C2 (n_26_81) );
AOI211_X1 g_13_87 (.ZN (n_13_87), .A (n_9_89), .B (n_14_85), .C1 (n_18_83), .C2 (n_24_80) );
AOI211_X1 g_11_86 (.ZN (n_11_86), .A (n_11_88), .B (n_12_86), .C1 (n_16_84), .C2 (n_22_81) );
AOI211_X1 g_13_85 (.ZN (n_13_85), .A (n_13_87), .B (n_10_87), .C1 (n_14_85), .C2 (n_20_82) );
AOI211_X1 g_15_84 (.ZN (n_15_84), .A (n_11_86), .B (n_9_89), .C1 (n_12_86), .C2 (n_18_83) );
AOI211_X1 g_17_83 (.ZN (n_17_83), .A (n_13_85), .B (n_11_88), .C1 (n_10_87), .C2 (n_16_84) );
AOI211_X1 g_19_82 (.ZN (n_19_82), .A (n_15_84), .B (n_13_87), .C1 (n_9_89), .C2 (n_14_85) );
AOI211_X1 g_21_81 (.ZN (n_21_81), .A (n_17_83), .B (n_11_86), .C1 (n_11_88), .C2 (n_12_86) );
AOI211_X1 g_23_80 (.ZN (n_23_80), .A (n_19_82), .B (n_13_85), .C1 (n_13_87), .C2 (n_10_87) );
AOI211_X1 g_24_82 (.ZN (n_24_82), .A (n_21_81), .B (n_15_84), .C1 (n_11_86), .C2 (n_9_89) );
AOI211_X1 g_22_83 (.ZN (n_22_83), .A (n_23_80), .B (n_17_83), .C1 (n_13_85), .C2 (n_11_88) );
AOI211_X1 g_20_84 (.ZN (n_20_84), .A (n_24_82), .B (n_19_82), .C1 (n_15_84), .C2 (n_13_87) );
AOI211_X1 g_18_85 (.ZN (n_18_85), .A (n_22_83), .B (n_21_81), .C1 (n_17_83), .C2 (n_11_86) );
AOI211_X1 g_16_86 (.ZN (n_16_86), .A (n_20_84), .B (n_23_80), .C1 (n_19_82), .C2 (n_13_85) );
AOI211_X1 g_14_87 (.ZN (n_14_87), .A (n_18_85), .B (n_24_82), .C1 (n_21_81), .C2 (n_15_84) );
AOI211_X1 g_12_88 (.ZN (n_12_88), .A (n_16_86), .B (n_22_83), .C1 (n_23_80), .C2 (n_17_83) );
AOI211_X1 g_10_89 (.ZN (n_10_89), .A (n_14_87), .B (n_20_84), .C1 (n_24_82), .C2 (n_19_82) );
AOI211_X1 g_11_87 (.ZN (n_11_87), .A (n_12_88), .B (n_18_85), .C1 (n_22_83), .C2 (n_21_81) );
AOI211_X1 g_9_88 (.ZN (n_9_88), .A (n_10_89), .B (n_16_86), .C1 (n_20_84), .C2 (n_23_80) );
AOI211_X1 g_7_89 (.ZN (n_7_89), .A (n_11_87), .B (n_14_87), .C1 (n_18_85), .C2 (n_24_82) );
AOI211_X1 g_6_91 (.ZN (n_6_91), .A (n_9_88), .B (n_12_88), .C1 (n_16_86), .C2 (n_22_83) );
AOI211_X1 g_8_90 (.ZN (n_8_90), .A (n_7_89), .B (n_10_89), .C1 (n_14_87), .C2 (n_20_84) );
AOI211_X1 g_7_92 (.ZN (n_7_92), .A (n_6_91), .B (n_11_87), .C1 (n_12_88), .C2 (n_18_85) );
AOI211_X1 g_5_93 (.ZN (n_5_93), .A (n_8_90), .B (n_9_88), .C1 (n_10_89), .C2 (n_16_86) );
AOI211_X1 g_4_95 (.ZN (n_4_95), .A (n_7_92), .B (n_7_89), .C1 (n_11_87), .C2 (n_14_87) );
AOI211_X1 g_3_97 (.ZN (n_3_97), .A (n_5_93), .B (n_6_91), .C1 (n_9_88), .C2 (n_12_88) );
AOI211_X1 g_4_99 (.ZN (n_4_99), .A (n_4_95), .B (n_8_90), .C1 (n_7_89), .C2 (n_10_89) );
AOI211_X1 g_6_100 (.ZN (n_6_100), .A (n_3_97), .B (n_7_92), .C1 (n_6_91), .C2 (n_11_87) );
AOI211_X1 g_5_98 (.ZN (n_5_98), .A (n_4_99), .B (n_5_93), .C1 (n_8_90), .C2 (n_9_88) );
AOI211_X1 g_6_96 (.ZN (n_6_96), .A (n_6_100), .B (n_4_95), .C1 (n_7_92), .C2 (n_7_89) );
AOI211_X1 g_7_94 (.ZN (n_7_94), .A (n_5_98), .B (n_3_97), .C1 (n_5_93), .C2 (n_6_91) );
AOI211_X1 g_8_92 (.ZN (n_8_92), .A (n_6_96), .B (n_4_99), .C1 (n_4_95), .C2 (n_8_90) );
AOI211_X1 g_9_90 (.ZN (n_9_90), .A (n_7_94), .B (n_6_100), .C1 (n_3_97), .C2 (n_7_92) );
AOI211_X1 g_10_88 (.ZN (n_10_88), .A (n_8_92), .B (n_5_98), .C1 (n_4_99), .C2 (n_5_93) );
AOI211_X1 g_12_87 (.ZN (n_12_87), .A (n_9_90), .B (n_6_96), .C1 (n_6_100), .C2 (n_4_95) );
AOI211_X1 g_14_86 (.ZN (n_14_86), .A (n_10_88), .B (n_7_94), .C1 (n_5_98), .C2 (n_3_97) );
AOI211_X1 g_16_85 (.ZN (n_16_85), .A (n_12_87), .B (n_8_92), .C1 (n_6_96), .C2 (n_4_99) );
AOI211_X1 g_18_84 (.ZN (n_18_84), .A (n_14_86), .B (n_9_90), .C1 (n_7_94), .C2 (n_6_100) );
AOI211_X1 g_20_83 (.ZN (n_20_83), .A (n_16_85), .B (n_10_88), .C1 (n_8_92), .C2 (n_5_98) );
AOI211_X1 g_22_82 (.ZN (n_22_82), .A (n_18_84), .B (n_12_87), .C1 (n_9_90), .C2 (n_6_96) );
AOI211_X1 g_24_81 (.ZN (n_24_81), .A (n_20_83), .B (n_14_86), .C1 (n_10_88), .C2 (n_7_94) );
AOI211_X1 g_26_80 (.ZN (n_26_80), .A (n_22_82), .B (n_16_85), .C1 (n_12_87), .C2 (n_8_92) );
AOI211_X1 g_25_82 (.ZN (n_25_82), .A (n_24_81), .B (n_18_84), .C1 (n_14_86), .C2 (n_9_90) );
AOI211_X1 g_23_83 (.ZN (n_23_83), .A (n_26_80), .B (n_20_83), .C1 (n_16_85), .C2 (n_10_88) );
AOI211_X1 g_21_84 (.ZN (n_21_84), .A (n_25_82), .B (n_22_82), .C1 (n_18_84), .C2 (n_12_87) );
AOI211_X1 g_19_85 (.ZN (n_19_85), .A (n_23_83), .B (n_24_81), .C1 (n_20_83), .C2 (n_14_86) );
AOI211_X1 g_17_86 (.ZN (n_17_86), .A (n_21_84), .B (n_26_80), .C1 (n_22_82), .C2 (n_16_85) );
AOI211_X1 g_15_87 (.ZN (n_15_87), .A (n_19_85), .B (n_25_82), .C1 (n_24_81), .C2 (n_18_84) );
AOI211_X1 g_13_88 (.ZN (n_13_88), .A (n_17_86), .B (n_23_83), .C1 (n_26_80), .C2 (n_20_83) );
AOI211_X1 g_11_89 (.ZN (n_11_89), .A (n_15_87), .B (n_21_84), .C1 (n_25_82), .C2 (n_22_82) );
AOI211_X1 g_10_91 (.ZN (n_10_91), .A (n_13_88), .B (n_19_85), .C1 (n_23_83), .C2 (n_24_81) );
AOI211_X1 g_12_90 (.ZN (n_12_90), .A (n_11_89), .B (n_17_86), .C1 (n_21_84), .C2 (n_26_80) );
AOI211_X1 g_14_89 (.ZN (n_14_89), .A (n_10_91), .B (n_15_87), .C1 (n_19_85), .C2 (n_25_82) );
AOI211_X1 g_16_88 (.ZN (n_16_88), .A (n_12_90), .B (n_13_88), .C1 (n_17_86), .C2 (n_23_83) );
AOI211_X1 g_15_86 (.ZN (n_15_86), .A (n_14_89), .B (n_11_89), .C1 (n_15_87), .C2 (n_21_84) );
AOI211_X1 g_17_85 (.ZN (n_17_85), .A (n_16_88), .B (n_10_91), .C1 (n_13_88), .C2 (n_19_85) );
AOI211_X1 g_19_84 (.ZN (n_19_84), .A (n_15_86), .B (n_12_90), .C1 (n_11_89), .C2 (n_17_86) );
AOI211_X1 g_21_83 (.ZN (n_21_83), .A (n_17_85), .B (n_14_89), .C1 (n_10_91), .C2 (n_15_87) );
AOI211_X1 g_23_82 (.ZN (n_23_82), .A (n_19_84), .B (n_16_88), .C1 (n_12_90), .C2 (n_13_88) );
AOI211_X1 g_25_81 (.ZN (n_25_81), .A (n_21_83), .B (n_15_86), .C1 (n_14_89), .C2 (n_11_89) );
AOI211_X1 g_27_80 (.ZN (n_27_80), .A (n_23_82), .B (n_17_85), .C1 (n_16_88), .C2 (n_10_91) );
AOI211_X1 g_29_79 (.ZN (n_29_79), .A (n_25_81), .B (n_19_84), .C1 (n_15_86), .C2 (n_12_90) );
AOI211_X1 g_28_81 (.ZN (n_28_81), .A (n_27_80), .B (n_21_83), .C1 (n_17_85), .C2 (n_14_89) );
AOI211_X1 g_30_80 (.ZN (n_30_80), .A (n_29_79), .B (n_23_82), .C1 (n_19_84), .C2 (n_16_88) );
AOI211_X1 g_32_79 (.ZN (n_32_79), .A (n_28_81), .B (n_25_81), .C1 (n_21_83), .C2 (n_15_86) );
AOI211_X1 g_34_78 (.ZN (n_34_78), .A (n_30_80), .B (n_27_80), .C1 (n_23_82), .C2 (n_17_85) );
AOI211_X1 g_36_77 (.ZN (n_36_77), .A (n_32_79), .B (n_29_79), .C1 (n_25_81), .C2 (n_19_84) );
AOI211_X1 g_38_76 (.ZN (n_38_76), .A (n_34_78), .B (n_28_81), .C1 (n_27_80), .C2 (n_21_83) );
AOI211_X1 g_40_75 (.ZN (n_40_75), .A (n_36_77), .B (n_30_80), .C1 (n_29_79), .C2 (n_23_82) );
AOI211_X1 g_42_74 (.ZN (n_42_74), .A (n_38_76), .B (n_32_79), .C1 (n_28_81), .C2 (n_25_81) );
AOI211_X1 g_44_73 (.ZN (n_44_73), .A (n_40_75), .B (n_34_78), .C1 (n_30_80), .C2 (n_27_80) );
AOI211_X1 g_46_72 (.ZN (n_46_72), .A (n_42_74), .B (n_36_77), .C1 (n_32_79), .C2 (n_29_79) );
AOI211_X1 g_48_71 (.ZN (n_48_71), .A (n_44_73), .B (n_38_76), .C1 (n_34_78), .C2 (n_28_81) );
AOI211_X1 g_50_70 (.ZN (n_50_70), .A (n_46_72), .B (n_40_75), .C1 (n_36_77), .C2 (n_30_80) );
AOI211_X1 g_52_69 (.ZN (n_52_69), .A (n_48_71), .B (n_42_74), .C1 (n_38_76), .C2 (n_32_79) );
AOI211_X1 g_51_71 (.ZN (n_51_71), .A (n_50_70), .B (n_44_73), .C1 (n_40_75), .C2 (n_34_78) );
AOI211_X1 g_49_72 (.ZN (n_49_72), .A (n_52_69), .B (n_46_72), .C1 (n_42_74), .C2 (n_36_77) );
AOI211_X1 g_47_71 (.ZN (n_47_71), .A (n_51_71), .B (n_48_71), .C1 (n_44_73), .C2 (n_38_76) );
AOI211_X1 g_45_72 (.ZN (n_45_72), .A (n_49_72), .B (n_50_70), .C1 (n_46_72), .C2 (n_40_75) );
AOI211_X1 g_43_73 (.ZN (n_43_73), .A (n_47_71), .B (n_52_69), .C1 (n_48_71), .C2 (n_42_74) );
AOI211_X1 g_41_74 (.ZN (n_41_74), .A (n_45_72), .B (n_51_71), .C1 (n_50_70), .C2 (n_44_73) );
AOI211_X1 g_39_75 (.ZN (n_39_75), .A (n_43_73), .B (n_49_72), .C1 (n_52_69), .C2 (n_46_72) );
AOI211_X1 g_37_76 (.ZN (n_37_76), .A (n_41_74), .B (n_47_71), .C1 (n_51_71), .C2 (n_48_71) );
AOI211_X1 g_35_77 (.ZN (n_35_77), .A (n_39_75), .B (n_45_72), .C1 (n_49_72), .C2 (n_50_70) );
AOI211_X1 g_33_78 (.ZN (n_33_78), .A (n_37_76), .B (n_43_73), .C1 (n_47_71), .C2 (n_52_69) );
AOI211_X1 g_31_79 (.ZN (n_31_79), .A (n_35_77), .B (n_41_74), .C1 (n_45_72), .C2 (n_51_71) );
AOI211_X1 g_29_80 (.ZN (n_29_80), .A (n_33_78), .B (n_39_75), .C1 (n_43_73), .C2 (n_49_72) );
AOI211_X1 g_28_82 (.ZN (n_28_82), .A (n_31_79), .B (n_37_76), .C1 (n_41_74), .C2 (n_47_71) );
AOI211_X1 g_30_81 (.ZN (n_30_81), .A (n_29_80), .B (n_35_77), .C1 (n_39_75), .C2 (n_45_72) );
AOI211_X1 g_32_80 (.ZN (n_32_80), .A (n_28_82), .B (n_33_78), .C1 (n_37_76), .C2 (n_43_73) );
AOI211_X1 g_34_79 (.ZN (n_34_79), .A (n_30_81), .B (n_31_79), .C1 (n_35_77), .C2 (n_41_74) );
AOI211_X1 g_36_78 (.ZN (n_36_78), .A (n_32_80), .B (n_29_80), .C1 (n_33_78), .C2 (n_39_75) );
AOI211_X1 g_38_77 (.ZN (n_38_77), .A (n_34_79), .B (n_28_82), .C1 (n_31_79), .C2 (n_37_76) );
AOI211_X1 g_40_76 (.ZN (n_40_76), .A (n_36_78), .B (n_30_81), .C1 (n_29_80), .C2 (n_35_77) );
AOI211_X1 g_42_75 (.ZN (n_42_75), .A (n_38_77), .B (n_32_80), .C1 (n_28_82), .C2 (n_33_78) );
AOI211_X1 g_44_74 (.ZN (n_44_74), .A (n_40_76), .B (n_34_79), .C1 (n_30_81), .C2 (n_31_79) );
AOI211_X1 g_46_73 (.ZN (n_46_73), .A (n_42_75), .B (n_36_78), .C1 (n_32_80), .C2 (n_29_80) );
AOI211_X1 g_48_72 (.ZN (n_48_72), .A (n_44_74), .B (n_38_77), .C1 (n_34_79), .C2 (n_28_82) );
AOI211_X1 g_47_74 (.ZN (n_47_74), .A (n_46_73), .B (n_40_76), .C1 (n_36_78), .C2 (n_30_81) );
AOI211_X1 g_49_73 (.ZN (n_49_73), .A (n_48_72), .B (n_42_75), .C1 (n_38_77), .C2 (n_32_80) );
AOI211_X1 g_51_72 (.ZN (n_51_72), .A (n_47_74), .B (n_44_74), .C1 (n_40_76), .C2 (n_34_79) );
AOI211_X1 g_53_71 (.ZN (n_53_71), .A (n_49_73), .B (n_46_73), .C1 (n_42_75), .C2 (n_36_78) );
AOI211_X1 g_55_70 (.ZN (n_55_70), .A (n_51_72), .B (n_48_72), .C1 (n_44_74), .C2 (n_38_77) );
AOI211_X1 g_57_69 (.ZN (n_57_69), .A (n_53_71), .B (n_47_74), .C1 (n_46_73), .C2 (n_40_76) );
AOI211_X1 g_59_70 (.ZN (n_59_70), .A (n_55_70), .B (n_49_73), .C1 (n_48_72), .C2 (n_42_75) );
AOI211_X1 g_58_68 (.ZN (n_58_68), .A (n_57_69), .B (n_51_72), .C1 (n_47_74), .C2 (n_44_74) );
AOI211_X1 g_56_69 (.ZN (n_56_69), .A (n_59_70), .B (n_53_71), .C1 (n_49_73), .C2 (n_46_73) );
AOI211_X1 g_54_70 (.ZN (n_54_70), .A (n_58_68), .B (n_55_70), .C1 (n_51_72), .C2 (n_48_72) );
AOI211_X1 g_52_71 (.ZN (n_52_71), .A (n_56_69), .B (n_57_69), .C1 (n_53_71), .C2 (n_47_74) );
AOI211_X1 g_50_72 (.ZN (n_50_72), .A (n_54_70), .B (n_59_70), .C1 (n_55_70), .C2 (n_49_73) );
AOI211_X1 g_48_73 (.ZN (n_48_73), .A (n_52_71), .B (n_58_68), .C1 (n_57_69), .C2 (n_51_72) );
AOI211_X1 g_46_74 (.ZN (n_46_74), .A (n_50_72), .B (n_56_69), .C1 (n_59_70), .C2 (n_53_71) );
AOI211_X1 g_44_75 (.ZN (n_44_75), .A (n_48_73), .B (n_54_70), .C1 (n_58_68), .C2 (n_55_70) );
AOI211_X1 g_42_76 (.ZN (n_42_76), .A (n_46_74), .B (n_52_71), .C1 (n_56_69), .C2 (n_57_69) );
AOI211_X1 g_40_77 (.ZN (n_40_77), .A (n_44_75), .B (n_50_72), .C1 (n_54_70), .C2 (n_59_70) );
AOI211_X1 g_41_75 (.ZN (n_41_75), .A (n_42_76), .B (n_48_73), .C1 (n_52_71), .C2 (n_58_68) );
AOI211_X1 g_39_76 (.ZN (n_39_76), .A (n_40_77), .B (n_46_74), .C1 (n_50_72), .C2 (n_56_69) );
AOI211_X1 g_37_77 (.ZN (n_37_77), .A (n_41_75), .B (n_44_75), .C1 (n_48_73), .C2 (n_54_70) );
AOI211_X1 g_35_78 (.ZN (n_35_78), .A (n_39_76), .B (n_42_76), .C1 (n_46_74), .C2 (n_52_71) );
AOI211_X1 g_33_79 (.ZN (n_33_79), .A (n_37_77), .B (n_40_77), .C1 (n_44_75), .C2 (n_50_72) );
AOI211_X1 g_31_80 (.ZN (n_31_80), .A (n_35_78), .B (n_41_75), .C1 (n_42_76), .C2 (n_48_73) );
AOI211_X1 g_29_81 (.ZN (n_29_81), .A (n_33_79), .B (n_39_76), .C1 (n_40_77), .C2 (n_46_74) );
AOI211_X1 g_27_82 (.ZN (n_27_82), .A (n_31_80), .B (n_37_77), .C1 (n_41_75), .C2 (n_44_75) );
AOI211_X1 g_25_83 (.ZN (n_25_83), .A (n_29_81), .B (n_35_78), .C1 (n_39_76), .C2 (n_42_76) );
AOI211_X1 g_23_84 (.ZN (n_23_84), .A (n_27_82), .B (n_33_79), .C1 (n_37_77), .C2 (n_40_77) );
AOI211_X1 g_21_85 (.ZN (n_21_85), .A (n_25_83), .B (n_31_80), .C1 (n_35_78), .C2 (n_41_75) );
AOI211_X1 g_19_86 (.ZN (n_19_86), .A (n_23_84), .B (n_29_81), .C1 (n_33_79), .C2 (n_39_76) );
AOI211_X1 g_17_87 (.ZN (n_17_87), .A (n_21_85), .B (n_27_82), .C1 (n_31_80), .C2 (n_37_77) );
AOI211_X1 g_15_88 (.ZN (n_15_88), .A (n_19_86), .B (n_25_83), .C1 (n_29_81), .C2 (n_35_78) );
AOI211_X1 g_13_89 (.ZN (n_13_89), .A (n_17_87), .B (n_23_84), .C1 (n_27_82), .C2 (n_33_79) );
AOI211_X1 g_11_90 (.ZN (n_11_90), .A (n_15_88), .B (n_21_85), .C1 (n_25_83), .C2 (n_31_80) );
AOI211_X1 g_9_91 (.ZN (n_9_91), .A (n_13_89), .B (n_19_86), .C1 (n_23_84), .C2 (n_29_81) );
AOI211_X1 g_8_93 (.ZN (n_8_93), .A (n_11_90), .B (n_17_87), .C1 (n_21_85), .C2 (n_27_82) );
AOI211_X1 g_6_94 (.ZN (n_6_94), .A (n_9_91), .B (n_15_88), .C1 (n_19_86), .C2 (n_25_83) );
AOI211_X1 g_5_96 (.ZN (n_5_96), .A (n_8_93), .B (n_13_89), .C1 (n_17_87), .C2 (n_23_84) );
AOI211_X1 g_4_98 (.ZN (n_4_98), .A (n_6_94), .B (n_11_90), .C1 (n_15_88), .C2 (n_21_85) );
AOI211_X1 g_5_100 (.ZN (n_5_100), .A (n_5_96), .B (n_9_91), .C1 (n_13_89), .C2 (n_19_86) );
AOI211_X1 g_6_98 (.ZN (n_6_98), .A (n_4_98), .B (n_8_93), .C1 (n_11_90), .C2 (n_17_87) );
AOI211_X1 g_8_99 (.ZN (n_8_99), .A (n_5_100), .B (n_6_94), .C1 (n_9_91), .C2 (n_15_88) );
AOI211_X1 g_10_100 (.ZN (n_10_100), .A (n_6_98), .B (n_5_96), .C1 (n_8_93), .C2 (n_13_89) );
AOI211_X1 g_12_99 (.ZN (n_12_99), .A (n_8_99), .B (n_4_98), .C1 (n_6_94), .C2 (n_11_90) );
AOI211_X1 g_14_100 (.ZN (n_14_100), .A (n_10_100), .B (n_5_100), .C1 (n_5_96), .C2 (n_9_91) );
AOI211_X1 g_16_99 (.ZN (n_16_99), .A (n_12_99), .B (n_6_98), .C1 (n_4_98), .C2 (n_8_93) );
AOI211_X1 g_18_100 (.ZN (n_18_100), .A (n_14_100), .B (n_8_99), .C1 (n_5_100), .C2 (n_6_94) );
AOI211_X1 g_20_99 (.ZN (n_20_99), .A (n_16_99), .B (n_10_100), .C1 (n_6_98), .C2 (n_5_96) );
AOI211_X1 g_22_100 (.ZN (n_22_100), .A (n_18_100), .B (n_12_99), .C1 (n_8_99), .C2 (n_4_98) );
AOI211_X1 g_24_99 (.ZN (n_24_99), .A (n_20_99), .B (n_14_100), .C1 (n_10_100), .C2 (n_5_100) );
AOI211_X1 g_26_100 (.ZN (n_26_100), .A (n_22_100), .B (n_16_99), .C1 (n_12_99), .C2 (n_6_98) );
AOI211_X1 g_28_99 (.ZN (n_28_99), .A (n_24_99), .B (n_18_100), .C1 (n_14_100), .C2 (n_8_99) );
AOI211_X1 g_30_100 (.ZN (n_30_100), .A (n_26_100), .B (n_20_99), .C1 (n_16_99), .C2 (n_10_100) );
AOI211_X1 g_32_99 (.ZN (n_32_99), .A (n_28_99), .B (n_22_100), .C1 (n_18_100), .C2 (n_12_99) );
AOI211_X1 g_34_100 (.ZN (n_34_100), .A (n_30_100), .B (n_24_99), .C1 (n_20_99), .C2 (n_14_100) );
AOI211_X1 g_36_99 (.ZN (n_36_99), .A (n_32_99), .B (n_26_100), .C1 (n_22_100), .C2 (n_16_99) );
AOI211_X1 g_38_100 (.ZN (n_38_100), .A (n_34_100), .B (n_28_99), .C1 (n_24_99), .C2 (n_18_100) );
AOI211_X1 g_40_99 (.ZN (n_40_99), .A (n_36_99), .B (n_30_100), .C1 (n_26_100), .C2 (n_20_99) );
AOI211_X1 g_42_100 (.ZN (n_42_100), .A (n_38_100), .B (n_32_99), .C1 (n_28_99), .C2 (n_22_100) );
AOI211_X1 g_44_99 (.ZN (n_44_99), .A (n_40_99), .B (n_34_100), .C1 (n_30_100), .C2 (n_24_99) );
AOI211_X1 g_46_100 (.ZN (n_46_100), .A (n_42_100), .B (n_36_99), .C1 (n_32_99), .C2 (n_26_100) );
AOI211_X1 g_48_99 (.ZN (n_48_99), .A (n_44_99), .B (n_38_100), .C1 (n_34_100), .C2 (n_28_99) );
AOI211_X1 g_50_100 (.ZN (n_50_100), .A (n_46_100), .B (n_40_99), .C1 (n_36_99), .C2 (n_30_100) );
AOI211_X1 g_52_99 (.ZN (n_52_99), .A (n_48_99), .B (n_42_100), .C1 (n_38_100), .C2 (n_32_99) );
AOI211_X1 g_54_100 (.ZN (n_54_100), .A (n_50_100), .B (n_44_99), .C1 (n_40_99), .C2 (n_34_100) );
AOI211_X1 g_56_99 (.ZN (n_56_99), .A (n_52_99), .B (n_46_100), .C1 (n_42_100), .C2 (n_36_99) );
AOI211_X1 g_58_100 (.ZN (n_58_100), .A (n_54_100), .B (n_48_99), .C1 (n_44_99), .C2 (n_38_100) );
AOI211_X1 g_60_99 (.ZN (n_60_99), .A (n_56_99), .B (n_50_100), .C1 (n_46_100), .C2 (n_40_99) );
AOI211_X1 g_62_100 (.ZN (n_62_100), .A (n_58_100), .B (n_52_99), .C1 (n_48_99), .C2 (n_42_100) );
AOI211_X1 g_64_99 (.ZN (n_64_99), .A (n_60_99), .B (n_54_100), .C1 (n_50_100), .C2 (n_44_99) );
AOI211_X1 g_66_100 (.ZN (n_66_100), .A (n_62_100), .B (n_56_99), .C1 (n_52_99), .C2 (n_46_100) );
AOI211_X1 g_68_99 (.ZN (n_68_99), .A (n_64_99), .B (n_58_100), .C1 (n_54_100), .C2 (n_48_99) );
AOI211_X1 g_70_100 (.ZN (n_70_100), .A (n_66_100), .B (n_60_99), .C1 (n_56_99), .C2 (n_50_100) );
AOI211_X1 g_72_99 (.ZN (n_72_99), .A (n_68_99), .B (n_62_100), .C1 (n_58_100), .C2 (n_52_99) );
AOI211_X1 g_74_100 (.ZN (n_74_100), .A (n_70_100), .B (n_64_99), .C1 (n_60_99), .C2 (n_54_100) );
AOI211_X1 g_76_99 (.ZN (n_76_99), .A (n_72_99), .B (n_66_100), .C1 (n_62_100), .C2 (n_56_99) );
AOI211_X1 g_78_100 (.ZN (n_78_100), .A (n_74_100), .B (n_68_99), .C1 (n_64_99), .C2 (n_58_100) );
AOI211_X1 g_80_99 (.ZN (n_80_99), .A (n_76_99), .B (n_70_100), .C1 (n_66_100), .C2 (n_60_99) );
AOI211_X1 g_82_100 (.ZN (n_82_100), .A (n_78_100), .B (n_72_99), .C1 (n_68_99), .C2 (n_62_100) );
AOI211_X1 g_84_99 (.ZN (n_84_99), .A (n_80_99), .B (n_74_100), .C1 (n_70_100), .C2 (n_64_99) );
AOI211_X1 g_86_100 (.ZN (n_86_100), .A (n_82_100), .B (n_76_99), .C1 (n_72_99), .C2 (n_66_100) );
AOI211_X1 g_88_99 (.ZN (n_88_99), .A (n_84_99), .B (n_78_100), .C1 (n_74_100), .C2 (n_68_99) );
AOI211_X1 g_90_100 (.ZN (n_90_100), .A (n_86_100), .B (n_80_99), .C1 (n_76_99), .C2 (n_70_100) );
AOI211_X1 g_92_99 (.ZN (n_92_99), .A (n_88_99), .B (n_82_100), .C1 (n_78_100), .C2 (n_72_99) );
AOI211_X1 g_94_100 (.ZN (n_94_100), .A (n_90_100), .B (n_84_99), .C1 (n_80_99), .C2 (n_74_100) );
AOI211_X1 g_96_99 (.ZN (n_96_99), .A (n_92_99), .B (n_86_100), .C1 (n_82_100), .C2 (n_76_99) );
AOI211_X1 g_98_100 (.ZN (n_98_100), .A (n_94_100), .B (n_88_99), .C1 (n_84_99), .C2 (n_78_100) );
AOI211_X1 g_100_99 (.ZN (n_100_99), .A (n_96_99), .B (n_90_100), .C1 (n_86_100), .C2 (n_80_99) );
AOI211_X1 g_98_98 (.ZN (n_98_98), .A (n_98_100), .B (n_92_99), .C1 (n_88_99), .C2 (n_82_100) );
AOI211_X1 g_100_97 (.ZN (n_100_97), .A (n_100_99), .B (n_94_100), .C1 (n_90_100), .C2 (n_84_99) );
AOI211_X1 g_99_99 (.ZN (n_99_99), .A (n_98_98), .B (n_96_99), .C1 (n_92_99), .C2 (n_86_100) );
AOI211_X1 g_97_100 (.ZN (n_97_100), .A (n_100_97), .B (n_98_100), .C1 (n_94_100), .C2 (n_88_99) );
AOI211_X1 g_95_99 (.ZN (n_95_99), .A (n_99_99), .B (n_100_99), .C1 (n_96_99), .C2 (n_90_100) );
AOI211_X1 g_93_100 (.ZN (n_93_100), .A (n_97_100), .B (n_98_98), .C1 (n_98_100), .C2 (n_92_99) );
AOI211_X1 g_94_98 (.ZN (n_94_98), .A (n_95_99), .B (n_100_97), .C1 (n_100_99), .C2 (n_94_100) );
AOI211_X1 g_96_97 (.ZN (n_96_97), .A (n_93_100), .B (n_99_99), .C1 (n_98_98), .C2 (n_96_99) );
AOI211_X1 g_98_96 (.ZN (n_98_96), .A (n_94_98), .B (n_97_100), .C1 (n_100_97), .C2 (n_98_100) );
AOI211_X1 g_100_95 (.ZN (n_100_95), .A (n_96_97), .B (n_95_99), .C1 (n_99_99), .C2 (n_100_99) );
AOI211_X1 g_99_97 (.ZN (n_99_97), .A (n_98_96), .B (n_93_100), .C1 (n_97_100), .C2 (n_98_98) );
AOI211_X1 g_97_98 (.ZN (n_97_98), .A (n_100_95), .B (n_94_98), .C1 (n_95_99), .C2 (n_100_97) );
AOI211_X1 g_96_100 (.ZN (n_96_100), .A (n_99_97), .B (n_96_97), .C1 (n_93_100), .C2 (n_99_99) );
AOI211_X1 g_98_99 (.ZN (n_98_99), .A (n_97_98), .B (n_98_96), .C1 (n_94_98), .C2 (n_97_100) );
AOI211_X1 g_100_100 (.ZN (n_100_100), .A (n_96_100), .B (n_100_95), .C1 (n_96_97), .C2 (n_95_99) );
AOI211_X1 g_99_98 (.ZN (n_99_98), .A (n_98_99), .B (n_99_97), .C1 (n_98_96), .C2 (n_93_100) );
AOI211_X1 g_100_96 (.ZN (n_100_96), .A (n_100_100), .B (n_97_98), .C1 (n_100_95), .C2 (n_94_98) );
AOI211_X1 g_99_94 (.ZN (n_99_94), .A (n_99_98), .B (n_96_100), .C1 (n_99_97), .C2 (n_96_97) );
AOI211_X1 g_100_92 (.ZN (n_100_92), .A (n_100_96), .B (n_98_99), .C1 (n_97_98), .C2 (n_98_96) );
AOI211_X1 g_99_90 (.ZN (n_99_90), .A (n_99_94), .B (n_100_100), .C1 (n_96_100), .C2 (n_100_95) );
AOI211_X1 g_100_88 (.ZN (n_100_88), .A (n_100_92), .B (n_99_98), .C1 (n_98_99), .C2 (n_99_97) );
AOI211_X1 g_99_86 (.ZN (n_99_86), .A (n_99_90), .B (n_100_96), .C1 (n_100_100), .C2 (n_97_98) );
AOI211_X1 g_100_84 (.ZN (n_100_84), .A (n_100_88), .B (n_99_94), .C1 (n_99_98), .C2 (n_96_100) );
AOI211_X1 g_99_82 (.ZN (n_99_82), .A (n_99_86), .B (n_100_92), .C1 (n_100_96), .C2 (n_98_99) );
AOI211_X1 g_100_80 (.ZN (n_100_80), .A (n_100_84), .B (n_99_90), .C1 (n_99_94), .C2 (n_100_100) );
AOI211_X1 g_99_78 (.ZN (n_99_78), .A (n_99_82), .B (n_100_88), .C1 (n_100_92), .C2 (n_99_98) );
AOI211_X1 g_100_76 (.ZN (n_100_76), .A (n_100_80), .B (n_99_86), .C1 (n_99_90), .C2 (n_100_96) );
AOI211_X1 g_99_74 (.ZN (n_99_74), .A (n_99_78), .B (n_100_84), .C1 (n_100_88), .C2 (n_99_94) );
AOI211_X1 g_100_72 (.ZN (n_100_72), .A (n_100_76), .B (n_99_82), .C1 (n_99_86), .C2 (n_100_92) );
AOI211_X1 g_99_70 (.ZN (n_99_70), .A (n_99_74), .B (n_100_80), .C1 (n_100_84), .C2 (n_99_90) );
AOI211_X1 g_98_68 (.ZN (n_98_68), .A (n_100_72), .B (n_99_78), .C1 (n_99_82), .C2 (n_100_88) );
AOI211_X1 g_97_66 (.ZN (n_97_66), .A (n_99_70), .B (n_100_76), .C1 (n_100_80), .C2 (n_99_86) );
AOI211_X1 g_96_64 (.ZN (n_96_64), .A (n_98_68), .B (n_99_74), .C1 (n_99_78), .C2 (n_100_84) );
AOI211_X1 g_95_62 (.ZN (n_95_62), .A (n_97_66), .B (n_100_72), .C1 (n_100_76), .C2 (n_99_82) );
AOI211_X1 g_97_61 (.ZN (n_97_61), .A (n_96_64), .B (n_99_70), .C1 (n_99_74), .C2 (n_100_80) );
AOI211_X1 g_96_59 (.ZN (n_96_59), .A (n_95_62), .B (n_98_68), .C1 (n_100_72), .C2 (n_99_78) );
AOI211_X1 g_95_57 (.ZN (n_95_57), .A (n_97_61), .B (n_97_66), .C1 (n_99_70), .C2 (n_100_76) );
AOI211_X1 g_93_56 (.ZN (n_93_56), .A (n_96_59), .B (n_96_64), .C1 (n_98_68), .C2 (n_99_74) );
AOI211_X1 g_91_57 (.ZN (n_91_57), .A (n_95_57), .B (n_95_62), .C1 (n_97_66), .C2 (n_100_72) );
AOI211_X1 g_93_58 (.ZN (n_93_58), .A (n_93_56), .B (n_97_61), .C1 (n_96_64), .C2 (n_99_70) );
AOI211_X1 g_94_60 (.ZN (n_94_60), .A (n_91_57), .B (n_96_59), .C1 (n_95_62), .C2 (n_98_68) );
AOI211_X1 g_92_59 (.ZN (n_92_59), .A (n_93_58), .B (n_95_57), .C1 (n_97_61), .C2 (n_97_66) );
AOI211_X1 g_94_58 (.ZN (n_94_58), .A (n_94_60), .B (n_93_56), .C1 (n_96_59), .C2 (n_96_64) );
AOI211_X1 g_95_60 (.ZN (n_95_60), .A (n_92_59), .B (n_91_57), .C1 (n_95_57), .C2 (n_95_62) );
AOI211_X1 g_93_59 (.ZN (n_93_59), .A (n_94_58), .B (n_93_58), .C1 (n_93_56), .C2 (n_97_61) );
AOI211_X1 g_91_58 (.ZN (n_91_58), .A (n_95_60), .B (n_94_60), .C1 (n_91_57), .C2 (n_96_59) );
AOI211_X1 g_89_57 (.ZN (n_89_57), .A (n_93_59), .B (n_92_59), .C1 (n_93_58), .C2 (n_95_57) );
AOI211_X1 g_87_58 (.ZN (n_87_58), .A (n_91_58), .B (n_94_58), .C1 (n_94_60), .C2 (n_93_56) );
AOI211_X1 g_85_59 (.ZN (n_85_59), .A (n_89_57), .B (n_95_60), .C1 (n_92_59), .C2 (n_91_57) );
AOI211_X1 g_83_60 (.ZN (n_83_60), .A (n_87_58), .B (n_93_59), .C1 (n_94_58), .C2 (n_93_58) );
AOI211_X1 g_81_61 (.ZN (n_81_61), .A (n_85_59), .B (n_91_58), .C1 (n_95_60), .C2 (n_94_60) );
AOI211_X1 g_79_62 (.ZN (n_79_62), .A (n_83_60), .B (n_89_57), .C1 (n_93_59), .C2 (n_92_59) );
AOI211_X1 g_80_60 (.ZN (n_80_60), .A (n_81_61), .B (n_87_58), .C1 (n_91_58), .C2 (n_94_58) );
AOI211_X1 g_78_61 (.ZN (n_78_61), .A (n_79_62), .B (n_85_59), .C1 (n_89_57), .C2 (n_95_60) );
AOI211_X1 g_76_62 (.ZN (n_76_62), .A (n_80_60), .B (n_83_60), .C1 (n_87_58), .C2 (n_93_59) );
AOI211_X1 g_74_63 (.ZN (n_74_63), .A (n_78_61), .B (n_81_61), .C1 (n_85_59), .C2 (n_91_58) );
AOI211_X1 g_72_64 (.ZN (n_72_64), .A (n_76_62), .B (n_79_62), .C1 (n_83_60), .C2 (n_89_57) );
AOI211_X1 g_70_65 (.ZN (n_70_65), .A (n_74_63), .B (n_80_60), .C1 (n_81_61), .C2 (n_87_58) );
AOI211_X1 g_69_67 (.ZN (n_69_67), .A (n_72_64), .B (n_78_61), .C1 (n_79_62), .C2 (n_85_59) );
AOI211_X1 g_67_68 (.ZN (n_67_68), .A (n_70_65), .B (n_76_62), .C1 (n_80_60), .C2 (n_83_60) );
AOI211_X1 g_66_70 (.ZN (n_66_70), .A (n_69_67), .B (n_74_63), .C1 (n_78_61), .C2 (n_81_61) );
AOI211_X1 g_65_68 (.ZN (n_65_68), .A (n_67_68), .B (n_72_64), .C1 (n_76_62), .C2 (n_79_62) );
AOI211_X1 g_67_67 (.ZN (n_67_67), .A (n_66_70), .B (n_70_65), .C1 (n_74_63), .C2 (n_80_60) );
AOI211_X1 g_69_66 (.ZN (n_69_66), .A (n_65_68), .B (n_69_67), .C1 (n_72_64), .C2 (n_78_61) );
AOI211_X1 g_71_65 (.ZN (n_71_65), .A (n_67_67), .B (n_67_68), .C1 (n_70_65), .C2 (n_76_62) );
AOI211_X1 g_73_64 (.ZN (n_73_64), .A (n_69_66), .B (n_66_70), .C1 (n_69_67), .C2 (n_74_63) );
AOI211_X1 g_72_66 (.ZN (n_72_66), .A (n_71_65), .B (n_65_68), .C1 (n_67_68), .C2 (n_72_64) );
AOI211_X1 g_74_65 (.ZN (n_74_65), .A (n_73_64), .B (n_67_67), .C1 (n_66_70), .C2 (n_70_65) );
AOI211_X1 g_76_64 (.ZN (n_76_64), .A (n_72_66), .B (n_69_66), .C1 (n_65_68), .C2 (n_69_67) );
AOI211_X1 g_78_63 (.ZN (n_78_63), .A (n_74_65), .B (n_71_65), .C1 (n_67_67), .C2 (n_67_68) );
AOI211_X1 g_80_62 (.ZN (n_80_62), .A (n_76_64), .B (n_73_64), .C1 (n_69_66), .C2 (n_66_70) );
AOI211_X1 g_82_61 (.ZN (n_82_61), .A (n_78_63), .B (n_72_66), .C1 (n_71_65), .C2 (n_65_68) );
AOI211_X1 g_84_60 (.ZN (n_84_60), .A (n_80_62), .B (n_74_65), .C1 (n_73_64), .C2 (n_67_67) );
AOI211_X1 g_86_59 (.ZN (n_86_59), .A (n_82_61), .B (n_76_64), .C1 (n_72_66), .C2 (n_69_66) );
AOI211_X1 g_88_58 (.ZN (n_88_58), .A (n_84_60), .B (n_78_63), .C1 (n_74_65), .C2 (n_71_65) );
AOI211_X1 g_90_57 (.ZN (n_90_57), .A (n_86_59), .B (n_80_62), .C1 (n_76_64), .C2 (n_73_64) );
AOI211_X1 g_89_59 (.ZN (n_89_59), .A (n_88_58), .B (n_82_61), .C1 (n_78_63), .C2 (n_72_66) );
AOI211_X1 g_87_60 (.ZN (n_87_60), .A (n_90_57), .B (n_84_60), .C1 (n_80_62), .C2 (n_74_65) );
AOI211_X1 g_85_61 (.ZN (n_85_61), .A (n_89_59), .B (n_86_59), .C1 (n_82_61), .C2 (n_76_64) );
AOI211_X1 g_83_62 (.ZN (n_83_62), .A (n_87_60), .B (n_88_58), .C1 (n_84_60), .C2 (n_78_63) );
AOI211_X1 g_81_63 (.ZN (n_81_63), .A (n_85_61), .B (n_90_57), .C1 (n_86_59), .C2 (n_80_62) );
AOI211_X1 g_80_61 (.ZN (n_80_61), .A (n_83_62), .B (n_89_59), .C1 (n_88_58), .C2 (n_82_61) );
AOI211_X1 g_78_62 (.ZN (n_78_62), .A (n_81_63), .B (n_87_60), .C1 (n_90_57), .C2 (n_84_60) );
AOI211_X1 g_76_63 (.ZN (n_76_63), .A (n_80_61), .B (n_85_61), .C1 (n_89_59), .C2 (n_86_59) );
AOI211_X1 g_74_64 (.ZN (n_74_64), .A (n_78_62), .B (n_83_62), .C1 (n_87_60), .C2 (n_88_58) );
AOI211_X1 g_72_65 (.ZN (n_72_65), .A (n_76_63), .B (n_81_63), .C1 (n_85_61), .C2 (n_90_57) );
AOI211_X1 g_70_66 (.ZN (n_70_66), .A (n_74_64), .B (n_80_61), .C1 (n_83_62), .C2 (n_89_59) );
AOI211_X1 g_68_67 (.ZN (n_68_67), .A (n_72_65), .B (n_78_62), .C1 (n_81_63), .C2 (n_87_60) );
AOI211_X1 g_66_68 (.ZN (n_66_68), .A (n_70_66), .B (n_76_63), .C1 (n_80_61), .C2 (n_85_61) );
AOI211_X1 g_64_69 (.ZN (n_64_69), .A (n_68_67), .B (n_74_64), .C1 (n_78_62), .C2 (n_83_62) );
AOI211_X1 g_62_68 (.ZN (n_62_68), .A (n_66_68), .B (n_72_65), .C1 (n_76_63), .C2 (n_81_63) );
AOI211_X1 g_60_69 (.ZN (n_60_69), .A (n_64_69), .B (n_70_66), .C1 (n_74_64), .C2 (n_80_61) );
AOI211_X1 g_58_70 (.ZN (n_58_70), .A (n_62_68), .B (n_68_67), .C1 (n_72_65), .C2 (n_78_62) );
AOI211_X1 g_56_71 (.ZN (n_56_71), .A (n_60_69), .B (n_66_68), .C1 (n_70_66), .C2 (n_76_63) );
AOI211_X1 g_54_72 (.ZN (n_54_72), .A (n_58_70), .B (n_64_69), .C1 (n_68_67), .C2 (n_74_64) );
AOI211_X1 g_52_73 (.ZN (n_52_73), .A (n_56_71), .B (n_62_68), .C1 (n_66_68), .C2 (n_72_65) );
AOI211_X1 g_50_74 (.ZN (n_50_74), .A (n_54_72), .B (n_60_69), .C1 (n_64_69), .C2 (n_70_66) );
AOI211_X1 g_48_75 (.ZN (n_48_75), .A (n_52_73), .B (n_58_70), .C1 (n_62_68), .C2 (n_68_67) );
AOI211_X1 g_47_73 (.ZN (n_47_73), .A (n_50_74), .B (n_56_71), .C1 (n_60_69), .C2 (n_66_68) );
AOI211_X1 g_45_74 (.ZN (n_45_74), .A (n_48_75), .B (n_54_72), .C1 (n_58_70), .C2 (n_64_69) );
AOI211_X1 g_43_75 (.ZN (n_43_75), .A (n_47_73), .B (n_52_73), .C1 (n_56_71), .C2 (n_62_68) );
AOI211_X1 g_41_76 (.ZN (n_41_76), .A (n_45_74), .B (n_50_74), .C1 (n_54_72), .C2 (n_60_69) );
AOI211_X1 g_39_77 (.ZN (n_39_77), .A (n_43_75), .B (n_48_75), .C1 (n_52_73), .C2 (n_58_70) );
AOI211_X1 g_37_78 (.ZN (n_37_78), .A (n_41_76), .B (n_47_73), .C1 (n_50_74), .C2 (n_56_71) );
AOI211_X1 g_35_79 (.ZN (n_35_79), .A (n_39_77), .B (n_45_74), .C1 (n_48_75), .C2 (n_54_72) );
AOI211_X1 g_33_80 (.ZN (n_33_80), .A (n_37_78), .B (n_43_75), .C1 (n_47_73), .C2 (n_52_73) );
AOI211_X1 g_31_81 (.ZN (n_31_81), .A (n_35_79), .B (n_41_76), .C1 (n_45_74), .C2 (n_50_74) );
AOI211_X1 g_29_82 (.ZN (n_29_82), .A (n_33_80), .B (n_39_77), .C1 (n_43_75), .C2 (n_48_75) );
AOI211_X1 g_27_83 (.ZN (n_27_83), .A (n_31_81), .B (n_37_78), .C1 (n_41_76), .C2 (n_47_73) );
AOI211_X1 g_25_84 (.ZN (n_25_84), .A (n_29_82), .B (n_35_79), .C1 (n_39_77), .C2 (n_45_74) );
AOI211_X1 g_26_82 (.ZN (n_26_82), .A (n_27_83), .B (n_33_80), .C1 (n_37_78), .C2 (n_43_75) );
AOI211_X1 g_24_83 (.ZN (n_24_83), .A (n_25_84), .B (n_31_81), .C1 (n_35_79), .C2 (n_41_76) );
AOI211_X1 g_22_84 (.ZN (n_22_84), .A (n_26_82), .B (n_29_82), .C1 (n_33_80), .C2 (n_39_77) );
AOI211_X1 g_20_85 (.ZN (n_20_85), .A (n_24_83), .B (n_27_83), .C1 (n_31_81), .C2 (n_37_78) );
AOI211_X1 g_18_86 (.ZN (n_18_86), .A (n_22_84), .B (n_25_84), .C1 (n_29_82), .C2 (n_35_79) );
AOI211_X1 g_16_87 (.ZN (n_16_87), .A (n_20_85), .B (n_26_82), .C1 (n_27_83), .C2 (n_33_80) );
AOI211_X1 g_14_88 (.ZN (n_14_88), .A (n_18_86), .B (n_24_83), .C1 (n_25_84), .C2 (n_31_81) );
AOI211_X1 g_12_89 (.ZN (n_12_89), .A (n_16_87), .B (n_22_84), .C1 (n_26_82), .C2 (n_29_82) );
AOI211_X1 g_10_90 (.ZN (n_10_90), .A (n_14_88), .B (n_20_85), .C1 (n_24_83), .C2 (n_27_83) );
AOI211_X1 g_8_91 (.ZN (n_8_91), .A (n_12_89), .B (n_18_86), .C1 (n_22_84), .C2 (n_25_84) );
AOI211_X1 g_7_93 (.ZN (n_7_93), .A (n_10_90), .B (n_16_87), .C1 (n_20_85), .C2 (n_26_82) );
AOI211_X1 g_9_92 (.ZN (n_9_92), .A (n_8_91), .B (n_14_88), .C1 (n_18_86), .C2 (n_24_83) );
AOI211_X1 g_11_91 (.ZN (n_11_91), .A (n_7_93), .B (n_12_89), .C1 (n_16_87), .C2 (n_22_84) );
AOI211_X1 g_13_90 (.ZN (n_13_90), .A (n_9_92), .B (n_10_90), .C1 (n_14_88), .C2 (n_20_85) );
AOI211_X1 g_15_89 (.ZN (n_15_89), .A (n_11_91), .B (n_8_91), .C1 (n_12_89), .C2 (n_18_86) );
AOI211_X1 g_17_88 (.ZN (n_17_88), .A (n_13_90), .B (n_7_93), .C1 (n_10_90), .C2 (n_16_87) );
AOI211_X1 g_19_87 (.ZN (n_19_87), .A (n_15_89), .B (n_9_92), .C1 (n_8_91), .C2 (n_14_88) );
AOI211_X1 g_21_86 (.ZN (n_21_86), .A (n_17_88), .B (n_11_91), .C1 (n_7_93), .C2 (n_12_89) );
AOI211_X1 g_23_85 (.ZN (n_23_85), .A (n_19_87), .B (n_13_90), .C1 (n_9_92), .C2 (n_10_90) );
AOI211_X1 g_22_87 (.ZN (n_22_87), .A (n_21_86), .B (n_15_89), .C1 (n_11_91), .C2 (n_8_91) );
AOI211_X1 g_20_86 (.ZN (n_20_86), .A (n_23_85), .B (n_17_88), .C1 (n_13_90), .C2 (n_7_93) );
AOI211_X1 g_18_87 (.ZN (n_18_87), .A (n_22_87), .B (n_19_87), .C1 (n_15_89), .C2 (n_9_92) );
AOI211_X1 g_20_88 (.ZN (n_20_88), .A (n_20_86), .B (n_21_86), .C1 (n_17_88), .C2 (n_11_91) );
AOI211_X1 g_18_89 (.ZN (n_18_89), .A (n_18_87), .B (n_23_85), .C1 (n_19_87), .C2 (n_13_90) );
AOI211_X1 g_16_90 (.ZN (n_16_90), .A (n_20_88), .B (n_22_87), .C1 (n_21_86), .C2 (n_15_89) );
AOI211_X1 g_14_91 (.ZN (n_14_91), .A (n_18_89), .B (n_20_86), .C1 (n_23_85), .C2 (n_17_88) );
AOI211_X1 g_12_92 (.ZN (n_12_92), .A (n_16_90), .B (n_18_87), .C1 (n_22_87), .C2 (n_19_87) );
AOI211_X1 g_10_93 (.ZN (n_10_93), .A (n_14_91), .B (n_20_88), .C1 (n_20_86), .C2 (n_21_86) );
AOI211_X1 g_8_94 (.ZN (n_8_94), .A (n_12_92), .B (n_18_89), .C1 (n_18_87), .C2 (n_23_85) );
AOI211_X1 g_6_95 (.ZN (n_6_95), .A (n_10_93), .B (n_16_90), .C1 (n_20_88), .C2 (n_22_87) );
AOI211_X1 g_5_97 (.ZN (n_5_97), .A (n_8_94), .B (n_14_91), .C1 (n_18_89), .C2 (n_20_86) );
AOI211_X1 g_7_96 (.ZN (n_7_96), .A (n_6_95), .B (n_12_92), .C1 (n_16_90), .C2 (n_18_87) );
AOI211_X1 g_9_95 (.ZN (n_9_95), .A (n_5_97), .B (n_10_93), .C1 (n_14_91), .C2 (n_20_88) );
AOI211_X1 g_8_97 (.ZN (n_8_97), .A (n_7_96), .B (n_8_94), .C1 (n_12_92), .C2 (n_18_89) );
AOI211_X1 g_7_95 (.ZN (n_7_95), .A (n_9_95), .B (n_6_95), .C1 (n_10_93), .C2 (n_16_90) );
AOI211_X1 g_6_97 (.ZN (n_6_97), .A (n_8_97), .B (n_5_97), .C1 (n_8_94), .C2 (n_14_91) );
AOI211_X1 g_7_99 (.ZN (n_7_99), .A (n_7_95), .B (n_7_96), .C1 (n_6_95), .C2 (n_12_92) );
AOI211_X1 g_9_100 (.ZN (n_9_100), .A (n_6_97), .B (n_9_95), .C1 (n_5_97), .C2 (n_10_93) );
AOI211_X1 g_10_98 (.ZN (n_10_98), .A (n_7_99), .B (n_8_97), .C1 (n_7_96), .C2 (n_8_94) );
AOI211_X1 g_9_96 (.ZN (n_9_96), .A (n_9_100), .B (n_7_95), .C1 (n_9_95), .C2 (n_6_95) );
AOI211_X1 g_7_97 (.ZN (n_7_97), .A (n_10_98), .B (n_6_97), .C1 (n_8_97), .C2 (n_5_97) );
AOI211_X1 g_6_99 (.ZN (n_6_99), .A (n_9_96), .B (n_7_99), .C1 (n_7_95), .C2 (n_7_96) );
AOI211_X1 g_8_98 (.ZN (n_8_98), .A (n_7_97), .B (n_9_100), .C1 (n_6_97), .C2 (n_9_95) );
AOI211_X1 g_10_97 (.ZN (n_10_97), .A (n_6_99), .B (n_10_98), .C1 (n_7_99), .C2 (n_8_97) );
AOI211_X1 g_8_96 (.ZN (n_8_96), .A (n_8_98), .B (n_9_96), .C1 (n_9_100), .C2 (n_7_95) );
AOI211_X1 g_7_98 (.ZN (n_7_98), .A (n_10_97), .B (n_7_97), .C1 (n_10_98), .C2 (n_6_97) );
AOI211_X1 g_8_100 (.ZN (n_8_100), .A (n_8_96), .B (n_6_99), .C1 (n_9_96), .C2 (n_7_99) );
AOI211_X1 g_9_98 (.ZN (n_9_98), .A (n_7_98), .B (n_8_98), .C1 (n_7_97), .C2 (n_9_100) );
AOI211_X1 g_11_99 (.ZN (n_11_99), .A (n_8_100), .B (n_10_97), .C1 (n_6_99), .C2 (n_10_98) );
AOI211_X1 g_13_100 (.ZN (n_13_100), .A (n_9_98), .B (n_8_96), .C1 (n_8_98), .C2 (n_9_96) );
AOI211_X1 g_14_98 (.ZN (n_14_98), .A (n_11_99), .B (n_7_98), .C1 (n_10_97), .C2 (n_7_97) );
AOI211_X1 g_12_97 (.ZN (n_12_97), .A (n_13_100), .B (n_8_100), .C1 (n_8_96), .C2 (n_6_99) );
AOI211_X1 g_11_95 (.ZN (n_11_95), .A (n_14_98), .B (n_9_98), .C1 (n_7_98), .C2 (n_8_98) );
AOI211_X1 g_9_94 (.ZN (n_9_94), .A (n_12_97), .B (n_11_99), .C1 (n_8_100), .C2 (n_10_97) );
AOI211_X1 g_10_92 (.ZN (n_10_92), .A (n_11_95), .B (n_13_100), .C1 (n_9_98), .C2 (n_8_96) );
AOI211_X1 g_12_91 (.ZN (n_12_91), .A (n_9_94), .B (n_14_98), .C1 (n_11_99), .C2 (n_7_98) );
AOI211_X1 g_14_90 (.ZN (n_14_90), .A (n_10_92), .B (n_12_97), .C1 (n_13_100), .C2 (n_8_100) );
AOI211_X1 g_16_89 (.ZN (n_16_89), .A (n_12_91), .B (n_11_95), .C1 (n_14_98), .C2 (n_9_98) );
AOI211_X1 g_18_88 (.ZN (n_18_88), .A (n_14_90), .B (n_9_94), .C1 (n_12_97), .C2 (n_11_99) );
AOI211_X1 g_20_87 (.ZN (n_20_87), .A (n_16_89), .B (n_10_92), .C1 (n_11_95), .C2 (n_13_100) );
AOI211_X1 g_22_86 (.ZN (n_22_86), .A (n_18_88), .B (n_12_91), .C1 (n_9_94), .C2 (n_14_98) );
AOI211_X1 g_24_85 (.ZN (n_24_85), .A (n_20_87), .B (n_14_90), .C1 (n_10_92), .C2 (n_12_97) );
AOI211_X1 g_26_84 (.ZN (n_26_84), .A (n_22_86), .B (n_16_89), .C1 (n_12_91), .C2 (n_11_95) );
AOI211_X1 g_28_83 (.ZN (n_28_83), .A (n_24_85), .B (n_18_88), .C1 (n_14_90), .C2 (n_9_94) );
AOI211_X1 g_30_82 (.ZN (n_30_82), .A (n_26_84), .B (n_20_87), .C1 (n_16_89), .C2 (n_10_92) );
AOI211_X1 g_32_81 (.ZN (n_32_81), .A (n_28_83), .B (n_22_86), .C1 (n_18_88), .C2 (n_12_91) );
AOI211_X1 g_34_80 (.ZN (n_34_80), .A (n_30_82), .B (n_24_85), .C1 (n_20_87), .C2 (n_14_90) );
AOI211_X1 g_36_79 (.ZN (n_36_79), .A (n_32_81), .B (n_26_84), .C1 (n_22_86), .C2 (n_16_89) );
AOI211_X1 g_38_78 (.ZN (n_38_78), .A (n_34_80), .B (n_28_83), .C1 (n_24_85), .C2 (n_18_88) );
AOI211_X1 g_37_80 (.ZN (n_37_80), .A (n_36_79), .B (n_30_82), .C1 (n_26_84), .C2 (n_20_87) );
AOI211_X1 g_39_79 (.ZN (n_39_79), .A (n_38_78), .B (n_32_81), .C1 (n_28_83), .C2 (n_22_86) );
AOI211_X1 g_41_78 (.ZN (n_41_78), .A (n_37_80), .B (n_34_80), .C1 (n_30_82), .C2 (n_24_85) );
AOI211_X1 g_43_77 (.ZN (n_43_77), .A (n_39_79), .B (n_36_79), .C1 (n_32_81), .C2 (n_26_84) );
AOI211_X1 g_45_76 (.ZN (n_45_76), .A (n_41_78), .B (n_38_78), .C1 (n_34_80), .C2 (n_28_83) );
AOI211_X1 g_47_75 (.ZN (n_47_75), .A (n_43_77), .B (n_37_80), .C1 (n_36_79), .C2 (n_30_82) );
AOI211_X1 g_49_74 (.ZN (n_49_74), .A (n_45_76), .B (n_39_79), .C1 (n_38_78), .C2 (n_32_81) );
AOI211_X1 g_51_73 (.ZN (n_51_73), .A (n_47_75), .B (n_41_78), .C1 (n_37_80), .C2 (n_34_80) );
AOI211_X1 g_53_72 (.ZN (n_53_72), .A (n_49_74), .B (n_43_77), .C1 (n_39_79), .C2 (n_36_79) );
AOI211_X1 g_55_71 (.ZN (n_55_71), .A (n_51_73), .B (n_45_76), .C1 (n_41_78), .C2 (n_38_78) );
AOI211_X1 g_57_70 (.ZN (n_57_70), .A (n_53_72), .B (n_47_75), .C1 (n_43_77), .C2 (n_37_80) );
AOI211_X1 g_59_69 (.ZN (n_59_69), .A (n_55_71), .B (n_49_74), .C1 (n_45_76), .C2 (n_39_79) );
AOI211_X1 g_61_68 (.ZN (n_61_68), .A (n_57_70), .B (n_51_73), .C1 (n_47_75), .C2 (n_41_78) );
AOI211_X1 g_62_70 (.ZN (n_62_70), .A (n_59_69), .B (n_53_72), .C1 (n_49_74), .C2 (n_43_77) );
AOI211_X1 g_60_71 (.ZN (n_60_71), .A (n_61_68), .B (n_55_71), .C1 (n_51_73), .C2 (n_45_76) );
AOI211_X1 g_58_72 (.ZN (n_58_72), .A (n_62_70), .B (n_57_70), .C1 (n_53_72), .C2 (n_47_75) );
AOI211_X1 g_56_73 (.ZN (n_56_73), .A (n_60_71), .B (n_59_69), .C1 (n_55_71), .C2 (n_49_74) );
AOI211_X1 g_57_71 (.ZN (n_57_71), .A (n_58_72), .B (n_61_68), .C1 (n_57_70), .C2 (n_51_73) );
AOI211_X1 g_58_69 (.ZN (n_58_69), .A (n_56_73), .B (n_62_70), .C1 (n_59_69), .C2 (n_53_72) );
AOI211_X1 g_56_70 (.ZN (n_56_70), .A (n_57_71), .B (n_60_71), .C1 (n_61_68), .C2 (n_55_71) );
AOI211_X1 g_54_71 (.ZN (n_54_71), .A (n_58_69), .B (n_58_72), .C1 (n_62_70), .C2 (n_57_70) );
AOI211_X1 g_52_72 (.ZN (n_52_72), .A (n_56_70), .B (n_56_73), .C1 (n_60_71), .C2 (n_59_69) );
AOI211_X1 g_50_73 (.ZN (n_50_73), .A (n_54_71), .B (n_57_71), .C1 (n_58_72), .C2 (n_61_68) );
AOI211_X1 g_48_74 (.ZN (n_48_74), .A (n_52_72), .B (n_58_69), .C1 (n_56_73), .C2 (n_62_70) );
AOI211_X1 g_46_75 (.ZN (n_46_75), .A (n_50_73), .B (n_56_70), .C1 (n_57_71), .C2 (n_60_71) );
AOI211_X1 g_44_76 (.ZN (n_44_76), .A (n_48_74), .B (n_54_71), .C1 (n_58_69), .C2 (n_58_72) );
AOI211_X1 g_42_77 (.ZN (n_42_77), .A (n_46_75), .B (n_52_72), .C1 (n_56_70), .C2 (n_56_73) );
AOI211_X1 g_40_78 (.ZN (n_40_78), .A (n_44_76), .B (n_50_73), .C1 (n_54_71), .C2 (n_57_71) );
AOI211_X1 g_38_79 (.ZN (n_38_79), .A (n_42_77), .B (n_48_74), .C1 (n_52_72), .C2 (n_58_69) );
AOI211_X1 g_36_80 (.ZN (n_36_80), .A (n_40_78), .B (n_46_75), .C1 (n_50_73), .C2 (n_56_70) );
AOI211_X1 g_34_81 (.ZN (n_34_81), .A (n_38_79), .B (n_44_76), .C1 (n_48_74), .C2 (n_54_71) );
AOI211_X1 g_32_82 (.ZN (n_32_82), .A (n_36_80), .B (n_42_77), .C1 (n_46_75), .C2 (n_52_72) );
AOI211_X1 g_30_83 (.ZN (n_30_83), .A (n_34_81), .B (n_40_78), .C1 (n_44_76), .C2 (n_50_73) );
AOI211_X1 g_28_84 (.ZN (n_28_84), .A (n_32_82), .B (n_38_79), .C1 (n_42_77), .C2 (n_48_74) );
AOI211_X1 g_26_83 (.ZN (n_26_83), .A (n_30_83), .B (n_36_80), .C1 (n_40_78), .C2 (n_46_75) );
AOI211_X1 g_24_84 (.ZN (n_24_84), .A (n_28_84), .B (n_34_81), .C1 (n_38_79), .C2 (n_44_76) );
AOI211_X1 g_22_85 (.ZN (n_22_85), .A (n_26_83), .B (n_32_82), .C1 (n_36_80), .C2 (n_42_77) );
AOI211_X1 g_24_86 (.ZN (n_24_86), .A (n_24_84), .B (n_30_83), .C1 (n_34_81), .C2 (n_40_78) );
AOI211_X1 g_26_85 (.ZN (n_26_85), .A (n_22_85), .B (n_28_84), .C1 (n_32_82), .C2 (n_38_79) );
AOI211_X1 g_25_87 (.ZN (n_25_87), .A (n_24_86), .B (n_26_83), .C1 (n_30_83), .C2 (n_36_80) );
AOI211_X1 g_23_86 (.ZN (n_23_86), .A (n_26_85), .B (n_24_84), .C1 (n_28_84), .C2 (n_34_81) );
AOI211_X1 g_25_85 (.ZN (n_25_85), .A (n_25_87), .B (n_22_85), .C1 (n_26_83), .C2 (n_32_82) );
AOI211_X1 g_27_84 (.ZN (n_27_84), .A (n_23_86), .B (n_24_86), .C1 (n_24_84), .C2 (n_30_83) );
AOI211_X1 g_29_83 (.ZN (n_29_83), .A (n_25_85), .B (n_26_85), .C1 (n_22_85), .C2 (n_28_84) );
AOI211_X1 g_31_82 (.ZN (n_31_82), .A (n_27_84), .B (n_25_87), .C1 (n_24_86), .C2 (n_26_83) );
AOI211_X1 g_33_81 (.ZN (n_33_81), .A (n_29_83), .B (n_23_86), .C1 (n_26_85), .C2 (n_24_84) );
AOI211_X1 g_35_80 (.ZN (n_35_80), .A (n_31_82), .B (n_25_85), .C1 (n_25_87), .C2 (n_22_85) );
AOI211_X1 g_37_79 (.ZN (n_37_79), .A (n_33_81), .B (n_27_84), .C1 (n_23_86), .C2 (n_24_86) );
AOI211_X1 g_39_78 (.ZN (n_39_78), .A (n_35_80), .B (n_29_83), .C1 (n_25_85), .C2 (n_26_85) );
AOI211_X1 g_41_77 (.ZN (n_41_77), .A (n_37_79), .B (n_31_82), .C1 (n_27_84), .C2 (n_25_87) );
AOI211_X1 g_43_76 (.ZN (n_43_76), .A (n_39_78), .B (n_33_81), .C1 (n_29_83), .C2 (n_23_86) );
AOI211_X1 g_45_75 (.ZN (n_45_75), .A (n_41_77), .B (n_35_80), .C1 (n_31_82), .C2 (n_25_85) );
AOI211_X1 g_44_77 (.ZN (n_44_77), .A (n_43_76), .B (n_37_79), .C1 (n_33_81), .C2 (n_27_84) );
AOI211_X1 g_46_76 (.ZN (n_46_76), .A (n_45_75), .B (n_39_78), .C1 (n_35_80), .C2 (n_29_83) );
AOI211_X1 g_45_78 (.ZN (n_45_78), .A (n_44_77), .B (n_41_77), .C1 (n_37_79), .C2 (n_31_82) );
AOI211_X1 g_47_77 (.ZN (n_47_77), .A (n_46_76), .B (n_43_76), .C1 (n_39_78), .C2 (n_33_81) );
AOI211_X1 g_49_76 (.ZN (n_49_76), .A (n_45_78), .B (n_45_75), .C1 (n_41_77), .C2 (n_35_80) );
AOI211_X1 g_51_75 (.ZN (n_51_75), .A (n_47_77), .B (n_44_77), .C1 (n_43_76), .C2 (n_37_79) );
AOI211_X1 g_53_74 (.ZN (n_53_74), .A (n_49_76), .B (n_46_76), .C1 (n_45_75), .C2 (n_39_78) );
AOI211_X1 g_55_73 (.ZN (n_55_73), .A (n_51_75), .B (n_45_78), .C1 (n_44_77), .C2 (n_41_77) );
AOI211_X1 g_57_72 (.ZN (n_57_72), .A (n_53_74), .B (n_47_77), .C1 (n_46_76), .C2 (n_43_76) );
AOI211_X1 g_59_71 (.ZN (n_59_71), .A (n_55_73), .B (n_49_76), .C1 (n_45_78), .C2 (n_45_75) );
AOI211_X1 g_61_70 (.ZN (n_61_70), .A (n_57_72), .B (n_51_75), .C1 (n_47_77), .C2 (n_44_77) );
AOI211_X1 g_63_69 (.ZN (n_63_69), .A (n_59_71), .B (n_53_74), .C1 (n_49_76), .C2 (n_46_76) );
AOI211_X1 g_64_71 (.ZN (n_64_71), .A (n_61_70), .B (n_55_73), .C1 (n_51_75), .C2 (n_45_78) );
AOI211_X1 g_62_72 (.ZN (n_62_72), .A (n_63_69), .B (n_57_72), .C1 (n_53_74), .C2 (n_47_77) );
AOI211_X1 g_63_70 (.ZN (n_63_70), .A (n_64_71), .B (n_59_71), .C1 (n_55_73), .C2 (n_49_76) );
AOI211_X1 g_61_71 (.ZN (n_61_71), .A (n_62_72), .B (n_61_70), .C1 (n_57_72), .C2 (n_51_75) );
AOI211_X1 g_62_69 (.ZN (n_62_69), .A (n_63_70), .B (n_63_69), .C1 (n_59_71), .C2 (n_53_74) );
AOI211_X1 g_60_70 (.ZN (n_60_70), .A (n_61_71), .B (n_64_71), .C1 (n_61_70), .C2 (n_55_73) );
AOI211_X1 g_58_71 (.ZN (n_58_71), .A (n_62_69), .B (n_62_72), .C1 (n_63_69), .C2 (n_57_72) );
AOI211_X1 g_56_72 (.ZN (n_56_72), .A (n_60_70), .B (n_63_70), .C1 (n_64_71), .C2 (n_59_71) );
AOI211_X1 g_54_73 (.ZN (n_54_73), .A (n_58_71), .B (n_61_71), .C1 (n_62_72), .C2 (n_61_70) );
AOI211_X1 g_52_74 (.ZN (n_52_74), .A (n_56_72), .B (n_62_69), .C1 (n_63_70), .C2 (n_63_69) );
AOI211_X1 g_50_75 (.ZN (n_50_75), .A (n_54_73), .B (n_60_70), .C1 (n_61_71), .C2 (n_64_71) );
AOI211_X1 g_48_76 (.ZN (n_48_76), .A (n_52_74), .B (n_58_71), .C1 (n_62_69), .C2 (n_62_72) );
AOI211_X1 g_46_77 (.ZN (n_46_77), .A (n_50_75), .B (n_56_72), .C1 (n_60_70), .C2 (n_63_70) );
AOI211_X1 g_44_78 (.ZN (n_44_78), .A (n_48_76), .B (n_54_73), .C1 (n_58_71), .C2 (n_61_71) );
AOI211_X1 g_42_79 (.ZN (n_42_79), .A (n_46_77), .B (n_52_74), .C1 (n_56_72), .C2 (n_62_69) );
AOI211_X1 g_40_80 (.ZN (n_40_80), .A (n_44_78), .B (n_50_75), .C1 (n_54_73), .C2 (n_60_70) );
AOI211_X1 g_38_81 (.ZN (n_38_81), .A (n_42_79), .B (n_48_76), .C1 (n_52_74), .C2 (n_58_71) );
AOI211_X1 g_36_82 (.ZN (n_36_82), .A (n_40_80), .B (n_46_77), .C1 (n_50_75), .C2 (n_56_72) );
AOI211_X1 g_34_83 (.ZN (n_34_83), .A (n_38_81), .B (n_44_78), .C1 (n_48_76), .C2 (n_54_73) );
AOI211_X1 g_35_81 (.ZN (n_35_81), .A (n_36_82), .B (n_42_79), .C1 (n_46_77), .C2 (n_52_74) );
AOI211_X1 g_33_82 (.ZN (n_33_82), .A (n_34_83), .B (n_40_80), .C1 (n_44_78), .C2 (n_50_75) );
AOI211_X1 g_31_83 (.ZN (n_31_83), .A (n_35_81), .B (n_38_81), .C1 (n_42_79), .C2 (n_48_76) );
AOI211_X1 g_29_84 (.ZN (n_29_84), .A (n_33_82), .B (n_36_82), .C1 (n_40_80), .C2 (n_46_77) );
AOI211_X1 g_27_85 (.ZN (n_27_85), .A (n_31_83), .B (n_34_83), .C1 (n_38_81), .C2 (n_44_78) );
AOI211_X1 g_25_86 (.ZN (n_25_86), .A (n_29_84), .B (n_35_81), .C1 (n_36_82), .C2 (n_42_79) );
AOI211_X1 g_23_87 (.ZN (n_23_87), .A (n_27_85), .B (n_33_82), .C1 (n_34_83), .C2 (n_40_80) );
AOI211_X1 g_21_88 (.ZN (n_21_88), .A (n_25_86), .B (n_31_83), .C1 (n_35_81), .C2 (n_38_81) );
AOI211_X1 g_19_89 (.ZN (n_19_89), .A (n_23_87), .B (n_29_84), .C1 (n_33_82), .C2 (n_36_82) );
AOI211_X1 g_17_90 (.ZN (n_17_90), .A (n_21_88), .B (n_27_85), .C1 (n_31_83), .C2 (n_34_83) );
AOI211_X1 g_15_91 (.ZN (n_15_91), .A (n_19_89), .B (n_25_86), .C1 (n_29_84), .C2 (n_35_81) );
AOI211_X1 g_13_92 (.ZN (n_13_92), .A (n_17_90), .B (n_23_87), .C1 (n_27_85), .C2 (n_33_82) );
AOI211_X1 g_11_93 (.ZN (n_11_93), .A (n_15_91), .B (n_21_88), .C1 (n_25_86), .C2 (n_31_83) );
AOI211_X1 g_10_95 (.ZN (n_10_95), .A (n_13_92), .B (n_19_89), .C1 (n_23_87), .C2 (n_29_84) );
AOI211_X1 g_9_93 (.ZN (n_9_93), .A (n_11_93), .B (n_17_90), .C1 (n_21_88), .C2 (n_27_85) );
AOI211_X1 g_8_95 (.ZN (n_8_95), .A (n_10_95), .B (n_15_91), .C1 (n_19_89), .C2 (n_25_86) );
AOI211_X1 g_9_97 (.ZN (n_9_97), .A (n_9_93), .B (n_13_92), .C1 (n_17_90), .C2 (n_23_87) );
AOI211_X1 g_10_99 (.ZN (n_10_99), .A (n_8_95), .B (n_11_93), .C1 (n_15_91), .C2 (n_21_88) );
AOI211_X1 g_11_97 (.ZN (n_11_97), .A (n_9_97), .B (n_10_95), .C1 (n_13_92), .C2 (n_19_89) );
AOI211_X1 g_13_96 (.ZN (n_13_96), .A (n_10_99), .B (n_9_93), .C1 (n_11_93), .C2 (n_17_90) );
AOI211_X1 g_12_98 (.ZN (n_12_98), .A (n_11_97), .B (n_8_95), .C1 (n_10_95), .C2 (n_15_91) );
AOI211_X1 g_11_96 (.ZN (n_11_96), .A (n_13_96), .B (n_9_97), .C1 (n_9_93), .C2 (n_13_92) );
AOI211_X1 g_12_94 (.ZN (n_12_94), .A (n_12_98), .B (n_10_99), .C1 (n_8_95), .C2 (n_11_93) );
AOI211_X1 g_11_92 (.ZN (n_11_92), .A (n_11_96), .B (n_11_97), .C1 (n_9_97), .C2 (n_10_95) );
AOI211_X1 g_10_94 (.ZN (n_10_94), .A (n_12_94), .B (n_13_96), .C1 (n_10_99), .C2 (n_9_93) );
AOI211_X1 g_12_93 (.ZN (n_12_93), .A (n_11_92), .B (n_12_98), .C1 (n_11_97), .C2 (n_8_95) );
AOI211_X1 g_13_91 (.ZN (n_13_91), .A (n_10_94), .B (n_11_96), .C1 (n_13_96), .C2 (n_9_97) );
AOI211_X1 g_15_90 (.ZN (n_15_90), .A (n_12_93), .B (n_12_94), .C1 (n_12_98), .C2 (n_10_99) );
AOI211_X1 g_17_89 (.ZN (n_17_89), .A (n_13_91), .B (n_11_92), .C1 (n_11_96), .C2 (n_11_97) );
AOI211_X1 g_19_88 (.ZN (n_19_88), .A (n_15_90), .B (n_10_94), .C1 (n_12_94), .C2 (n_13_96) );
AOI211_X1 g_21_87 (.ZN (n_21_87), .A (n_17_89), .B (n_12_93), .C1 (n_11_92), .C2 (n_12_98) );
AOI211_X1 g_23_88 (.ZN (n_23_88), .A (n_19_88), .B (n_13_91), .C1 (n_10_94), .C2 (n_11_96) );
AOI211_X1 g_21_89 (.ZN (n_21_89), .A (n_21_87), .B (n_15_90), .C1 (n_12_93), .C2 (n_12_94) );
AOI211_X1 g_19_90 (.ZN (n_19_90), .A (n_23_88), .B (n_17_89), .C1 (n_13_91), .C2 (n_11_92) );
AOI211_X1 g_17_91 (.ZN (n_17_91), .A (n_21_89), .B (n_19_88), .C1 (n_15_90), .C2 (n_10_94) );
AOI211_X1 g_15_92 (.ZN (n_15_92), .A (n_19_90), .B (n_21_87), .C1 (n_17_89), .C2 (n_12_93) );
AOI211_X1 g_13_93 (.ZN (n_13_93), .A (n_17_91), .B (n_23_88), .C1 (n_19_88), .C2 (n_13_91) );
AOI211_X1 g_11_94 (.ZN (n_11_94), .A (n_15_92), .B (n_21_89), .C1 (n_21_87), .C2 (n_15_90) );
AOI211_X1 g_10_96 (.ZN (n_10_96), .A (n_13_93), .B (n_19_90), .C1 (n_23_88), .C2 (n_17_89) );
AOI211_X1 g_12_95 (.ZN (n_12_95), .A (n_11_94), .B (n_17_91), .C1 (n_21_89), .C2 (n_19_88) );
AOI211_X1 g_14_94 (.ZN (n_14_94), .A (n_10_96), .B (n_15_92), .C1 (n_19_90), .C2 (n_21_87) );
AOI211_X1 g_16_93 (.ZN (n_16_93), .A (n_12_95), .B (n_13_93), .C1 (n_17_91), .C2 (n_23_88) );
AOI211_X1 g_14_92 (.ZN (n_14_92), .A (n_14_94), .B (n_11_94), .C1 (n_15_92), .C2 (n_21_89) );
AOI211_X1 g_16_91 (.ZN (n_16_91), .A (n_16_93), .B (n_10_96), .C1 (n_13_93), .C2 (n_19_90) );
AOI211_X1 g_18_90 (.ZN (n_18_90), .A (n_14_92), .B (n_12_95), .C1 (n_11_94), .C2 (n_17_91) );
AOI211_X1 g_20_89 (.ZN (n_20_89), .A (n_16_91), .B (n_14_94), .C1 (n_10_96), .C2 (n_15_92) );
AOI211_X1 g_22_88 (.ZN (n_22_88), .A (n_18_90), .B (n_16_93), .C1 (n_12_95), .C2 (n_13_93) );
AOI211_X1 g_24_87 (.ZN (n_24_87), .A (n_20_89), .B (n_14_92), .C1 (n_14_94), .C2 (n_11_94) );
AOI211_X1 g_26_86 (.ZN (n_26_86), .A (n_22_88), .B (n_16_91), .C1 (n_16_93), .C2 (n_10_96) );
AOI211_X1 g_28_85 (.ZN (n_28_85), .A (n_24_87), .B (n_18_90), .C1 (n_14_92), .C2 (n_12_95) );
AOI211_X1 g_30_84 (.ZN (n_30_84), .A (n_26_86), .B (n_20_89), .C1 (n_16_91), .C2 (n_14_94) );
AOI211_X1 g_32_83 (.ZN (n_32_83), .A (n_28_85), .B (n_22_88), .C1 (n_18_90), .C2 (n_16_93) );
AOI211_X1 g_34_82 (.ZN (n_34_82), .A (n_30_84), .B (n_24_87), .C1 (n_20_89), .C2 (n_14_92) );
AOI211_X1 g_36_81 (.ZN (n_36_81), .A (n_32_83), .B (n_26_86), .C1 (n_22_88), .C2 (n_16_91) );
AOI211_X1 g_38_80 (.ZN (n_38_80), .A (n_34_82), .B (n_28_85), .C1 (n_24_87), .C2 (n_18_90) );
AOI211_X1 g_40_79 (.ZN (n_40_79), .A (n_36_81), .B (n_30_84), .C1 (n_26_86), .C2 (n_20_89) );
AOI211_X1 g_42_78 (.ZN (n_42_78), .A (n_38_80), .B (n_32_83), .C1 (n_28_85), .C2 (n_22_88) );
AOI211_X1 g_41_80 (.ZN (n_41_80), .A (n_40_79), .B (n_34_82), .C1 (n_30_84), .C2 (n_24_87) );
AOI211_X1 g_43_79 (.ZN (n_43_79), .A (n_42_78), .B (n_36_81), .C1 (n_32_83), .C2 (n_26_86) );
AOI211_X1 g_42_81 (.ZN (n_42_81), .A (n_41_80), .B (n_38_80), .C1 (n_34_82), .C2 (n_28_85) );
AOI211_X1 g_41_79 (.ZN (n_41_79), .A (n_43_79), .B (n_40_79), .C1 (n_36_81), .C2 (n_30_84) );
AOI211_X1 g_43_78 (.ZN (n_43_78), .A (n_42_81), .B (n_42_78), .C1 (n_38_80), .C2 (n_32_83) );
AOI211_X1 g_45_77 (.ZN (n_45_77), .A (n_41_79), .B (n_41_80), .C1 (n_40_79), .C2 (n_34_82) );
AOI211_X1 g_47_76 (.ZN (n_47_76), .A (n_43_78), .B (n_43_79), .C1 (n_42_78), .C2 (n_36_81) );
AOI211_X1 g_49_75 (.ZN (n_49_75), .A (n_45_77), .B (n_42_81), .C1 (n_41_80), .C2 (n_38_80) );
AOI211_X1 g_51_74 (.ZN (n_51_74), .A (n_47_76), .B (n_41_79), .C1 (n_43_79), .C2 (n_40_79) );
AOI211_X1 g_53_73 (.ZN (n_53_73), .A (n_49_75), .B (n_43_78), .C1 (n_42_81), .C2 (n_42_78) );
AOI211_X1 g_55_72 (.ZN (n_55_72), .A (n_51_74), .B (n_45_77), .C1 (n_41_79), .C2 (n_41_80) );
AOI211_X1 g_54_74 (.ZN (n_54_74), .A (n_53_73), .B (n_47_76), .C1 (n_43_78), .C2 (n_43_79) );
AOI211_X1 g_52_75 (.ZN (n_52_75), .A (n_55_72), .B (n_49_75), .C1 (n_45_77), .C2 (n_42_81) );
AOI211_X1 g_50_76 (.ZN (n_50_76), .A (n_54_74), .B (n_51_74), .C1 (n_47_76), .C2 (n_41_79) );
AOI211_X1 g_48_77 (.ZN (n_48_77), .A (n_52_75), .B (n_53_73), .C1 (n_49_75), .C2 (n_43_78) );
AOI211_X1 g_46_78 (.ZN (n_46_78), .A (n_50_76), .B (n_55_72), .C1 (n_51_74), .C2 (n_45_77) );
AOI211_X1 g_44_79 (.ZN (n_44_79), .A (n_48_77), .B (n_54_74), .C1 (n_53_73), .C2 (n_47_76) );
AOI211_X1 g_42_80 (.ZN (n_42_80), .A (n_46_78), .B (n_52_75), .C1 (n_55_72), .C2 (n_49_75) );
AOI211_X1 g_40_81 (.ZN (n_40_81), .A (n_44_79), .B (n_50_76), .C1 (n_54_74), .C2 (n_51_74) );
AOI211_X1 g_38_82 (.ZN (n_38_82), .A (n_42_80), .B (n_48_77), .C1 (n_52_75), .C2 (n_53_73) );
AOI211_X1 g_39_80 (.ZN (n_39_80), .A (n_40_81), .B (n_46_78), .C1 (n_50_76), .C2 (n_55_72) );
AOI211_X1 g_37_81 (.ZN (n_37_81), .A (n_38_82), .B (n_44_79), .C1 (n_48_77), .C2 (n_54_74) );
AOI211_X1 g_35_82 (.ZN (n_35_82), .A (n_39_80), .B (n_42_80), .C1 (n_46_78), .C2 (n_52_75) );
AOI211_X1 g_33_83 (.ZN (n_33_83), .A (n_37_81), .B (n_40_81), .C1 (n_44_79), .C2 (n_50_76) );
AOI211_X1 g_31_84 (.ZN (n_31_84), .A (n_35_82), .B (n_38_82), .C1 (n_42_80), .C2 (n_48_77) );
AOI211_X1 g_29_85 (.ZN (n_29_85), .A (n_33_83), .B (n_39_80), .C1 (n_40_81), .C2 (n_46_78) );
AOI211_X1 g_27_86 (.ZN (n_27_86), .A (n_31_84), .B (n_37_81), .C1 (n_38_82), .C2 (n_44_79) );
AOI211_X1 g_26_88 (.ZN (n_26_88), .A (n_29_85), .B (n_35_82), .C1 (n_39_80), .C2 (n_42_80) );
AOI211_X1 g_28_87 (.ZN (n_28_87), .A (n_27_86), .B (n_33_83), .C1 (n_37_81), .C2 (n_40_81) );
AOI211_X1 g_30_86 (.ZN (n_30_86), .A (n_26_88), .B (n_31_84), .C1 (n_35_82), .C2 (n_38_82) );
AOI211_X1 g_32_85 (.ZN (n_32_85), .A (n_28_87), .B (n_29_85), .C1 (n_33_83), .C2 (n_39_80) );
AOI211_X1 g_34_84 (.ZN (n_34_84), .A (n_30_86), .B (n_27_86), .C1 (n_31_84), .C2 (n_37_81) );
AOI211_X1 g_36_83 (.ZN (n_36_83), .A (n_32_85), .B (n_26_88), .C1 (n_29_85), .C2 (n_35_82) );
AOI211_X1 g_35_85 (.ZN (n_35_85), .A (n_34_84), .B (n_28_87), .C1 (n_27_86), .C2 (n_33_83) );
AOI211_X1 g_33_84 (.ZN (n_33_84), .A (n_36_83), .B (n_30_86), .C1 (n_26_88), .C2 (n_31_84) );
AOI211_X1 g_35_83 (.ZN (n_35_83), .A (n_35_85), .B (n_32_85), .C1 (n_28_87), .C2 (n_29_85) );
AOI211_X1 g_37_82 (.ZN (n_37_82), .A (n_33_84), .B (n_34_84), .C1 (n_30_86), .C2 (n_27_86) );
AOI211_X1 g_39_81 (.ZN (n_39_81), .A (n_35_83), .B (n_36_83), .C1 (n_32_85), .C2 (n_26_88) );
AOI211_X1 g_38_83 (.ZN (n_38_83), .A (n_37_82), .B (n_35_85), .C1 (n_34_84), .C2 (n_28_87) );
AOI211_X1 g_40_82 (.ZN (n_40_82), .A (n_39_81), .B (n_33_84), .C1 (n_36_83), .C2 (n_30_86) );
AOI211_X1 g_39_84 (.ZN (n_39_84), .A (n_38_83), .B (n_35_83), .C1 (n_35_85), .C2 (n_32_85) );
AOI211_X1 g_37_83 (.ZN (n_37_83), .A (n_40_82), .B (n_37_82), .C1 (n_33_84), .C2 (n_34_84) );
AOI211_X1 g_39_82 (.ZN (n_39_82), .A (n_39_84), .B (n_39_81), .C1 (n_35_83), .C2 (n_36_83) );
AOI211_X1 g_41_81 (.ZN (n_41_81), .A (n_37_83), .B (n_38_83), .C1 (n_37_82), .C2 (n_35_85) );
AOI211_X1 g_43_80 (.ZN (n_43_80), .A (n_39_82), .B (n_40_82), .C1 (n_39_81), .C2 (n_33_84) );
AOI211_X1 g_45_79 (.ZN (n_45_79), .A (n_41_81), .B (n_39_84), .C1 (n_38_83), .C2 (n_35_83) );
AOI211_X1 g_47_78 (.ZN (n_47_78), .A (n_43_80), .B (n_37_83), .C1 (n_40_82), .C2 (n_37_82) );
AOI211_X1 g_49_77 (.ZN (n_49_77), .A (n_45_79), .B (n_39_82), .C1 (n_39_84), .C2 (n_39_81) );
AOI211_X1 g_51_76 (.ZN (n_51_76), .A (n_47_78), .B (n_41_81), .C1 (n_37_83), .C2 (n_38_83) );
AOI211_X1 g_53_75 (.ZN (n_53_75), .A (n_49_77), .B (n_43_80), .C1 (n_39_82), .C2 (n_40_82) );
AOI211_X1 g_55_74 (.ZN (n_55_74), .A (n_51_76), .B (n_45_79), .C1 (n_41_81), .C2 (n_39_84) );
AOI211_X1 g_57_73 (.ZN (n_57_73), .A (n_53_75), .B (n_47_78), .C1 (n_43_80), .C2 (n_37_83) );
AOI211_X1 g_59_72 (.ZN (n_59_72), .A (n_55_74), .B (n_49_77), .C1 (n_45_79), .C2 (n_39_82) );
AOI211_X1 g_58_74 (.ZN (n_58_74), .A (n_57_73), .B (n_51_76), .C1 (n_47_78), .C2 (n_41_81) );
AOI211_X1 g_60_73 (.ZN (n_60_73), .A (n_59_72), .B (n_53_75), .C1 (n_49_77), .C2 (n_43_80) );
AOI211_X1 g_59_75 (.ZN (n_59_75), .A (n_58_74), .B (n_55_74), .C1 (n_51_76), .C2 (n_45_79) );
AOI211_X1 g_58_73 (.ZN (n_58_73), .A (n_60_73), .B (n_57_73), .C1 (n_53_75), .C2 (n_47_78) );
AOI211_X1 g_60_72 (.ZN (n_60_72), .A (n_59_75), .B (n_59_72), .C1 (n_55_74), .C2 (n_49_77) );
AOI211_X1 g_62_71 (.ZN (n_62_71), .A (n_58_73), .B (n_58_74), .C1 (n_57_73), .C2 (n_51_76) );
AOI211_X1 g_64_70 (.ZN (n_64_70), .A (n_60_72), .B (n_60_73), .C1 (n_59_72), .C2 (n_53_75) );
AOI211_X1 g_66_69 (.ZN (n_66_69), .A (n_62_71), .B (n_59_75), .C1 (n_58_74), .C2 (n_55_74) );
AOI211_X1 g_68_68 (.ZN (n_68_68), .A (n_64_70), .B (n_58_73), .C1 (n_60_73), .C2 (n_57_73) );
AOI211_X1 g_70_67 (.ZN (n_70_67), .A (n_66_69), .B (n_60_72), .C1 (n_59_75), .C2 (n_59_72) );
AOI211_X1 g_69_69 (.ZN (n_69_69), .A (n_68_68), .B (n_62_71), .C1 (n_58_73), .C2 (n_58_74) );
AOI211_X1 g_71_68 (.ZN (n_71_68), .A (n_70_67), .B (n_64_70), .C1 (n_60_72), .C2 (n_60_73) );
AOI211_X1 g_73_67 (.ZN (n_73_67), .A (n_69_69), .B (n_66_69), .C1 (n_62_71), .C2 (n_59_75) );
AOI211_X1 g_71_66 (.ZN (n_71_66), .A (n_71_68), .B (n_68_68), .C1 (n_64_70), .C2 (n_58_73) );
AOI211_X1 g_73_65 (.ZN (n_73_65), .A (n_73_67), .B (n_70_67), .C1 (n_66_69), .C2 (n_60_72) );
AOI211_X1 g_75_64 (.ZN (n_75_64), .A (n_71_66), .B (n_69_69), .C1 (n_68_68), .C2 (n_62_71) );
AOI211_X1 g_77_63 (.ZN (n_77_63), .A (n_73_65), .B (n_71_68), .C1 (n_70_67), .C2 (n_64_70) );
AOI211_X1 g_79_64 (.ZN (n_79_64), .A (n_75_64), .B (n_73_67), .C1 (n_69_69), .C2 (n_66_69) );
AOI211_X1 g_77_65 (.ZN (n_77_65), .A (n_77_63), .B (n_71_66), .C1 (n_71_68), .C2 (n_68_68) );
AOI211_X1 g_75_66 (.ZN (n_75_66), .A (n_79_64), .B (n_73_65), .C1 (n_73_67), .C2 (n_70_67) );
AOI211_X1 g_74_68 (.ZN (n_74_68), .A (n_77_65), .B (n_75_64), .C1 (n_71_66), .C2 (n_69_69) );
AOI211_X1 g_73_66 (.ZN (n_73_66), .A (n_75_66), .B (n_77_63), .C1 (n_73_65), .C2 (n_71_68) );
AOI211_X1 g_75_65 (.ZN (n_75_65), .A (n_74_68), .B (n_79_64), .C1 (n_75_64), .C2 (n_73_67) );
AOI211_X1 g_77_64 (.ZN (n_77_64), .A (n_73_66), .B (n_77_65), .C1 (n_77_63), .C2 (n_71_66) );
AOI211_X1 g_79_63 (.ZN (n_79_63), .A (n_75_65), .B (n_75_66), .C1 (n_79_64), .C2 (n_73_65) );
AOI211_X1 g_81_62 (.ZN (n_81_62), .A (n_77_64), .B (n_74_68), .C1 (n_77_65), .C2 (n_75_64) );
AOI211_X1 g_80_64 (.ZN (n_80_64), .A (n_79_63), .B (n_73_66), .C1 (n_75_66), .C2 (n_77_63) );
AOI211_X1 g_82_63 (.ZN (n_82_63), .A (n_81_62), .B (n_75_65), .C1 (n_74_68), .C2 (n_79_64) );
AOI211_X1 g_84_62 (.ZN (n_84_62), .A (n_80_64), .B (n_77_64), .C1 (n_73_66), .C2 (n_77_65) );
AOI211_X1 g_86_61 (.ZN (n_86_61), .A (n_82_63), .B (n_79_63), .C1 (n_75_65), .C2 (n_75_66) );
AOI211_X1 g_88_60 (.ZN (n_88_60), .A (n_84_62), .B (n_81_62), .C1 (n_77_64), .C2 (n_74_68) );
AOI211_X1 g_90_59 (.ZN (n_90_59), .A (n_86_61), .B (n_80_64), .C1 (n_79_63), .C2 (n_73_66) );
AOI211_X1 g_92_58 (.ZN (n_92_58), .A (n_88_60), .B (n_82_63), .C1 (n_81_62), .C2 (n_75_65) );
AOI211_X1 g_94_59 (.ZN (n_94_59), .A (n_90_59), .B (n_84_62), .C1 (n_80_64), .C2 (n_77_64) );
AOI211_X1 g_92_60 (.ZN (n_92_60), .A (n_92_58), .B (n_86_61), .C1 (n_82_63), .C2 (n_79_63) );
AOI211_X1 g_94_61 (.ZN (n_94_61), .A (n_94_59), .B (n_88_60), .C1 (n_84_62), .C2 (n_81_62) );
AOI211_X1 g_95_63 (.ZN (n_95_63), .A (n_92_60), .B (n_90_59), .C1 (n_86_61), .C2 (n_80_64) );
AOI211_X1 g_96_65 (.ZN (n_96_65), .A (n_94_61), .B (n_92_58), .C1 (n_88_60), .C2 (n_82_63) );
AOI211_X1 g_97_67 (.ZN (n_97_67), .A (n_95_63), .B (n_94_59), .C1 (n_90_59), .C2 (n_84_62) );
AOI211_X1 g_98_69 (.ZN (n_98_69), .A (n_96_65), .B (n_92_60), .C1 (n_92_58), .C2 (n_86_61) );
AOI211_X1 g_99_71 (.ZN (n_99_71), .A (n_97_67), .B (n_94_61), .C1 (n_94_59), .C2 (n_88_60) );
AOI211_X1 g_100_73 (.ZN (n_100_73), .A (n_98_69), .B (n_95_63), .C1 (n_92_60), .C2 (n_90_59) );
AOI211_X1 g_98_72 (.ZN (n_98_72), .A (n_99_71), .B (n_96_65), .C1 (n_94_61), .C2 (n_92_58) );
AOI211_X1 g_97_70 (.ZN (n_97_70), .A (n_100_73), .B (n_97_67), .C1 (n_95_63), .C2 (n_94_59) );
AOI211_X1 g_96_68 (.ZN (n_96_68), .A (n_98_72), .B (n_98_69), .C1 (n_96_65), .C2 (n_92_60) );
AOI211_X1 g_95_66 (.ZN (n_95_66), .A (n_97_70), .B (n_99_71), .C1 (n_97_67), .C2 (n_94_61) );
AOI211_X1 g_97_65 (.ZN (n_97_65), .A (n_96_68), .B (n_100_73), .C1 (n_98_69), .C2 (n_95_63) );
AOI211_X1 g_96_63 (.ZN (n_96_63), .A (n_95_66), .B (n_98_72), .C1 (n_99_71), .C2 (n_96_65) );
AOI211_X1 g_95_61 (.ZN (n_95_61), .A (n_97_65), .B (n_97_70), .C1 (n_100_73), .C2 (n_97_67) );
AOI211_X1 g_93_60 (.ZN (n_93_60), .A (n_96_63), .B (n_96_68), .C1 (n_98_72), .C2 (n_98_69) );
AOI211_X1 g_91_59 (.ZN (n_91_59), .A (n_95_61), .B (n_95_66), .C1 (n_97_70), .C2 (n_99_71) );
AOI211_X1 g_90_61 (.ZN (n_90_61), .A (n_93_60), .B (n_97_65), .C1 (n_96_68), .C2 (n_100_73) );
AOI211_X1 g_88_62 (.ZN (n_88_62), .A (n_91_59), .B (n_96_63), .C1 (n_95_66), .C2 (n_98_72) );
AOI211_X1 g_89_60 (.ZN (n_89_60), .A (n_90_61), .B (n_95_61), .C1 (n_97_65), .C2 (n_97_70) );
AOI211_X1 g_90_58 (.ZN (n_90_58), .A (n_88_62), .B (n_93_60), .C1 (n_96_63), .C2 (n_96_68) );
AOI211_X1 g_88_59 (.ZN (n_88_59), .A (n_89_60), .B (n_91_59), .C1 (n_95_61), .C2 (n_95_66) );
AOI211_X1 g_86_60 (.ZN (n_86_60), .A (n_90_58), .B (n_90_61), .C1 (n_93_60), .C2 (n_97_65) );
AOI211_X1 g_84_61 (.ZN (n_84_61), .A (n_88_59), .B (n_88_62), .C1 (n_91_59), .C2 (n_96_63) );
AOI211_X1 g_82_62 (.ZN (n_82_62), .A (n_86_60), .B (n_89_60), .C1 (n_90_61), .C2 (n_95_61) );
AOI211_X1 g_80_63 (.ZN (n_80_63), .A (n_84_61), .B (n_90_58), .C1 (n_88_62), .C2 (n_93_60) );
AOI211_X1 g_78_64 (.ZN (n_78_64), .A (n_82_62), .B (n_88_59), .C1 (n_89_60), .C2 (n_91_59) );
AOI211_X1 g_76_65 (.ZN (n_76_65), .A (n_80_63), .B (n_86_60), .C1 (n_90_58), .C2 (n_90_61) );
AOI211_X1 g_74_66 (.ZN (n_74_66), .A (n_78_64), .B (n_84_61), .C1 (n_88_59), .C2 (n_88_62) );
AOI211_X1 g_72_67 (.ZN (n_72_67), .A (n_76_65), .B (n_82_62), .C1 (n_86_60), .C2 (n_89_60) );
AOI211_X1 g_70_68 (.ZN (n_70_68), .A (n_74_66), .B (n_80_63), .C1 (n_84_61), .C2 (n_90_58) );
AOI211_X1 g_68_69 (.ZN (n_68_69), .A (n_72_67), .B (n_78_64), .C1 (n_82_62), .C2 (n_88_59) );
AOI211_X1 g_67_71 (.ZN (n_67_71), .A (n_70_68), .B (n_76_65), .C1 (n_80_63), .C2 (n_86_60) );
AOI211_X1 g_65_70 (.ZN (n_65_70), .A (n_68_69), .B (n_74_66), .C1 (n_78_64), .C2 (n_84_61) );
AOI211_X1 g_67_69 (.ZN (n_67_69), .A (n_67_71), .B (n_72_67), .C1 (n_76_65), .C2 (n_82_62) );
AOI211_X1 g_69_68 (.ZN (n_69_68), .A (n_65_70), .B (n_70_68), .C1 (n_74_66), .C2 (n_80_63) );
AOI211_X1 g_71_67 (.ZN (n_71_67), .A (n_67_69), .B (n_68_69), .C1 (n_72_67), .C2 (n_78_64) );
AOI211_X1 g_72_69 (.ZN (n_72_69), .A (n_69_68), .B (n_67_71), .C1 (n_70_68), .C2 (n_76_65) );
AOI211_X1 g_70_70 (.ZN (n_70_70), .A (n_71_67), .B (n_65_70), .C1 (n_68_69), .C2 (n_74_66) );
AOI211_X1 g_68_71 (.ZN (n_68_71), .A (n_72_69), .B (n_67_69), .C1 (n_67_71), .C2 (n_72_67) );
AOI211_X1 g_66_72 (.ZN (n_66_72), .A (n_70_70), .B (n_69_68), .C1 (n_65_70), .C2 (n_70_68) );
AOI211_X1 g_67_70 (.ZN (n_67_70), .A (n_68_71), .B (n_71_67), .C1 (n_67_69), .C2 (n_68_69) );
AOI211_X1 g_65_71 (.ZN (n_65_71), .A (n_66_72), .B (n_72_69), .C1 (n_69_68), .C2 (n_67_71) );
AOI211_X1 g_63_72 (.ZN (n_63_72), .A (n_67_70), .B (n_70_70), .C1 (n_71_67), .C2 (n_65_70) );
AOI211_X1 g_61_73 (.ZN (n_61_73), .A (n_65_71), .B (n_68_71), .C1 (n_72_69), .C2 (n_67_69) );
AOI211_X1 g_59_74 (.ZN (n_59_74), .A (n_63_72), .B (n_66_72), .C1 (n_70_70), .C2 (n_69_68) );
AOI211_X1 g_57_75 (.ZN (n_57_75), .A (n_61_73), .B (n_67_70), .C1 (n_68_71), .C2 (n_71_67) );
AOI211_X1 g_55_76 (.ZN (n_55_76), .A (n_59_74), .B (n_65_71), .C1 (n_66_72), .C2 (n_72_69) );
AOI211_X1 g_56_74 (.ZN (n_56_74), .A (n_57_75), .B (n_63_72), .C1 (n_67_70), .C2 (n_70_70) );
AOI211_X1 g_54_75 (.ZN (n_54_75), .A (n_55_76), .B (n_61_73), .C1 (n_65_71), .C2 (n_68_71) );
AOI211_X1 g_52_76 (.ZN (n_52_76), .A (n_56_74), .B (n_59_74), .C1 (n_63_72), .C2 (n_66_72) );
AOI211_X1 g_50_77 (.ZN (n_50_77), .A (n_54_75), .B (n_57_75), .C1 (n_61_73), .C2 (n_67_70) );
AOI211_X1 g_48_78 (.ZN (n_48_78), .A (n_52_76), .B (n_55_76), .C1 (n_59_74), .C2 (n_65_71) );
AOI211_X1 g_46_79 (.ZN (n_46_79), .A (n_50_77), .B (n_56_74), .C1 (n_57_75), .C2 (n_63_72) );
AOI211_X1 g_44_80 (.ZN (n_44_80), .A (n_48_78), .B (n_54_75), .C1 (n_55_76), .C2 (n_61_73) );
AOI211_X1 g_43_82 (.ZN (n_43_82), .A (n_46_79), .B (n_52_76), .C1 (n_56_74), .C2 (n_59_74) );
AOI211_X1 g_41_83 (.ZN (n_41_83), .A (n_44_80), .B (n_50_77), .C1 (n_54_75), .C2 (n_57_75) );
AOI211_X1 g_40_85 (.ZN (n_40_85), .A (n_43_82), .B (n_48_78), .C1 (n_52_76), .C2 (n_55_76) );
AOI211_X1 g_39_83 (.ZN (n_39_83), .A (n_41_83), .B (n_46_79), .C1 (n_50_77), .C2 (n_56_74) );
AOI211_X1 g_37_84 (.ZN (n_37_84), .A (n_40_85), .B (n_44_80), .C1 (n_48_78), .C2 (n_54_75) );
AOI211_X1 g_38_86 (.ZN (n_38_86), .A (n_39_83), .B (n_43_82), .C1 (n_46_79), .C2 (n_52_76) );
AOI211_X1 g_36_85 (.ZN (n_36_85), .A (n_37_84), .B (n_41_83), .C1 (n_44_80), .C2 (n_50_77) );
AOI211_X1 g_38_84 (.ZN (n_38_84), .A (n_38_86), .B (n_40_85), .C1 (n_43_82), .C2 (n_48_78) );
AOI211_X1 g_40_83 (.ZN (n_40_83), .A (n_36_85), .B (n_39_83), .C1 (n_41_83), .C2 (n_46_79) );
AOI211_X1 g_42_82 (.ZN (n_42_82), .A (n_38_84), .B (n_37_84), .C1 (n_40_85), .C2 (n_44_80) );
AOI211_X1 g_44_81 (.ZN (n_44_81), .A (n_40_83), .B (n_38_86), .C1 (n_39_83), .C2 (n_43_82) );
AOI211_X1 g_46_80 (.ZN (n_46_80), .A (n_42_82), .B (n_36_85), .C1 (n_37_84), .C2 (n_41_83) );
AOI211_X1 g_48_79 (.ZN (n_48_79), .A (n_44_81), .B (n_38_84), .C1 (n_38_86), .C2 (n_40_85) );
AOI211_X1 g_50_78 (.ZN (n_50_78), .A (n_46_80), .B (n_40_83), .C1 (n_36_85), .C2 (n_39_83) );
AOI211_X1 g_52_77 (.ZN (n_52_77), .A (n_48_79), .B (n_42_82), .C1 (n_38_84), .C2 (n_37_84) );
AOI211_X1 g_54_76 (.ZN (n_54_76), .A (n_50_78), .B (n_44_81), .C1 (n_40_83), .C2 (n_38_86) );
AOI211_X1 g_56_75 (.ZN (n_56_75), .A (n_52_77), .B (n_46_80), .C1 (n_42_82), .C2 (n_36_85) );
AOI211_X1 g_55_77 (.ZN (n_55_77), .A (n_54_76), .B (n_48_79), .C1 (n_44_81), .C2 (n_38_84) );
AOI211_X1 g_57_76 (.ZN (n_57_76), .A (n_56_75), .B (n_50_78), .C1 (n_46_80), .C2 (n_40_83) );
AOI211_X1 g_55_75 (.ZN (n_55_75), .A (n_55_77), .B (n_52_77), .C1 (n_48_79), .C2 (n_42_82) );
AOI211_X1 g_57_74 (.ZN (n_57_74), .A (n_57_76), .B (n_54_76), .C1 (n_50_78), .C2 (n_44_81) );
AOI211_X1 g_59_73 (.ZN (n_59_73), .A (n_55_75), .B (n_56_75), .C1 (n_52_77), .C2 (n_46_80) );
AOI211_X1 g_61_72 (.ZN (n_61_72), .A (n_57_74), .B (n_55_77), .C1 (n_54_76), .C2 (n_48_79) );
AOI211_X1 g_63_71 (.ZN (n_63_71), .A (n_59_73), .B (n_57_76), .C1 (n_56_75), .C2 (n_50_78) );
AOI211_X1 g_64_73 (.ZN (n_64_73), .A (n_61_72), .B (n_55_75), .C1 (n_55_77), .C2 (n_52_77) );
AOI211_X1 g_62_74 (.ZN (n_62_74), .A (n_63_71), .B (n_57_74), .C1 (n_57_76), .C2 (n_54_76) );
AOI211_X1 g_60_75 (.ZN (n_60_75), .A (n_64_73), .B (n_59_73), .C1 (n_55_75), .C2 (n_56_75) );
AOI211_X1 g_58_76 (.ZN (n_58_76), .A (n_62_74), .B (n_61_72), .C1 (n_57_74), .C2 (n_55_77) );
AOI211_X1 g_56_77 (.ZN (n_56_77), .A (n_60_75), .B (n_63_71), .C1 (n_59_73), .C2 (n_57_76) );
AOI211_X1 g_54_78 (.ZN (n_54_78), .A (n_58_76), .B (n_64_73), .C1 (n_61_72), .C2 (n_55_75) );
AOI211_X1 g_53_76 (.ZN (n_53_76), .A (n_56_77), .B (n_62_74), .C1 (n_63_71), .C2 (n_57_74) );
AOI211_X1 g_51_77 (.ZN (n_51_77), .A (n_54_78), .B (n_60_75), .C1 (n_64_73), .C2 (n_59_73) );
AOI211_X1 g_49_78 (.ZN (n_49_78), .A (n_53_76), .B (n_58_76), .C1 (n_62_74), .C2 (n_61_72) );
AOI211_X1 g_47_79 (.ZN (n_47_79), .A (n_51_77), .B (n_56_77), .C1 (n_60_75), .C2 (n_63_71) );
AOI211_X1 g_45_80 (.ZN (n_45_80), .A (n_49_78), .B (n_54_78), .C1 (n_58_76), .C2 (n_64_73) );
AOI211_X1 g_43_81 (.ZN (n_43_81), .A (n_47_79), .B (n_53_76), .C1 (n_56_77), .C2 (n_62_74) );
AOI211_X1 g_41_82 (.ZN (n_41_82), .A (n_45_80), .B (n_51_77), .C1 (n_54_78), .C2 (n_60_75) );
AOI211_X1 g_42_84 (.ZN (n_42_84), .A (n_43_81), .B (n_49_78), .C1 (n_53_76), .C2 (n_58_76) );
AOI211_X1 g_44_83 (.ZN (n_44_83), .A (n_41_82), .B (n_47_79), .C1 (n_51_77), .C2 (n_56_77) );
AOI211_X1 g_45_81 (.ZN (n_45_81), .A (n_42_84), .B (n_45_80), .C1 (n_49_78), .C2 (n_54_78) );
AOI211_X1 g_47_80 (.ZN (n_47_80), .A (n_44_83), .B (n_43_81), .C1 (n_47_79), .C2 (n_53_76) );
AOI211_X1 g_49_79 (.ZN (n_49_79), .A (n_45_81), .B (n_41_82), .C1 (n_45_80), .C2 (n_51_77) );
AOI211_X1 g_51_78 (.ZN (n_51_78), .A (n_47_80), .B (n_42_84), .C1 (n_43_81), .C2 (n_49_78) );
AOI211_X1 g_53_77 (.ZN (n_53_77), .A (n_49_79), .B (n_44_83), .C1 (n_41_82), .C2 (n_47_79) );
AOI211_X1 g_52_79 (.ZN (n_52_79), .A (n_51_78), .B (n_45_81), .C1 (n_42_84), .C2 (n_45_80) );
AOI211_X1 g_50_80 (.ZN (n_50_80), .A (n_53_77), .B (n_47_80), .C1 (n_44_83), .C2 (n_43_81) );
AOI211_X1 g_48_81 (.ZN (n_48_81), .A (n_52_79), .B (n_49_79), .C1 (n_45_81), .C2 (n_41_82) );
AOI211_X1 g_46_82 (.ZN (n_46_82), .A (n_50_80), .B (n_51_78), .C1 (n_47_80), .C2 (n_42_84) );
AOI211_X1 g_45_84 (.ZN (n_45_84), .A (n_48_81), .B (n_53_77), .C1 (n_49_79), .C2 (n_44_83) );
AOI211_X1 g_44_82 (.ZN (n_44_82), .A (n_46_82), .B (n_52_79), .C1 (n_51_78), .C2 (n_45_81) );
AOI211_X1 g_46_81 (.ZN (n_46_81), .A (n_45_84), .B (n_50_80), .C1 (n_53_77), .C2 (n_47_80) );
AOI211_X1 g_48_80 (.ZN (n_48_80), .A (n_44_82), .B (n_48_81), .C1 (n_52_79), .C2 (n_49_79) );
AOI211_X1 g_50_79 (.ZN (n_50_79), .A (n_46_81), .B (n_46_82), .C1 (n_50_80), .C2 (n_51_78) );
AOI211_X1 g_52_78 (.ZN (n_52_78), .A (n_48_80), .B (n_45_84), .C1 (n_48_81), .C2 (n_53_77) );
AOI211_X1 g_54_77 (.ZN (n_54_77), .A (n_50_79), .B (n_44_82), .C1 (n_46_82), .C2 (n_52_79) );
AOI211_X1 g_56_76 (.ZN (n_56_76), .A (n_52_78), .B (n_46_81), .C1 (n_45_84), .C2 (n_50_80) );
AOI211_X1 g_58_75 (.ZN (n_58_75), .A (n_54_77), .B (n_48_80), .C1 (n_44_82), .C2 (n_48_81) );
AOI211_X1 g_60_74 (.ZN (n_60_74), .A (n_56_76), .B (n_50_79), .C1 (n_46_81), .C2 (n_46_82) );
AOI211_X1 g_62_73 (.ZN (n_62_73), .A (n_58_75), .B (n_52_78), .C1 (n_48_80), .C2 (n_45_84) );
AOI211_X1 g_64_72 (.ZN (n_64_72), .A (n_60_74), .B (n_54_77), .C1 (n_50_79), .C2 (n_44_82) );
AOI211_X1 g_66_71 (.ZN (n_66_71), .A (n_62_73), .B (n_56_76), .C1 (n_52_78), .C2 (n_46_81) );
AOI211_X1 g_68_70 (.ZN (n_68_70), .A (n_64_72), .B (n_58_75), .C1 (n_54_77), .C2 (n_48_80) );
AOI211_X1 g_70_69 (.ZN (n_70_69), .A (n_66_71), .B (n_60_74), .C1 (n_56_76), .C2 (n_50_79) );
AOI211_X1 g_72_68 (.ZN (n_72_68), .A (n_68_70), .B (n_62_73), .C1 (n_58_75), .C2 (n_52_78) );
AOI211_X1 g_74_67 (.ZN (n_74_67), .A (n_70_69), .B (n_64_72), .C1 (n_60_74), .C2 (n_54_77) );
AOI211_X1 g_76_66 (.ZN (n_76_66), .A (n_72_68), .B (n_66_71), .C1 (n_62_73), .C2 (n_56_76) );
AOI211_X1 g_78_65 (.ZN (n_78_65), .A (n_74_67), .B (n_68_70), .C1 (n_64_72), .C2 (n_58_75) );
AOI211_X1 g_77_67 (.ZN (n_77_67), .A (n_76_66), .B (n_70_69), .C1 (n_66_71), .C2 (n_60_74) );
AOI211_X1 g_79_66 (.ZN (n_79_66), .A (n_78_65), .B (n_72_68), .C1 (n_68_70), .C2 (n_62_73) );
AOI211_X1 g_81_65 (.ZN (n_81_65), .A (n_77_67), .B (n_74_67), .C1 (n_70_69), .C2 (n_64_72) );
AOI211_X1 g_83_64 (.ZN (n_83_64), .A (n_79_66), .B (n_76_66), .C1 (n_72_68), .C2 (n_66_71) );
AOI211_X1 g_85_63 (.ZN (n_85_63), .A (n_81_65), .B (n_78_65), .C1 (n_74_67), .C2 (n_68_70) );
AOI211_X1 g_87_62 (.ZN (n_87_62), .A (n_83_64), .B (n_77_67), .C1 (n_76_66), .C2 (n_70_69) );
AOI211_X1 g_89_61 (.ZN (n_89_61), .A (n_85_63), .B (n_79_66), .C1 (n_78_65), .C2 (n_72_68) );
AOI211_X1 g_91_60 (.ZN (n_91_60), .A (n_87_62), .B (n_81_65), .C1 (n_77_67), .C2 (n_74_67) );
AOI211_X1 g_93_61 (.ZN (n_93_61), .A (n_89_61), .B (n_83_64), .C1 (n_79_66), .C2 (n_76_66) );
AOI211_X1 g_94_63 (.ZN (n_94_63), .A (n_91_60), .B (n_85_63), .C1 (n_81_65), .C2 (n_78_65) );
AOI211_X1 g_92_62 (.ZN (n_92_62), .A (n_93_61), .B (n_87_62), .C1 (n_83_64), .C2 (n_77_67) );
AOI211_X1 g_90_63 (.ZN (n_90_63), .A (n_94_63), .B (n_89_61), .C1 (n_85_63), .C2 (n_79_66) );
AOI211_X1 g_91_61 (.ZN (n_91_61), .A (n_92_62), .B (n_91_60), .C1 (n_87_62), .C2 (n_81_65) );
AOI211_X1 g_93_62 (.ZN (n_93_62), .A (n_90_63), .B (n_93_61), .C1 (n_89_61), .C2 (n_83_64) );
AOI211_X1 g_94_64 (.ZN (n_94_64), .A (n_91_61), .B (n_94_63), .C1 (n_91_60), .C2 (n_85_63) );
AOI211_X1 g_92_63 (.ZN (n_92_63), .A (n_93_62), .B (n_92_62), .C1 (n_93_61), .C2 (n_87_62) );
AOI211_X1 g_94_62 (.ZN (n_94_62), .A (n_94_64), .B (n_90_63), .C1 (n_94_63), .C2 (n_89_61) );
AOI211_X1 g_95_64 (.ZN (n_95_64), .A (n_92_63), .B (n_91_61), .C1 (n_92_62), .C2 (n_91_60) );
AOI211_X1 g_93_65 (.ZN (n_93_65), .A (n_94_62), .B (n_93_62), .C1 (n_90_63), .C2 (n_93_61) );
AOI211_X1 g_94_67 (.ZN (n_94_67), .A (n_95_64), .B (n_94_64), .C1 (n_91_61), .C2 (n_94_63) );
AOI211_X1 g_95_65 (.ZN (n_95_65), .A (n_93_65), .B (n_92_63), .C1 (n_93_62), .C2 (n_92_62) );
AOI211_X1 g_93_64 (.ZN (n_93_64), .A (n_94_67), .B (n_94_62), .C1 (n_94_64), .C2 (n_90_63) );
AOI211_X1 g_91_63 (.ZN (n_91_63), .A (n_95_65), .B (n_95_64), .C1 (n_92_63), .C2 (n_91_61) );
AOI211_X1 g_92_61 (.ZN (n_92_61), .A (n_93_64), .B (n_93_65), .C1 (n_94_62), .C2 (n_93_62) );
AOI211_X1 g_90_60 (.ZN (n_90_60), .A (n_91_63), .B (n_94_67), .C1 (n_95_64), .C2 (n_94_64) );
AOI211_X1 g_88_61 (.ZN (n_88_61), .A (n_92_61), .B (n_95_65), .C1 (n_93_65), .C2 (n_92_63) );
AOI211_X1 g_90_62 (.ZN (n_90_62), .A (n_90_60), .B (n_93_64), .C1 (n_94_67), .C2 (n_94_62) );
AOI211_X1 g_89_64 (.ZN (n_89_64), .A (n_88_61), .B (n_91_63), .C1 (n_95_65), .C2 (n_95_64) );
AOI211_X1 g_91_65 (.ZN (n_91_65), .A (n_90_62), .B (n_92_61), .C1 (n_93_64), .C2 (n_93_65) );
AOI211_X1 g_93_66 (.ZN (n_93_66), .A (n_89_64), .B (n_90_60), .C1 (n_91_63), .C2 (n_94_67) );
AOI211_X1 g_92_64 (.ZN (n_92_64), .A (n_91_65), .B (n_88_61), .C1 (n_92_61), .C2 (n_95_65) );
AOI211_X1 g_91_62 (.ZN (n_91_62), .A (n_93_66), .B (n_90_62), .C1 (n_90_60), .C2 (n_93_64) );
AOI211_X1 g_93_63 (.ZN (n_93_63), .A (n_92_64), .B (n_89_64), .C1 (n_88_61), .C2 (n_91_63) );
AOI211_X1 g_94_65 (.ZN (n_94_65), .A (n_91_62), .B (n_91_65), .C1 (n_90_62), .C2 (n_92_61) );
AOI211_X1 g_95_67 (.ZN (n_95_67), .A (n_93_63), .B (n_93_66), .C1 (n_89_64), .C2 (n_90_60) );
AOI211_X1 g_96_69 (.ZN (n_96_69), .A (n_94_65), .B (n_92_64), .C1 (n_91_65), .C2 (n_88_61) );
AOI211_X1 g_97_71 (.ZN (n_97_71), .A (n_95_67), .B (n_91_62), .C1 (n_93_66), .C2 (n_90_62) );
AOI211_X1 g_98_73 (.ZN (n_98_73), .A (n_96_69), .B (n_93_63), .C1 (n_92_64), .C2 (n_89_64) );
AOI211_X1 g_99_75 (.ZN (n_99_75), .A (n_97_71), .B (n_94_65), .C1 (n_91_62), .C2 (n_91_65) );
AOI211_X1 g_100_77 (.ZN (n_100_77), .A (n_98_73), .B (n_95_67), .C1 (n_93_63), .C2 (n_93_66) );
AOI211_X1 g_98_76 (.ZN (n_98_76), .A (n_99_75), .B (n_96_69), .C1 (n_94_65), .C2 (n_92_64) );
AOI211_X1 g_100_75 (.ZN (n_100_75), .A (n_100_77), .B (n_97_71), .C1 (n_95_67), .C2 (n_91_62) );
AOI211_X1 g_99_73 (.ZN (n_99_73), .A (n_98_76), .B (n_98_73), .C1 (n_96_69), .C2 (n_93_63) );
AOI211_X1 g_98_71 (.ZN (n_98_71), .A (n_100_75), .B (n_99_75), .C1 (n_97_71), .C2 (n_94_65) );
AOI211_X1 g_97_69 (.ZN (n_97_69), .A (n_99_73), .B (n_100_77), .C1 (n_98_73), .C2 (n_95_67) );
AOI211_X1 g_96_67 (.ZN (n_96_67), .A (n_98_71), .B (n_98_76), .C1 (n_99_75), .C2 (n_96_69) );
AOI211_X1 g_94_66 (.ZN (n_94_66), .A (n_97_69), .B (n_100_75), .C1 (n_100_77), .C2 (n_97_71) );
AOI211_X1 g_92_65 (.ZN (n_92_65), .A (n_96_67), .B (n_99_73), .C1 (n_98_76), .C2 (n_98_73) );
AOI211_X1 g_90_64 (.ZN (n_90_64), .A (n_94_66), .B (n_98_71), .C1 (n_100_75), .C2 (n_99_75) );
AOI211_X1 g_89_62 (.ZN (n_89_62), .A (n_92_65), .B (n_97_69), .C1 (n_99_73), .C2 (n_100_77) );
AOI211_X1 g_87_61 (.ZN (n_87_61), .A (n_90_64), .B (n_96_67), .C1 (n_98_71), .C2 (n_98_76) );
AOI211_X1 g_85_62 (.ZN (n_85_62), .A (n_89_62), .B (n_94_66), .C1 (n_97_69), .C2 (n_100_75) );
AOI211_X1 g_87_63 (.ZN (n_87_63), .A (n_87_61), .B (n_92_65), .C1 (n_96_67), .C2 (n_99_73) );
AOI211_X1 g_85_64 (.ZN (n_85_64), .A (n_85_62), .B (n_90_64), .C1 (n_94_66), .C2 (n_98_71) );
AOI211_X1 g_86_62 (.ZN (n_86_62), .A (n_87_63), .B (n_89_62), .C1 (n_92_65), .C2 (n_97_69) );
AOI211_X1 g_88_63 (.ZN (n_88_63), .A (n_85_64), .B (n_87_61), .C1 (n_90_64), .C2 (n_96_67) );
AOI211_X1 g_86_64 (.ZN (n_86_64), .A (n_86_62), .B (n_85_62), .C1 (n_89_62), .C2 (n_94_66) );
AOI211_X1 g_84_63 (.ZN (n_84_63), .A (n_88_63), .B (n_87_63), .C1 (n_87_61), .C2 (n_92_65) );
AOI211_X1 g_82_64 (.ZN (n_82_64), .A (n_86_64), .B (n_85_64), .C1 (n_85_62), .C2 (n_90_64) );
AOI211_X1 g_80_65 (.ZN (n_80_65), .A (n_84_63), .B (n_86_62), .C1 (n_87_63), .C2 (n_89_62) );
AOI211_X1 g_78_66 (.ZN (n_78_66), .A (n_82_64), .B (n_88_63), .C1 (n_85_64), .C2 (n_87_61) );
AOI211_X1 g_76_67 (.ZN (n_76_67), .A (n_80_65), .B (n_86_64), .C1 (n_86_62), .C2 (n_85_62) );
AOI211_X1 g_75_69 (.ZN (n_75_69), .A (n_78_66), .B (n_84_63), .C1 (n_88_63), .C2 (n_87_63) );
AOI211_X1 g_73_68 (.ZN (n_73_68), .A (n_76_67), .B (n_82_64), .C1 (n_86_64), .C2 (n_85_64) );
AOI211_X1 g_75_67 (.ZN (n_75_67), .A (n_75_69), .B (n_80_65), .C1 (n_84_63), .C2 (n_86_62) );
AOI211_X1 g_77_66 (.ZN (n_77_66), .A (n_73_68), .B (n_78_66), .C1 (n_82_64), .C2 (n_88_63) );
AOI211_X1 g_79_65 (.ZN (n_79_65), .A (n_75_67), .B (n_76_67), .C1 (n_80_65), .C2 (n_86_64) );
AOI211_X1 g_81_64 (.ZN (n_81_64), .A (n_77_66), .B (n_75_69), .C1 (n_78_66), .C2 (n_84_63) );
AOI211_X1 g_83_63 (.ZN (n_83_63), .A (n_79_65), .B (n_73_68), .C1 (n_76_67), .C2 (n_82_64) );
AOI211_X1 g_84_65 (.ZN (n_84_65), .A (n_81_64), .B (n_75_67), .C1 (n_75_69), .C2 (n_80_65) );
AOI211_X1 g_82_66 (.ZN (n_82_66), .A (n_83_63), .B (n_77_66), .C1 (n_73_68), .C2 (n_78_66) );
AOI211_X1 g_80_67 (.ZN (n_80_67), .A (n_84_65), .B (n_79_65), .C1 (n_75_67), .C2 (n_76_67) );
AOI211_X1 g_78_68 (.ZN (n_78_68), .A (n_82_66), .B (n_81_64), .C1 (n_77_66), .C2 (n_75_69) );
AOI211_X1 g_76_69 (.ZN (n_76_69), .A (n_80_67), .B (n_83_63), .C1 (n_79_65), .C2 (n_73_68) );
AOI211_X1 g_74_70 (.ZN (n_74_70), .A (n_78_68), .B (n_84_65), .C1 (n_81_64), .C2 (n_75_67) );
AOI211_X1 g_75_68 (.ZN (n_75_68), .A (n_76_69), .B (n_82_66), .C1 (n_83_63), .C2 (n_77_66) );
AOI211_X1 g_73_69 (.ZN (n_73_69), .A (n_74_70), .B (n_80_67), .C1 (n_84_65), .C2 (n_79_65) );
AOI211_X1 g_71_70 (.ZN (n_71_70), .A (n_75_68), .B (n_78_68), .C1 (n_82_66), .C2 (n_81_64) );
AOI211_X1 g_69_71 (.ZN (n_69_71), .A (n_73_69), .B (n_76_69), .C1 (n_80_67), .C2 (n_83_63) );
AOI211_X1 g_67_72 (.ZN (n_67_72), .A (n_71_70), .B (n_74_70), .C1 (n_78_68), .C2 (n_84_65) );
AOI211_X1 g_65_73 (.ZN (n_65_73), .A (n_69_71), .B (n_75_68), .C1 (n_76_69), .C2 (n_82_66) );
AOI211_X1 g_63_74 (.ZN (n_63_74), .A (n_67_72), .B (n_73_69), .C1 (n_74_70), .C2 (n_80_67) );
AOI211_X1 g_61_75 (.ZN (n_61_75), .A (n_65_73), .B (n_71_70), .C1 (n_75_68), .C2 (n_78_68) );
AOI211_X1 g_59_76 (.ZN (n_59_76), .A (n_63_74), .B (n_69_71), .C1 (n_73_69), .C2 (n_76_69) );
AOI211_X1 g_57_77 (.ZN (n_57_77), .A (n_61_75), .B (n_67_72), .C1 (n_71_70), .C2 (n_74_70) );
AOI211_X1 g_55_78 (.ZN (n_55_78), .A (n_59_76), .B (n_65_73), .C1 (n_69_71), .C2 (n_75_68) );
AOI211_X1 g_53_79 (.ZN (n_53_79), .A (n_57_77), .B (n_63_74), .C1 (n_67_72), .C2 (n_73_69) );
AOI211_X1 g_51_80 (.ZN (n_51_80), .A (n_55_78), .B (n_61_75), .C1 (n_65_73), .C2 (n_71_70) );
AOI211_X1 g_49_81 (.ZN (n_49_81), .A (n_53_79), .B (n_59_76), .C1 (n_63_74), .C2 (n_69_71) );
AOI211_X1 g_47_82 (.ZN (n_47_82), .A (n_51_80), .B (n_57_77), .C1 (n_61_75), .C2 (n_67_72) );
AOI211_X1 g_45_83 (.ZN (n_45_83), .A (n_49_81), .B (n_55_78), .C1 (n_59_76), .C2 (n_65_73) );
AOI211_X1 g_43_84 (.ZN (n_43_84), .A (n_47_82), .B (n_53_79), .C1 (n_57_77), .C2 (n_63_74) );
AOI211_X1 g_41_85 (.ZN (n_41_85), .A (n_45_83), .B (n_51_80), .C1 (n_55_78), .C2 (n_61_75) );
AOI211_X1 g_42_83 (.ZN (n_42_83), .A (n_43_84), .B (n_49_81), .C1 (n_53_79), .C2 (n_59_76) );
AOI211_X1 g_40_84 (.ZN (n_40_84), .A (n_41_85), .B (n_47_82), .C1 (n_51_80), .C2 (n_57_77) );
AOI211_X1 g_38_85 (.ZN (n_38_85), .A (n_42_83), .B (n_45_83), .C1 (n_49_81), .C2 (n_55_78) );
AOI211_X1 g_36_84 (.ZN (n_36_84), .A (n_40_84), .B (n_43_84), .C1 (n_47_82), .C2 (n_53_79) );
AOI211_X1 g_34_85 (.ZN (n_34_85), .A (n_38_85), .B (n_41_85), .C1 (n_45_83), .C2 (n_51_80) );
AOI211_X1 g_32_84 (.ZN (n_32_84), .A (n_36_84), .B (n_42_83), .C1 (n_43_84), .C2 (n_49_81) );
AOI211_X1 g_30_85 (.ZN (n_30_85), .A (n_34_85), .B (n_40_84), .C1 (n_41_85), .C2 (n_47_82) );
AOI211_X1 g_28_86 (.ZN (n_28_86), .A (n_32_84), .B (n_38_85), .C1 (n_42_83), .C2 (n_45_83) );
AOI211_X1 g_26_87 (.ZN (n_26_87), .A (n_30_85), .B (n_36_84), .C1 (n_40_84), .C2 (n_43_84) );
AOI211_X1 g_24_88 (.ZN (n_24_88), .A (n_28_86), .B (n_34_85), .C1 (n_38_85), .C2 (n_41_85) );
AOI211_X1 g_22_89 (.ZN (n_22_89), .A (n_26_87), .B (n_32_84), .C1 (n_36_84), .C2 (n_42_83) );
AOI211_X1 g_20_90 (.ZN (n_20_90), .A (n_24_88), .B (n_30_85), .C1 (n_34_85), .C2 (n_40_84) );
AOI211_X1 g_18_91 (.ZN (n_18_91), .A (n_22_89), .B (n_28_86), .C1 (n_32_84), .C2 (n_38_85) );
AOI211_X1 g_16_92 (.ZN (n_16_92), .A (n_20_90), .B (n_26_87), .C1 (n_30_85), .C2 (n_36_84) );
AOI211_X1 g_14_93 (.ZN (n_14_93), .A (n_18_91), .B (n_24_88), .C1 (n_28_86), .C2 (n_34_85) );
AOI211_X1 g_13_95 (.ZN (n_13_95), .A (n_16_92), .B (n_22_89), .C1 (n_26_87), .C2 (n_32_84) );
AOI211_X1 g_15_94 (.ZN (n_15_94), .A (n_14_93), .B (n_20_90), .C1 (n_24_88), .C2 (n_30_85) );
AOI211_X1 g_17_93 (.ZN (n_17_93), .A (n_13_95), .B (n_18_91), .C1 (n_22_89), .C2 (n_28_86) );
AOI211_X1 g_19_92 (.ZN (n_19_92), .A (n_15_94), .B (n_16_92), .C1 (n_20_90), .C2 (n_26_87) );
AOI211_X1 g_21_91 (.ZN (n_21_91), .A (n_17_93), .B (n_14_93), .C1 (n_18_91), .C2 (n_24_88) );
AOI211_X1 g_23_90 (.ZN (n_23_90), .A (n_19_92), .B (n_13_95), .C1 (n_16_92), .C2 (n_22_89) );
AOI211_X1 g_25_89 (.ZN (n_25_89), .A (n_21_91), .B (n_15_94), .C1 (n_14_93), .C2 (n_20_90) );
AOI211_X1 g_27_88 (.ZN (n_27_88), .A (n_23_90), .B (n_17_93), .C1 (n_13_95), .C2 (n_18_91) );
AOI211_X1 g_29_87 (.ZN (n_29_87), .A (n_25_89), .B (n_19_92), .C1 (n_15_94), .C2 (n_16_92) );
AOI211_X1 g_31_86 (.ZN (n_31_86), .A (n_27_88), .B (n_21_91), .C1 (n_17_93), .C2 (n_14_93) );
AOI211_X1 g_33_85 (.ZN (n_33_85), .A (n_29_87), .B (n_23_90), .C1 (n_19_92), .C2 (n_13_95) );
AOI211_X1 g_35_84 (.ZN (n_35_84), .A (n_31_86), .B (n_25_89), .C1 (n_21_91), .C2 (n_15_94) );
AOI211_X1 g_34_86 (.ZN (n_34_86), .A (n_33_85), .B (n_27_88), .C1 (n_23_90), .C2 (n_17_93) );
AOI211_X1 g_32_87 (.ZN (n_32_87), .A (n_35_84), .B (n_29_87), .C1 (n_25_89), .C2 (n_19_92) );
AOI211_X1 g_31_85 (.ZN (n_31_85), .A (n_34_86), .B (n_31_86), .C1 (n_27_88), .C2 (n_21_91) );
AOI211_X1 g_29_86 (.ZN (n_29_86), .A (n_32_87), .B (n_33_85), .C1 (n_29_87), .C2 (n_23_90) );
AOI211_X1 g_27_87 (.ZN (n_27_87), .A (n_31_85), .B (n_35_84), .C1 (n_31_86), .C2 (n_25_89) );
AOI211_X1 g_25_88 (.ZN (n_25_88), .A (n_29_86), .B (n_34_86), .C1 (n_33_85), .C2 (n_27_88) );
AOI211_X1 g_23_89 (.ZN (n_23_89), .A (n_27_87), .B (n_32_87), .C1 (n_35_84), .C2 (n_29_87) );
AOI211_X1 g_21_90 (.ZN (n_21_90), .A (n_25_88), .B (n_31_85), .C1 (n_34_86), .C2 (n_31_86) );
AOI211_X1 g_19_91 (.ZN (n_19_91), .A (n_23_89), .B (n_29_86), .C1 (n_32_87), .C2 (n_33_85) );
AOI211_X1 g_17_92 (.ZN (n_17_92), .A (n_21_90), .B (n_27_87), .C1 (n_31_85), .C2 (n_35_84) );
AOI211_X1 g_15_93 (.ZN (n_15_93), .A (n_19_91), .B (n_25_88), .C1 (n_29_86), .C2 (n_34_86) );
AOI211_X1 g_13_94 (.ZN (n_13_94), .A (n_17_92), .B (n_23_89), .C1 (n_27_87), .C2 (n_32_87) );
AOI211_X1 g_12_96 (.ZN (n_12_96), .A (n_15_93), .B (n_21_90), .C1 (n_25_88), .C2 (n_31_85) );
AOI211_X1 g_11_98 (.ZN (n_11_98), .A (n_13_94), .B (n_19_91), .C1 (n_23_89), .C2 (n_29_86) );
AOI211_X1 g_12_100 (.ZN (n_12_100), .A (n_12_96), .B (n_17_92), .C1 (n_21_90), .C2 (n_27_87) );
AOI211_X1 g_13_98 (.ZN (n_13_98), .A (n_11_98), .B (n_15_93), .C1 (n_19_91), .C2 (n_25_88) );
AOI211_X1 g_14_96 (.ZN (n_14_96), .A (n_12_100), .B (n_13_94), .C1 (n_17_92), .C2 (n_23_89) );
AOI211_X1 g_16_95 (.ZN (n_16_95), .A (n_13_98), .B (n_12_96), .C1 (n_15_93), .C2 (n_21_90) );
AOI211_X1 g_18_94 (.ZN (n_18_94), .A (n_14_96), .B (n_11_98), .C1 (n_13_94), .C2 (n_19_91) );
AOI211_X1 g_20_93 (.ZN (n_20_93), .A (n_16_95), .B (n_12_100), .C1 (n_12_96), .C2 (n_17_92) );
AOI211_X1 g_18_92 (.ZN (n_18_92), .A (n_18_94), .B (n_13_98), .C1 (n_11_98), .C2 (n_15_93) );
AOI211_X1 g_20_91 (.ZN (n_20_91), .A (n_20_93), .B (n_14_96), .C1 (n_12_100), .C2 (n_13_94) );
AOI211_X1 g_22_90 (.ZN (n_22_90), .A (n_18_92), .B (n_16_95), .C1 (n_13_98), .C2 (n_12_96) );
AOI211_X1 g_24_89 (.ZN (n_24_89), .A (n_20_91), .B (n_18_94), .C1 (n_14_96), .C2 (n_11_98) );
AOI211_X1 g_23_91 (.ZN (n_23_91), .A (n_22_90), .B (n_20_93), .C1 (n_16_95), .C2 (n_12_100) );
AOI211_X1 g_25_90 (.ZN (n_25_90), .A (n_24_89), .B (n_18_92), .C1 (n_18_94), .C2 (n_13_98) );
AOI211_X1 g_27_89 (.ZN (n_27_89), .A (n_23_91), .B (n_20_91), .C1 (n_20_93), .C2 (n_14_96) );
AOI211_X1 g_29_88 (.ZN (n_29_88), .A (n_25_90), .B (n_22_90), .C1 (n_18_92), .C2 (n_16_95) );
AOI211_X1 g_31_87 (.ZN (n_31_87), .A (n_27_89), .B (n_24_89), .C1 (n_20_91), .C2 (n_18_94) );
AOI211_X1 g_33_86 (.ZN (n_33_86), .A (n_29_88), .B (n_23_91), .C1 (n_22_90), .C2 (n_20_93) );
AOI211_X1 g_35_87 (.ZN (n_35_87), .A (n_31_87), .B (n_25_90), .C1 (n_24_89), .C2 (n_18_92) );
AOI211_X1 g_37_86 (.ZN (n_37_86), .A (n_33_86), .B (n_27_89), .C1 (n_23_91), .C2 (n_20_91) );
AOI211_X1 g_39_85 (.ZN (n_39_85), .A (n_35_87), .B (n_29_88), .C1 (n_25_90), .C2 (n_22_90) );
AOI211_X1 g_41_84 (.ZN (n_41_84), .A (n_37_86), .B (n_31_87), .C1 (n_27_89), .C2 (n_24_89) );
AOI211_X1 g_43_83 (.ZN (n_43_83), .A (n_39_85), .B (n_33_86), .C1 (n_29_88), .C2 (n_23_91) );
AOI211_X1 g_45_82 (.ZN (n_45_82), .A (n_41_84), .B (n_35_87), .C1 (n_31_87), .C2 (n_25_90) );
AOI211_X1 g_47_81 (.ZN (n_47_81), .A (n_43_83), .B (n_37_86), .C1 (n_33_86), .C2 (n_27_89) );
AOI211_X1 g_49_80 (.ZN (n_49_80), .A (n_45_82), .B (n_39_85), .C1 (n_35_87), .C2 (n_29_88) );
AOI211_X1 g_51_79 (.ZN (n_51_79), .A (n_47_81), .B (n_41_84), .C1 (n_37_86), .C2 (n_31_87) );
AOI211_X1 g_53_78 (.ZN (n_53_78), .A (n_49_80), .B (n_43_83), .C1 (n_39_85), .C2 (n_33_86) );
AOI211_X1 g_52_80 (.ZN (n_52_80), .A (n_51_79), .B (n_45_82), .C1 (n_41_84), .C2 (n_35_87) );
AOI211_X1 g_54_79 (.ZN (n_54_79), .A (n_53_78), .B (n_47_81), .C1 (n_43_83), .C2 (n_37_86) );
AOI211_X1 g_56_78 (.ZN (n_56_78), .A (n_52_80), .B (n_49_80), .C1 (n_45_82), .C2 (n_39_85) );
AOI211_X1 g_58_77 (.ZN (n_58_77), .A (n_54_79), .B (n_51_79), .C1 (n_47_81), .C2 (n_41_84) );
AOI211_X1 g_60_76 (.ZN (n_60_76), .A (n_56_78), .B (n_53_78), .C1 (n_49_80), .C2 (n_43_83) );
AOI211_X1 g_61_74 (.ZN (n_61_74), .A (n_58_77), .B (n_52_80), .C1 (n_51_79), .C2 (n_45_82) );
AOI211_X1 g_63_73 (.ZN (n_63_73), .A (n_60_76), .B (n_54_79), .C1 (n_53_78), .C2 (n_47_81) );
AOI211_X1 g_65_72 (.ZN (n_65_72), .A (n_61_74), .B (n_56_78), .C1 (n_52_80), .C2 (n_49_80) );
AOI211_X1 g_64_74 (.ZN (n_64_74), .A (n_63_73), .B (n_58_77), .C1 (n_54_79), .C2 (n_51_79) );
AOI211_X1 g_62_75 (.ZN (n_62_75), .A (n_65_72), .B (n_60_76), .C1 (n_56_78), .C2 (n_53_78) );
AOI211_X1 g_61_77 (.ZN (n_61_77), .A (n_64_74), .B (n_61_74), .C1 (n_58_77), .C2 (n_52_80) );
AOI211_X1 g_63_76 (.ZN (n_63_76), .A (n_62_75), .B (n_63_73), .C1 (n_60_76), .C2 (n_54_79) );
AOI211_X1 g_65_75 (.ZN (n_65_75), .A (n_61_77), .B (n_65_72), .C1 (n_61_74), .C2 (n_56_78) );
AOI211_X1 g_66_73 (.ZN (n_66_73), .A (n_63_76), .B (n_64_74), .C1 (n_63_73), .C2 (n_58_77) );
AOI211_X1 g_68_72 (.ZN (n_68_72), .A (n_65_75), .B (n_62_75), .C1 (n_65_72), .C2 (n_60_76) );
AOI211_X1 g_69_70 (.ZN (n_69_70), .A (n_66_73), .B (n_61_77), .C1 (n_64_74), .C2 (n_61_74) );
AOI211_X1 g_71_69 (.ZN (n_71_69), .A (n_68_72), .B (n_63_76), .C1 (n_62_75), .C2 (n_63_73) );
AOI211_X1 g_70_71 (.ZN (n_70_71), .A (n_69_70), .B (n_65_75), .C1 (n_61_77), .C2 (n_65_72) );
AOI211_X1 g_72_70 (.ZN (n_72_70), .A (n_71_69), .B (n_66_73), .C1 (n_63_76), .C2 (n_64_74) );
AOI211_X1 g_74_69 (.ZN (n_74_69), .A (n_70_71), .B (n_68_72), .C1 (n_65_75), .C2 (n_62_75) );
AOI211_X1 g_76_68 (.ZN (n_76_68), .A (n_72_70), .B (n_69_70), .C1 (n_66_73), .C2 (n_61_77) );
AOI211_X1 g_78_67 (.ZN (n_78_67), .A (n_74_69), .B (n_71_69), .C1 (n_68_72), .C2 (n_63_76) );
AOI211_X1 g_80_66 (.ZN (n_80_66), .A (n_76_68), .B (n_70_71), .C1 (n_69_70), .C2 (n_65_75) );
AOI211_X1 g_82_65 (.ZN (n_82_65), .A (n_78_67), .B (n_72_70), .C1 (n_71_69), .C2 (n_66_73) );
AOI211_X1 g_84_64 (.ZN (n_84_64), .A (n_80_66), .B (n_74_69), .C1 (n_70_71), .C2 (n_68_72) );
AOI211_X1 g_86_63 (.ZN (n_86_63), .A (n_82_65), .B (n_76_68), .C1 (n_72_70), .C2 (n_69_70) );
AOI211_X1 g_87_65 (.ZN (n_87_65), .A (n_84_64), .B (n_78_67), .C1 (n_74_69), .C2 (n_71_69) );
AOI211_X1 g_85_66 (.ZN (n_85_66), .A (n_86_63), .B (n_80_66), .C1 (n_76_68), .C2 (n_70_71) );
AOI211_X1 g_83_65 (.ZN (n_83_65), .A (n_87_65), .B (n_82_65), .C1 (n_78_67), .C2 (n_72_70) );
AOI211_X1 g_81_66 (.ZN (n_81_66), .A (n_85_66), .B (n_84_64), .C1 (n_80_66), .C2 (n_74_69) );
AOI211_X1 g_79_67 (.ZN (n_79_67), .A (n_83_65), .B (n_86_63), .C1 (n_82_65), .C2 (n_76_68) );
AOI211_X1 g_77_68 (.ZN (n_77_68), .A (n_81_66), .B (n_87_65), .C1 (n_84_64), .C2 (n_78_67) );
AOI211_X1 g_76_70 (.ZN (n_76_70), .A (n_79_67), .B (n_85_66), .C1 (n_86_63), .C2 (n_80_66) );
AOI211_X1 g_78_69 (.ZN (n_78_69), .A (n_77_68), .B (n_83_65), .C1 (n_87_65), .C2 (n_82_65) );
AOI211_X1 g_80_68 (.ZN (n_80_68), .A (n_76_70), .B (n_81_66), .C1 (n_85_66), .C2 (n_84_64) );
AOI211_X1 g_82_67 (.ZN (n_82_67), .A (n_78_69), .B (n_79_67), .C1 (n_83_65), .C2 (n_86_63) );
AOI211_X1 g_84_66 (.ZN (n_84_66), .A (n_80_68), .B (n_77_68), .C1 (n_81_66), .C2 (n_87_65) );
AOI211_X1 g_86_65 (.ZN (n_86_65), .A (n_82_67), .B (n_76_70), .C1 (n_79_67), .C2 (n_85_66) );
AOI211_X1 g_88_64 (.ZN (n_88_64), .A (n_84_66), .B (n_78_69), .C1 (n_77_68), .C2 (n_83_65) );
AOI211_X1 g_89_66 (.ZN (n_89_66), .A (n_86_65), .B (n_80_68), .C1 (n_76_70), .C2 (n_81_66) );
AOI211_X1 g_87_67 (.ZN (n_87_67), .A (n_88_64), .B (n_82_67), .C1 (n_78_69), .C2 (n_79_67) );
AOI211_X1 g_88_65 (.ZN (n_88_65), .A (n_89_66), .B (n_84_66), .C1 (n_80_68), .C2 (n_77_68) );
AOI211_X1 g_89_63 (.ZN (n_89_63), .A (n_87_67), .B (n_86_65), .C1 (n_82_67), .C2 (n_76_70) );
AOI211_X1 g_91_64 (.ZN (n_91_64), .A (n_88_65), .B (n_88_64), .C1 (n_84_66), .C2 (n_78_69) );
AOI211_X1 g_90_66 (.ZN (n_90_66), .A (n_89_63), .B (n_89_66), .C1 (n_86_65), .C2 (n_80_68) );
AOI211_X1 g_92_67 (.ZN (n_92_67), .A (n_91_64), .B (n_87_67), .C1 (n_88_64), .C2 (n_82_67) );
AOI211_X1 g_94_68 (.ZN (n_94_68), .A (n_90_66), .B (n_88_65), .C1 (n_89_66), .C2 (n_84_66) );
AOI211_X1 g_95_70 (.ZN (n_95_70), .A (n_92_67), .B (n_89_63), .C1 (n_87_67), .C2 (n_86_65) );
AOI211_X1 g_96_72 (.ZN (n_96_72), .A (n_94_68), .B (n_91_64), .C1 (n_88_65), .C2 (n_88_64) );
AOI211_X1 g_97_74 (.ZN (n_97_74), .A (n_95_70), .B (n_90_66), .C1 (n_89_63), .C2 (n_89_66) );
AOI211_X1 g_95_73 (.ZN (n_95_73), .A (n_96_72), .B (n_92_67), .C1 (n_91_64), .C2 (n_87_67) );
AOI211_X1 g_97_72 (.ZN (n_97_72), .A (n_97_74), .B (n_94_68), .C1 (n_90_66), .C2 (n_88_65) );
AOI211_X1 g_98_74 (.ZN (n_98_74), .A (n_95_73), .B (n_95_70), .C1 (n_92_67), .C2 (n_89_63) );
AOI211_X1 g_96_73 (.ZN (n_96_73), .A (n_97_72), .B (n_96_72), .C1 (n_94_68), .C2 (n_91_64) );
AOI211_X1 g_95_71 (.ZN (n_95_71), .A (n_98_74), .B (n_97_74), .C1 (n_95_70), .C2 (n_90_66) );
AOI211_X1 g_94_69 (.ZN (n_94_69), .A (n_96_73), .B (n_95_73), .C1 (n_96_72), .C2 (n_92_67) );
AOI211_X1 g_96_70 (.ZN (n_96_70), .A (n_95_71), .B (n_97_72), .C1 (n_97_74), .C2 (n_94_68) );
AOI211_X1 g_95_68 (.ZN (n_95_68), .A (n_94_69), .B (n_98_74), .C1 (n_95_73), .C2 (n_95_70) );
AOI211_X1 g_93_67 (.ZN (n_93_67), .A (n_96_70), .B (n_96_73), .C1 (n_97_72), .C2 (n_96_72) );
AOI211_X1 g_91_66 (.ZN (n_91_66), .A (n_95_68), .B (n_95_71), .C1 (n_98_74), .C2 (n_97_74) );
AOI211_X1 g_89_65 (.ZN (n_89_65), .A (n_93_67), .B (n_94_69), .C1 (n_96_73), .C2 (n_95_73) );
AOI211_X1 g_87_64 (.ZN (n_87_64), .A (n_91_66), .B (n_96_70), .C1 (n_95_71), .C2 (n_97_72) );
AOI211_X1 g_85_65 (.ZN (n_85_65), .A (n_89_65), .B (n_95_68), .C1 (n_94_69), .C2 (n_98_74) );
AOI211_X1 g_83_66 (.ZN (n_83_66), .A (n_87_64), .B (n_93_67), .C1 (n_96_70), .C2 (n_96_73) );
AOI211_X1 g_81_67 (.ZN (n_81_67), .A (n_85_65), .B (n_91_66), .C1 (n_95_68), .C2 (n_95_71) );
AOI211_X1 g_79_68 (.ZN (n_79_68), .A (n_83_66), .B (n_89_65), .C1 (n_93_67), .C2 (n_94_69) );
AOI211_X1 g_77_69 (.ZN (n_77_69), .A (n_81_67), .B (n_87_64), .C1 (n_91_66), .C2 (n_96_70) );
AOI211_X1 g_75_70 (.ZN (n_75_70), .A (n_79_68), .B (n_85_65), .C1 (n_89_65), .C2 (n_95_68) );
AOI211_X1 g_73_71 (.ZN (n_73_71), .A (n_77_69), .B (n_83_66), .C1 (n_87_64), .C2 (n_93_67) );
AOI211_X1 g_71_72 (.ZN (n_71_72), .A (n_75_70), .B (n_81_67), .C1 (n_85_65), .C2 (n_91_66) );
AOI211_X1 g_69_73 (.ZN (n_69_73), .A (n_73_71), .B (n_79_68), .C1 (n_83_66), .C2 (n_89_65) );
AOI211_X1 g_67_74 (.ZN (n_67_74), .A (n_71_72), .B (n_77_69), .C1 (n_81_67), .C2 (n_87_64) );
AOI211_X1 g_66_76 (.ZN (n_66_76), .A (n_69_73), .B (n_75_70), .C1 (n_79_68), .C2 (n_85_65) );
AOI211_X1 g_65_74 (.ZN (n_65_74), .A (n_67_74), .B (n_73_71), .C1 (n_77_69), .C2 (n_83_66) );
AOI211_X1 g_67_73 (.ZN (n_67_73), .A (n_66_76), .B (n_71_72), .C1 (n_75_70), .C2 (n_81_67) );
AOI211_X1 g_69_72 (.ZN (n_69_72), .A (n_65_74), .B (n_69_73), .C1 (n_73_71), .C2 (n_79_68) );
AOI211_X1 g_71_71 (.ZN (n_71_71), .A (n_67_73), .B (n_67_74), .C1 (n_71_72), .C2 (n_77_69) );
AOI211_X1 g_73_70 (.ZN (n_73_70), .A (n_69_72), .B (n_66_76), .C1 (n_69_73), .C2 (n_75_70) );
AOI211_X1 g_72_72 (.ZN (n_72_72), .A (n_71_71), .B (n_65_74), .C1 (n_67_74), .C2 (n_73_71) );
AOI211_X1 g_74_71 (.ZN (n_74_71), .A (n_73_70), .B (n_67_73), .C1 (n_66_76), .C2 (n_71_72) );
AOI211_X1 g_73_73 (.ZN (n_73_73), .A (n_72_72), .B (n_69_72), .C1 (n_65_74), .C2 (n_69_73) );
AOI211_X1 g_72_71 (.ZN (n_72_71), .A (n_74_71), .B (n_71_71), .C1 (n_67_73), .C2 (n_67_74) );
AOI211_X1 g_70_72 (.ZN (n_70_72), .A (n_73_73), .B (n_73_70), .C1 (n_69_72), .C2 (n_66_76) );
AOI211_X1 g_68_73 (.ZN (n_68_73), .A (n_72_71), .B (n_72_72), .C1 (n_71_71), .C2 (n_65_74) );
AOI211_X1 g_66_74 (.ZN (n_66_74), .A (n_70_72), .B (n_74_71), .C1 (n_73_70), .C2 (n_67_73) );
AOI211_X1 g_64_75 (.ZN (n_64_75), .A (n_68_73), .B (n_73_73), .C1 (n_72_72), .C2 (n_69_72) );
AOI211_X1 g_62_76 (.ZN (n_62_76), .A (n_66_74), .B (n_72_71), .C1 (n_74_71), .C2 (n_71_71) );
AOI211_X1 g_60_77 (.ZN (n_60_77), .A (n_64_75), .B (n_70_72), .C1 (n_73_73), .C2 (n_73_70) );
AOI211_X1 g_58_78 (.ZN (n_58_78), .A (n_62_76), .B (n_68_73), .C1 (n_72_71), .C2 (n_72_72) );
AOI211_X1 g_56_79 (.ZN (n_56_79), .A (n_60_77), .B (n_66_74), .C1 (n_70_72), .C2 (n_74_71) );
AOI211_X1 g_54_80 (.ZN (n_54_80), .A (n_58_78), .B (n_64_75), .C1 (n_68_73), .C2 (n_73_73) );
AOI211_X1 g_52_81 (.ZN (n_52_81), .A (n_56_79), .B (n_62_76), .C1 (n_66_74), .C2 (n_72_71) );
AOI211_X1 g_50_82 (.ZN (n_50_82), .A (n_54_80), .B (n_60_77), .C1 (n_64_75), .C2 (n_70_72) );
AOI211_X1 g_48_83 (.ZN (n_48_83), .A (n_52_81), .B (n_58_78), .C1 (n_62_76), .C2 (n_68_73) );
AOI211_X1 g_46_84 (.ZN (n_46_84), .A (n_50_82), .B (n_56_79), .C1 (n_60_77), .C2 (n_66_74) );
AOI211_X1 g_44_85 (.ZN (n_44_85), .A (n_48_83), .B (n_54_80), .C1 (n_58_78), .C2 (n_64_75) );
AOI211_X1 g_42_86 (.ZN (n_42_86), .A (n_46_84), .B (n_52_81), .C1 (n_56_79), .C2 (n_62_76) );
AOI211_X1 g_40_87 (.ZN (n_40_87), .A (n_44_85), .B (n_50_82), .C1 (n_54_80), .C2 (n_60_77) );
AOI211_X1 g_38_88 (.ZN (n_38_88), .A (n_42_86), .B (n_48_83), .C1 (n_52_81), .C2 (n_58_78) );
AOI211_X1 g_39_86 (.ZN (n_39_86), .A (n_40_87), .B (n_46_84), .C1 (n_50_82), .C2 (n_56_79) );
AOI211_X1 g_37_85 (.ZN (n_37_85), .A (n_38_88), .B (n_44_85), .C1 (n_48_83), .C2 (n_54_80) );
AOI211_X1 g_36_87 (.ZN (n_36_87), .A (n_39_86), .B (n_42_86), .C1 (n_46_84), .C2 (n_52_81) );
AOI211_X1 g_34_88 (.ZN (n_34_88), .A (n_37_85), .B (n_40_87), .C1 (n_44_85), .C2 (n_50_82) );
AOI211_X1 g_35_86 (.ZN (n_35_86), .A (n_36_87), .B (n_38_88), .C1 (n_42_86), .C2 (n_48_83) );
AOI211_X1 g_33_87 (.ZN (n_33_87), .A (n_34_88), .B (n_39_86), .C1 (n_40_87), .C2 (n_46_84) );
AOI211_X1 g_31_88 (.ZN (n_31_88), .A (n_35_86), .B (n_37_85), .C1 (n_38_88), .C2 (n_44_85) );
AOI211_X1 g_32_86 (.ZN (n_32_86), .A (n_33_87), .B (n_36_87), .C1 (n_39_86), .C2 (n_42_86) );
AOI211_X1 g_30_87 (.ZN (n_30_87), .A (n_31_88), .B (n_34_88), .C1 (n_37_85), .C2 (n_40_87) );
AOI211_X1 g_28_88 (.ZN (n_28_88), .A (n_32_86), .B (n_35_86), .C1 (n_36_87), .C2 (n_38_88) );
AOI211_X1 g_26_89 (.ZN (n_26_89), .A (n_30_87), .B (n_33_87), .C1 (n_34_88), .C2 (n_39_86) );
AOI211_X1 g_24_90 (.ZN (n_24_90), .A (n_28_88), .B (n_31_88), .C1 (n_35_86), .C2 (n_37_85) );
AOI211_X1 g_22_91 (.ZN (n_22_91), .A (n_26_89), .B (n_32_86), .C1 (n_33_87), .C2 (n_36_87) );
AOI211_X1 g_20_92 (.ZN (n_20_92), .A (n_24_90), .B (n_30_87), .C1 (n_31_88), .C2 (n_34_88) );
AOI211_X1 g_18_93 (.ZN (n_18_93), .A (n_22_91), .B (n_28_88), .C1 (n_32_86), .C2 (n_35_86) );
AOI211_X1 g_16_94 (.ZN (n_16_94), .A (n_20_92), .B (n_26_89), .C1 (n_30_87), .C2 (n_33_87) );
AOI211_X1 g_14_95 (.ZN (n_14_95), .A (n_18_93), .B (n_24_90), .C1 (n_28_88), .C2 (n_31_88) );
AOI211_X1 g_13_97 (.ZN (n_13_97), .A (n_16_94), .B (n_22_91), .C1 (n_26_89), .C2 (n_32_86) );
AOI211_X1 g_15_96 (.ZN (n_15_96), .A (n_14_95), .B (n_20_92), .C1 (n_24_90), .C2 (n_30_87) );
AOI211_X1 g_17_95 (.ZN (n_17_95), .A (n_13_97), .B (n_18_93), .C1 (n_22_91), .C2 (n_28_88) );
AOI211_X1 g_19_94 (.ZN (n_19_94), .A (n_15_96), .B (n_16_94), .C1 (n_20_92), .C2 (n_26_89) );
AOI211_X1 g_21_93 (.ZN (n_21_93), .A (n_17_95), .B (n_14_95), .C1 (n_18_93), .C2 (n_24_90) );
AOI211_X1 g_23_92 (.ZN (n_23_92), .A (n_19_94), .B (n_13_97), .C1 (n_16_94), .C2 (n_22_91) );
AOI211_X1 g_25_91 (.ZN (n_25_91), .A (n_21_93), .B (n_15_96), .C1 (n_14_95), .C2 (n_20_92) );
AOI211_X1 g_27_90 (.ZN (n_27_90), .A (n_23_92), .B (n_17_95), .C1 (n_13_97), .C2 (n_18_93) );
AOI211_X1 g_29_89 (.ZN (n_29_89), .A (n_25_91), .B (n_19_94), .C1 (n_15_96), .C2 (n_16_94) );
AOI211_X1 g_28_91 (.ZN (n_28_91), .A (n_27_90), .B (n_21_93), .C1 (n_17_95), .C2 (n_14_95) );
AOI211_X1 g_26_90 (.ZN (n_26_90), .A (n_29_89), .B (n_23_92), .C1 (n_19_94), .C2 (n_13_97) );
AOI211_X1 g_28_89 (.ZN (n_28_89), .A (n_28_91), .B (n_25_91), .C1 (n_21_93), .C2 (n_15_96) );
AOI211_X1 g_30_88 (.ZN (n_30_88), .A (n_26_90), .B (n_27_90), .C1 (n_23_92), .C2 (n_17_95) );
AOI211_X1 g_32_89 (.ZN (n_32_89), .A (n_28_89), .B (n_29_89), .C1 (n_25_91), .C2 (n_19_94) );
AOI211_X1 g_30_90 (.ZN (n_30_90), .A (n_30_88), .B (n_28_91), .C1 (n_27_90), .C2 (n_21_93) );
AOI211_X1 g_29_92 (.ZN (n_29_92), .A (n_32_89), .B (n_26_90), .C1 (n_29_89), .C2 (n_23_92) );
AOI211_X1 g_28_90 (.ZN (n_28_90), .A (n_30_90), .B (n_28_89), .C1 (n_28_91), .C2 (n_25_91) );
AOI211_X1 g_30_89 (.ZN (n_30_89), .A (n_29_92), .B (n_30_88), .C1 (n_26_90), .C2 (n_27_90) );
AOI211_X1 g_32_88 (.ZN (n_32_88), .A (n_28_90), .B (n_32_89), .C1 (n_28_89), .C2 (n_29_89) );
AOI211_X1 g_34_87 (.ZN (n_34_87), .A (n_30_89), .B (n_30_90), .C1 (n_30_88), .C2 (n_28_91) );
AOI211_X1 g_36_86 (.ZN (n_36_86), .A (n_32_88), .B (n_29_92), .C1 (n_32_89), .C2 (n_26_90) );
AOI211_X1 g_35_88 (.ZN (n_35_88), .A (n_34_87), .B (n_28_90), .C1 (n_30_90), .C2 (n_28_89) );
AOI211_X1 g_37_87 (.ZN (n_37_87), .A (n_36_86), .B (n_30_89), .C1 (n_29_92), .C2 (n_30_88) );
AOI211_X1 g_36_89 (.ZN (n_36_89), .A (n_35_88), .B (n_32_88), .C1 (n_28_90), .C2 (n_32_89) );
AOI211_X1 g_34_90 (.ZN (n_34_90), .A (n_37_87), .B (n_34_87), .C1 (n_30_89), .C2 (n_30_90) );
AOI211_X1 g_33_88 (.ZN (n_33_88), .A (n_36_89), .B (n_36_86), .C1 (n_32_88), .C2 (n_29_92) );
AOI211_X1 g_31_89 (.ZN (n_31_89), .A (n_34_90), .B (n_35_88), .C1 (n_34_87), .C2 (n_28_90) );
AOI211_X1 g_29_90 (.ZN (n_29_90), .A (n_33_88), .B (n_37_87), .C1 (n_36_86), .C2 (n_30_89) );
AOI211_X1 g_27_91 (.ZN (n_27_91), .A (n_31_89), .B (n_36_89), .C1 (n_35_88), .C2 (n_32_88) );
AOI211_X1 g_25_92 (.ZN (n_25_92), .A (n_29_90), .B (n_34_90), .C1 (n_37_87), .C2 (n_34_87) );
AOI211_X1 g_27_93 (.ZN (n_27_93), .A (n_27_91), .B (n_33_88), .C1 (n_36_89), .C2 (n_36_86) );
AOI211_X1 g_26_91 (.ZN (n_26_91), .A (n_25_92), .B (n_31_89), .C1 (n_34_90), .C2 (n_35_88) );
AOI211_X1 g_24_92 (.ZN (n_24_92), .A (n_27_93), .B (n_29_90), .C1 (n_33_88), .C2 (n_37_87) );
AOI211_X1 g_22_93 (.ZN (n_22_93), .A (n_26_91), .B (n_27_91), .C1 (n_31_89), .C2 (n_36_89) );
AOI211_X1 g_20_94 (.ZN (n_20_94), .A (n_24_92), .B (n_25_92), .C1 (n_29_90), .C2 (n_34_90) );
AOI211_X1 g_21_92 (.ZN (n_21_92), .A (n_22_93), .B (n_27_93), .C1 (n_27_91), .C2 (n_33_88) );
AOI211_X1 g_19_93 (.ZN (n_19_93), .A (n_20_94), .B (n_26_91), .C1 (n_25_92), .C2 (n_31_89) );
AOI211_X1 g_17_94 (.ZN (n_17_94), .A (n_21_92), .B (n_24_92), .C1 (n_27_93), .C2 (n_29_90) );
AOI211_X1 g_15_95 (.ZN (n_15_95), .A (n_19_93), .B (n_22_93), .C1 (n_26_91), .C2 (n_27_91) );
AOI211_X1 g_14_97 (.ZN (n_14_97), .A (n_17_94), .B (n_20_94), .C1 (n_24_92), .C2 (n_25_92) );
AOI211_X1 g_15_99 (.ZN (n_15_99), .A (n_15_95), .B (n_21_92), .C1 (n_22_93), .C2 (n_27_93) );
AOI211_X1 g_16_97 (.ZN (n_16_97), .A (n_14_97), .B (n_19_93), .C1 (n_20_94), .C2 (n_26_91) );
AOI211_X1 g_18_96 (.ZN (n_18_96), .A (n_15_99), .B (n_17_94), .C1 (n_21_92), .C2 (n_24_92) );
AOI211_X1 g_20_95 (.ZN (n_20_95), .A (n_16_97), .B (n_15_95), .C1 (n_19_93), .C2 (n_22_93) );
AOI211_X1 g_22_94 (.ZN (n_22_94), .A (n_18_96), .B (n_14_97), .C1 (n_17_94), .C2 (n_20_94) );
AOI211_X1 g_24_93 (.ZN (n_24_93), .A (n_20_95), .B (n_15_99), .C1 (n_15_95), .C2 (n_21_92) );
AOI211_X1 g_22_92 (.ZN (n_22_92), .A (n_22_94), .B (n_16_97), .C1 (n_14_97), .C2 (n_19_93) );
AOI211_X1 g_24_91 (.ZN (n_24_91), .A (n_24_93), .B (n_18_96), .C1 (n_15_99), .C2 (n_17_94) );
AOI211_X1 g_26_92 (.ZN (n_26_92), .A (n_22_92), .B (n_20_95), .C1 (n_16_97), .C2 (n_15_95) );
AOI211_X1 g_25_94 (.ZN (n_25_94), .A (n_24_91), .B (n_22_94), .C1 (n_18_96), .C2 (n_14_97) );
AOI211_X1 g_23_93 (.ZN (n_23_93), .A (n_26_92), .B (n_24_93), .C1 (n_20_95), .C2 (n_15_99) );
AOI211_X1 g_21_94 (.ZN (n_21_94), .A (n_25_94), .B (n_22_92), .C1 (n_22_94), .C2 (n_16_97) );
AOI211_X1 g_19_95 (.ZN (n_19_95), .A (n_23_93), .B (n_24_91), .C1 (n_24_93), .C2 (n_18_96) );
AOI211_X1 g_17_96 (.ZN (n_17_96), .A (n_21_94), .B (n_26_92), .C1 (n_22_92), .C2 (n_20_95) );
AOI211_X1 g_15_97 (.ZN (n_15_97), .A (n_19_95), .B (n_25_94), .C1 (n_24_91), .C2 (n_22_94) );
AOI211_X1 g_14_99 (.ZN (n_14_99), .A (n_17_96), .B (n_23_93), .C1 (n_26_92), .C2 (n_24_93) );
AOI211_X1 g_16_98 (.ZN (n_16_98), .A (n_15_97), .B (n_21_94), .C1 (n_25_94), .C2 (n_22_92) );
AOI211_X1 g_17_100 (.ZN (n_17_100), .A (n_14_99), .B (n_19_95), .C1 (n_23_93), .C2 (n_24_91) );
AOI211_X1 g_18_98 (.ZN (n_18_98), .A (n_16_98), .B (n_17_96), .C1 (n_21_94), .C2 (n_26_92) );
AOI211_X1 g_20_97 (.ZN (n_20_97), .A (n_17_100), .B (n_15_97), .C1 (n_19_95), .C2 (n_25_94) );
AOI211_X1 g_21_95 (.ZN (n_21_95), .A (n_18_98), .B (n_14_99), .C1 (n_17_96), .C2 (n_23_93) );
AOI211_X1 g_19_96 (.ZN (n_19_96), .A (n_20_97), .B (n_16_98), .C1 (n_15_97), .C2 (n_21_94) );
AOI211_X1 g_17_97 (.ZN (n_17_97), .A (n_21_95), .B (n_17_100), .C1 (n_14_99), .C2 (n_19_95) );
AOI211_X1 g_15_98 (.ZN (n_15_98), .A (n_19_96), .B (n_18_98), .C1 (n_16_98), .C2 (n_17_96) );
AOI211_X1 g_16_100 (.ZN (n_16_100), .A (n_17_97), .B (n_20_97), .C1 (n_17_100), .C2 (n_15_97) );
AOI211_X1 g_18_99 (.ZN (n_18_99), .A (n_15_98), .B (n_21_95), .C1 (n_18_98), .C2 (n_14_99) );
AOI211_X1 g_20_100 (.ZN (n_20_100), .A (n_16_100), .B (n_19_96), .C1 (n_20_97), .C2 (n_16_98) );
AOI211_X1 g_19_98 (.ZN (n_19_98), .A (n_18_99), .B (n_17_97), .C1 (n_21_95), .C2 (n_17_100) );
AOI211_X1 g_21_97 (.ZN (n_21_97), .A (n_20_100), .B (n_15_98), .C1 (n_19_96), .C2 (n_18_98) );
AOI211_X1 g_22_95 (.ZN (n_22_95), .A (n_19_98), .B (n_16_100), .C1 (n_17_97), .C2 (n_20_97) );
AOI211_X1 g_24_94 (.ZN (n_24_94), .A (n_21_97), .B (n_18_99), .C1 (n_15_98), .C2 (n_21_95) );
AOI211_X1 g_26_93 (.ZN (n_26_93), .A (n_22_95), .B (n_20_100), .C1 (n_16_100), .C2 (n_19_96) );
AOI211_X1 g_28_92 (.ZN (n_28_92), .A (n_24_94), .B (n_19_98), .C1 (n_18_99), .C2 (n_17_97) );
AOI211_X1 g_30_91 (.ZN (n_30_91), .A (n_26_93), .B (n_21_97), .C1 (n_20_100), .C2 (n_15_98) );
AOI211_X1 g_32_90 (.ZN (n_32_90), .A (n_28_92), .B (n_22_95), .C1 (n_19_98), .C2 (n_16_100) );
AOI211_X1 g_34_89 (.ZN (n_34_89), .A (n_30_91), .B (n_24_94), .C1 (n_21_97), .C2 (n_18_99) );
AOI211_X1 g_36_88 (.ZN (n_36_88), .A (n_32_90), .B (n_26_93), .C1 (n_22_95), .C2 (n_20_100) );
AOI211_X1 g_38_87 (.ZN (n_38_87), .A (n_34_89), .B (n_28_92), .C1 (n_24_94), .C2 (n_19_98) );
AOI211_X1 g_40_86 (.ZN (n_40_86), .A (n_36_88), .B (n_30_91), .C1 (n_26_93), .C2 (n_21_97) );
AOI211_X1 g_42_85 (.ZN (n_42_85), .A (n_38_87), .B (n_32_90), .C1 (n_28_92), .C2 (n_22_95) );
AOI211_X1 g_44_84 (.ZN (n_44_84), .A (n_40_86), .B (n_34_89), .C1 (n_30_91), .C2 (n_24_94) );
AOI211_X1 g_46_83 (.ZN (n_46_83), .A (n_42_85), .B (n_36_88), .C1 (n_32_90), .C2 (n_26_93) );
AOI211_X1 g_48_82 (.ZN (n_48_82), .A (n_44_84), .B (n_38_87), .C1 (n_34_89), .C2 (n_28_92) );
AOI211_X1 g_50_81 (.ZN (n_50_81), .A (n_46_83), .B (n_40_86), .C1 (n_36_88), .C2 (n_30_91) );
AOI211_X1 g_49_83 (.ZN (n_49_83), .A (n_48_82), .B (n_42_85), .C1 (n_38_87), .C2 (n_32_90) );
AOI211_X1 g_51_82 (.ZN (n_51_82), .A (n_50_81), .B (n_44_84), .C1 (n_40_86), .C2 (n_34_89) );
AOI211_X1 g_53_81 (.ZN (n_53_81), .A (n_49_83), .B (n_46_83), .C1 (n_42_85), .C2 (n_36_88) );
AOI211_X1 g_55_80 (.ZN (n_55_80), .A (n_51_82), .B (n_48_82), .C1 (n_44_84), .C2 (n_38_87) );
AOI211_X1 g_57_79 (.ZN (n_57_79), .A (n_53_81), .B (n_50_81), .C1 (n_46_83), .C2 (n_40_86) );
AOI211_X1 g_59_78 (.ZN (n_59_78), .A (n_55_80), .B (n_49_83), .C1 (n_48_82), .C2 (n_42_85) );
AOI211_X1 g_58_80 (.ZN (n_58_80), .A (n_57_79), .B (n_51_82), .C1 (n_50_81), .C2 (n_44_84) );
AOI211_X1 g_57_78 (.ZN (n_57_78), .A (n_59_78), .B (n_53_81), .C1 (n_49_83), .C2 (n_46_83) );
AOI211_X1 g_59_77 (.ZN (n_59_77), .A (n_58_80), .B (n_55_80), .C1 (n_51_82), .C2 (n_48_82) );
AOI211_X1 g_61_76 (.ZN (n_61_76), .A (n_57_78), .B (n_57_79), .C1 (n_53_81), .C2 (n_50_81) );
AOI211_X1 g_63_75 (.ZN (n_63_75), .A (n_59_77), .B (n_59_78), .C1 (n_55_80), .C2 (n_49_83) );
AOI211_X1 g_64_77 (.ZN (n_64_77), .A (n_61_76), .B (n_58_80), .C1 (n_57_79), .C2 (n_51_82) );
AOI211_X1 g_62_78 (.ZN (n_62_78), .A (n_63_75), .B (n_57_78), .C1 (n_59_78), .C2 (n_53_81) );
AOI211_X1 g_60_79 (.ZN (n_60_79), .A (n_64_77), .B (n_59_77), .C1 (n_58_80), .C2 (n_55_80) );
AOI211_X1 g_59_81 (.ZN (n_59_81), .A (n_62_78), .B (n_61_76), .C1 (n_57_78), .C2 (n_57_79) );
AOI211_X1 g_58_79 (.ZN (n_58_79), .A (n_60_79), .B (n_63_75), .C1 (n_59_77), .C2 (n_59_78) );
AOI211_X1 g_60_78 (.ZN (n_60_78), .A (n_59_81), .B (n_64_77), .C1 (n_61_76), .C2 (n_58_80) );
AOI211_X1 g_62_77 (.ZN (n_62_77), .A (n_58_79), .B (n_62_78), .C1 (n_63_75), .C2 (n_57_78) );
AOI211_X1 g_64_76 (.ZN (n_64_76), .A (n_60_78), .B (n_60_79), .C1 (n_64_77), .C2 (n_59_77) );
AOI211_X1 g_66_75 (.ZN (n_66_75), .A (n_62_77), .B (n_59_81), .C1 (n_62_78), .C2 (n_61_76) );
AOI211_X1 g_68_74 (.ZN (n_68_74), .A (n_64_76), .B (n_58_79), .C1 (n_60_79), .C2 (n_63_75) );
AOI211_X1 g_70_73 (.ZN (n_70_73), .A (n_66_75), .B (n_60_78), .C1 (n_59_81), .C2 (n_64_77) );
AOI211_X1 g_69_75 (.ZN (n_69_75), .A (n_68_74), .B (n_62_77), .C1 (n_58_79), .C2 (n_62_78) );
AOI211_X1 g_71_74 (.ZN (n_71_74), .A (n_70_73), .B (n_64_76), .C1 (n_60_78), .C2 (n_60_79) );
AOI211_X1 g_70_76 (.ZN (n_70_76), .A (n_69_75), .B (n_66_75), .C1 (n_62_77), .C2 (n_59_81) );
AOI211_X1 g_68_75 (.ZN (n_68_75), .A (n_71_74), .B (n_68_74), .C1 (n_64_76), .C2 (n_58_79) );
AOI211_X1 g_70_74 (.ZN (n_70_74), .A (n_70_76), .B (n_70_73), .C1 (n_66_75), .C2 (n_60_78) );
AOI211_X1 g_72_73 (.ZN (n_72_73), .A (n_68_75), .B (n_69_75), .C1 (n_68_74), .C2 (n_62_77) );
AOI211_X1 g_74_72 (.ZN (n_74_72), .A (n_70_74), .B (n_71_74), .C1 (n_70_73), .C2 (n_64_76) );
AOI211_X1 g_76_71 (.ZN (n_76_71), .A (n_72_73), .B (n_70_76), .C1 (n_69_75), .C2 (n_66_75) );
AOI211_X1 g_78_70 (.ZN (n_78_70), .A (n_74_72), .B (n_68_75), .C1 (n_71_74), .C2 (n_68_74) );
AOI211_X1 g_80_69 (.ZN (n_80_69), .A (n_76_71), .B (n_70_74), .C1 (n_70_76), .C2 (n_70_73) );
AOI211_X1 g_82_68 (.ZN (n_82_68), .A (n_78_70), .B (n_72_73), .C1 (n_68_75), .C2 (n_69_75) );
AOI211_X1 g_84_67 (.ZN (n_84_67), .A (n_80_69), .B (n_74_72), .C1 (n_70_74), .C2 (n_71_74) );
AOI211_X1 g_86_66 (.ZN (n_86_66), .A (n_82_68), .B (n_76_71), .C1 (n_72_73), .C2 (n_70_76) );
AOI211_X1 g_88_67 (.ZN (n_88_67), .A (n_84_67), .B (n_78_70), .C1 (n_74_72), .C2 (n_68_75) );
AOI211_X1 g_90_68 (.ZN (n_90_68), .A (n_86_66), .B (n_80_69), .C1 (n_76_71), .C2 (n_70_74) );
AOI211_X1 g_92_69 (.ZN (n_92_69), .A (n_88_67), .B (n_82_68), .C1 (n_78_70), .C2 (n_72_73) );
AOI211_X1 g_91_67 (.ZN (n_91_67), .A (n_90_68), .B (n_84_67), .C1 (n_80_69), .C2 (n_74_72) );
AOI211_X1 g_90_65 (.ZN (n_90_65), .A (n_92_69), .B (n_86_66), .C1 (n_82_68), .C2 (n_76_71) );
AOI211_X1 g_92_66 (.ZN (n_92_66), .A (n_91_67), .B (n_88_67), .C1 (n_84_67), .C2 (n_78_70) );
AOI211_X1 g_93_68 (.ZN (n_93_68), .A (n_90_65), .B (n_90_68), .C1 (n_86_66), .C2 (n_80_69) );
AOI211_X1 g_95_69 (.ZN (n_95_69), .A (n_92_66), .B (n_92_69), .C1 (n_88_67), .C2 (n_82_68) );
AOI211_X1 g_96_71 (.ZN (n_96_71), .A (n_93_68), .B (n_91_67), .C1 (n_90_68), .C2 (n_84_67) );
AOI211_X1 g_94_70 (.ZN (n_94_70), .A (n_95_69), .B (n_90_65), .C1 (n_92_69), .C2 (n_86_66) );
AOI211_X1 g_93_72 (.ZN (n_93_72), .A (n_96_71), .B (n_92_66), .C1 (n_91_67), .C2 (n_88_67) );
AOI211_X1 g_92_70 (.ZN (n_92_70), .A (n_94_70), .B (n_93_68), .C1 (n_90_65), .C2 (n_90_68) );
AOI211_X1 g_94_71 (.ZN (n_94_71), .A (n_93_72), .B (n_95_69), .C1 (n_92_66), .C2 (n_92_69) );
AOI211_X1 g_93_69 (.ZN (n_93_69), .A (n_92_70), .B (n_96_71), .C1 (n_93_68), .C2 (n_91_67) );
AOI211_X1 g_91_68 (.ZN (n_91_68), .A (n_94_71), .B (n_94_70), .C1 (n_95_69), .C2 (n_90_65) );
AOI211_X1 g_89_67 (.ZN (n_89_67), .A (n_93_69), .B (n_93_72), .C1 (n_96_71), .C2 (n_92_66) );
AOI211_X1 g_87_66 (.ZN (n_87_66), .A (n_91_68), .B (n_92_70), .C1 (n_94_70), .C2 (n_93_68) );
AOI211_X1 g_85_67 (.ZN (n_85_67), .A (n_89_67), .B (n_94_71), .C1 (n_93_72), .C2 (n_95_69) );
AOI211_X1 g_83_68 (.ZN (n_83_68), .A (n_87_66), .B (n_93_69), .C1 (n_92_70), .C2 (n_96_71) );
AOI211_X1 g_81_69 (.ZN (n_81_69), .A (n_85_67), .B (n_91_68), .C1 (n_94_71), .C2 (n_94_70) );
AOI211_X1 g_79_70 (.ZN (n_79_70), .A (n_83_68), .B (n_89_67), .C1 (n_93_69), .C2 (n_93_72) );
AOI211_X1 g_77_71 (.ZN (n_77_71), .A (n_81_69), .B (n_87_66), .C1 (n_91_68), .C2 (n_92_70) );
AOI211_X1 g_75_72 (.ZN (n_75_72), .A (n_79_70), .B (n_85_67), .C1 (n_89_67), .C2 (n_94_71) );
AOI211_X1 g_74_74 (.ZN (n_74_74), .A (n_77_71), .B (n_83_68), .C1 (n_87_66), .C2 (n_93_69) );
AOI211_X1 g_73_72 (.ZN (n_73_72), .A (n_75_72), .B (n_81_69), .C1 (n_85_67), .C2 (n_91_68) );
AOI211_X1 g_75_71 (.ZN (n_75_71), .A (n_74_74), .B (n_79_70), .C1 (n_83_68), .C2 (n_89_67) );
AOI211_X1 g_77_70 (.ZN (n_77_70), .A (n_73_72), .B (n_77_71), .C1 (n_81_69), .C2 (n_87_66) );
AOI211_X1 g_79_69 (.ZN (n_79_69), .A (n_75_71), .B (n_75_72), .C1 (n_79_70), .C2 (n_85_67) );
AOI211_X1 g_81_68 (.ZN (n_81_68), .A (n_77_70), .B (n_74_74), .C1 (n_77_71), .C2 (n_83_68) );
AOI211_X1 g_83_67 (.ZN (n_83_67), .A (n_79_69), .B (n_73_72), .C1 (n_75_72), .C2 (n_81_69) );
AOI211_X1 g_85_68 (.ZN (n_85_68), .A (n_81_68), .B (n_75_71), .C1 (n_74_74), .C2 (n_79_70) );
AOI211_X1 g_83_69 (.ZN (n_83_69), .A (n_83_67), .B (n_77_70), .C1 (n_73_72), .C2 (n_77_71) );
AOI211_X1 g_81_70 (.ZN (n_81_70), .A (n_85_68), .B (n_79_69), .C1 (n_75_71), .C2 (n_75_72) );
AOI211_X1 g_79_71 (.ZN (n_79_71), .A (n_83_69), .B (n_81_68), .C1 (n_77_70), .C2 (n_74_74) );
AOI211_X1 g_77_72 (.ZN (n_77_72), .A (n_81_70), .B (n_83_67), .C1 (n_79_69), .C2 (n_73_72) );
AOI211_X1 g_75_73 (.ZN (n_75_73), .A (n_79_71), .B (n_85_68), .C1 (n_81_68), .C2 (n_75_71) );
AOI211_X1 g_73_74 (.ZN (n_73_74), .A (n_77_72), .B (n_83_69), .C1 (n_83_67), .C2 (n_77_70) );
AOI211_X1 g_71_73 (.ZN (n_71_73), .A (n_75_73), .B (n_81_70), .C1 (n_85_68), .C2 (n_79_69) );
AOI211_X1 g_69_74 (.ZN (n_69_74), .A (n_73_74), .B (n_79_71), .C1 (n_83_69), .C2 (n_81_68) );
AOI211_X1 g_67_75 (.ZN (n_67_75), .A (n_71_73), .B (n_77_72), .C1 (n_81_70), .C2 (n_83_67) );
AOI211_X1 g_65_76 (.ZN (n_65_76), .A (n_69_74), .B (n_75_73), .C1 (n_79_71), .C2 (n_85_68) );
AOI211_X1 g_63_77 (.ZN (n_63_77), .A (n_67_75), .B (n_73_74), .C1 (n_77_72), .C2 (n_83_69) );
AOI211_X1 g_61_78 (.ZN (n_61_78), .A (n_65_76), .B (n_71_73), .C1 (n_75_73), .C2 (n_81_70) );
AOI211_X1 g_59_79 (.ZN (n_59_79), .A (n_63_77), .B (n_69_74), .C1 (n_73_74), .C2 (n_79_71) );
AOI211_X1 g_57_80 (.ZN (n_57_80), .A (n_61_78), .B (n_67_75), .C1 (n_71_73), .C2 (n_77_72) );
AOI211_X1 g_55_79 (.ZN (n_55_79), .A (n_59_79), .B (n_65_76), .C1 (n_69_74), .C2 (n_75_73) );
AOI211_X1 g_53_80 (.ZN (n_53_80), .A (n_57_80), .B (n_63_77), .C1 (n_67_75), .C2 (n_73_74) );
AOI211_X1 g_51_81 (.ZN (n_51_81), .A (n_55_79), .B (n_61_78), .C1 (n_65_76), .C2 (n_71_73) );
AOI211_X1 g_49_82 (.ZN (n_49_82), .A (n_53_80), .B (n_59_79), .C1 (n_63_77), .C2 (n_69_74) );
AOI211_X1 g_47_83 (.ZN (n_47_83), .A (n_51_81), .B (n_57_80), .C1 (n_61_78), .C2 (n_67_75) );
AOI211_X1 g_46_85 (.ZN (n_46_85), .A (n_49_82), .B (n_55_79), .C1 (n_59_79), .C2 (n_65_76) );
AOI211_X1 g_48_84 (.ZN (n_48_84), .A (n_47_83), .B (n_53_80), .C1 (n_57_80), .C2 (n_63_77) );
AOI211_X1 g_50_83 (.ZN (n_50_83), .A (n_46_85), .B (n_51_81), .C1 (n_55_79), .C2 (n_61_78) );
AOI211_X1 g_52_82 (.ZN (n_52_82), .A (n_48_84), .B (n_49_82), .C1 (n_53_80), .C2 (n_59_79) );
AOI211_X1 g_54_81 (.ZN (n_54_81), .A (n_50_83), .B (n_47_83), .C1 (n_51_81), .C2 (n_57_80) );
AOI211_X1 g_56_80 (.ZN (n_56_80), .A (n_52_82), .B (n_46_85), .C1 (n_49_82), .C2 (n_55_79) );
AOI211_X1 g_55_82 (.ZN (n_55_82), .A (n_54_81), .B (n_48_84), .C1 (n_47_83), .C2 (n_53_80) );
AOI211_X1 g_57_81 (.ZN (n_57_81), .A (n_56_80), .B (n_50_83), .C1 (n_46_85), .C2 (n_51_81) );
AOI211_X1 g_59_80 (.ZN (n_59_80), .A (n_55_82), .B (n_52_82), .C1 (n_48_84), .C2 (n_49_82) );
AOI211_X1 g_61_79 (.ZN (n_61_79), .A (n_57_81), .B (n_54_81), .C1 (n_50_83), .C2 (n_47_83) );
AOI211_X1 g_63_78 (.ZN (n_63_78), .A (n_59_80), .B (n_56_80), .C1 (n_52_82), .C2 (n_46_85) );
AOI211_X1 g_65_77 (.ZN (n_65_77), .A (n_61_79), .B (n_55_82), .C1 (n_54_81), .C2 (n_48_84) );
AOI211_X1 g_67_76 (.ZN (n_67_76), .A (n_63_78), .B (n_57_81), .C1 (n_56_80), .C2 (n_50_83) );
AOI211_X1 g_66_78 (.ZN (n_66_78), .A (n_65_77), .B (n_59_80), .C1 (n_55_82), .C2 (n_52_82) );
AOI211_X1 g_68_77 (.ZN (n_68_77), .A (n_67_76), .B (n_61_79), .C1 (n_57_81), .C2 (n_54_81) );
AOI211_X1 g_67_79 (.ZN (n_67_79), .A (n_66_78), .B (n_63_78), .C1 (n_59_80), .C2 (n_56_80) );
AOI211_X1 g_66_77 (.ZN (n_66_77), .A (n_68_77), .B (n_65_77), .C1 (n_61_79), .C2 (n_55_82) );
AOI211_X1 g_68_76 (.ZN (n_68_76), .A (n_67_79), .B (n_67_76), .C1 (n_63_78), .C2 (n_57_81) );
AOI211_X1 g_70_75 (.ZN (n_70_75), .A (n_66_77), .B (n_66_78), .C1 (n_65_77), .C2 (n_59_80) );
AOI211_X1 g_72_74 (.ZN (n_72_74), .A (n_68_76), .B (n_68_77), .C1 (n_67_76), .C2 (n_61_79) );
AOI211_X1 g_74_73 (.ZN (n_74_73), .A (n_70_75), .B (n_67_79), .C1 (n_66_78), .C2 (n_63_78) );
AOI211_X1 g_76_72 (.ZN (n_76_72), .A (n_72_74), .B (n_66_77), .C1 (n_68_77), .C2 (n_65_77) );
AOI211_X1 g_78_71 (.ZN (n_78_71), .A (n_74_73), .B (n_68_76), .C1 (n_67_79), .C2 (n_67_76) );
AOI211_X1 g_80_70 (.ZN (n_80_70), .A (n_76_72), .B (n_70_75), .C1 (n_66_77), .C2 (n_66_78) );
AOI211_X1 g_82_69 (.ZN (n_82_69), .A (n_78_71), .B (n_72_74), .C1 (n_68_76), .C2 (n_68_77) );
AOI211_X1 g_84_68 (.ZN (n_84_68), .A (n_80_70), .B (n_74_73), .C1 (n_70_75), .C2 (n_67_79) );
AOI211_X1 g_86_67 (.ZN (n_86_67), .A (n_82_69), .B (n_76_72), .C1 (n_72_74), .C2 (n_66_77) );
AOI211_X1 g_88_66 (.ZN (n_88_66), .A (n_84_68), .B (n_78_71), .C1 (n_74_73), .C2 (n_68_76) );
AOI211_X1 g_87_68 (.ZN (n_87_68), .A (n_86_67), .B (n_80_70), .C1 (n_76_72), .C2 (n_70_75) );
AOI211_X1 g_85_69 (.ZN (n_85_69), .A (n_88_66), .B (n_82_69), .C1 (n_78_71), .C2 (n_72_74) );
AOI211_X1 g_83_70 (.ZN (n_83_70), .A (n_87_68), .B (n_84_68), .C1 (n_80_70), .C2 (n_74_73) );
AOI211_X1 g_81_71 (.ZN (n_81_71), .A (n_85_69), .B (n_86_67), .C1 (n_82_69), .C2 (n_76_72) );
AOI211_X1 g_79_72 (.ZN (n_79_72), .A (n_83_70), .B (n_88_66), .C1 (n_84_68), .C2 (n_78_71) );
AOI211_X1 g_77_73 (.ZN (n_77_73), .A (n_81_71), .B (n_87_68), .C1 (n_86_67), .C2 (n_80_70) );
AOI211_X1 g_75_74 (.ZN (n_75_74), .A (n_79_72), .B (n_85_69), .C1 (n_88_66), .C2 (n_82_69) );
AOI211_X1 g_73_75 (.ZN (n_73_75), .A (n_77_73), .B (n_83_70), .C1 (n_87_68), .C2 (n_84_68) );
AOI211_X1 g_71_76 (.ZN (n_71_76), .A (n_75_74), .B (n_81_71), .C1 (n_85_69), .C2 (n_86_67) );
AOI211_X1 g_69_77 (.ZN (n_69_77), .A (n_73_75), .B (n_79_72), .C1 (n_83_70), .C2 (n_88_66) );
AOI211_X1 g_67_78 (.ZN (n_67_78), .A (n_71_76), .B (n_77_73), .C1 (n_81_71), .C2 (n_87_68) );
AOI211_X1 g_65_79 (.ZN (n_65_79), .A (n_69_77), .B (n_75_74), .C1 (n_79_72), .C2 (n_85_69) );
AOI211_X1 g_63_80 (.ZN (n_63_80), .A (n_67_78), .B (n_73_75), .C1 (n_77_73), .C2 (n_83_70) );
AOI211_X1 g_64_78 (.ZN (n_64_78), .A (n_65_79), .B (n_71_76), .C1 (n_75_74), .C2 (n_81_71) );
AOI211_X1 g_62_79 (.ZN (n_62_79), .A (n_63_80), .B (n_69_77), .C1 (n_73_75), .C2 (n_79_72) );
AOI211_X1 g_60_80 (.ZN (n_60_80), .A (n_64_78), .B (n_67_78), .C1 (n_71_76), .C2 (n_77_73) );
AOI211_X1 g_58_81 (.ZN (n_58_81), .A (n_62_79), .B (n_65_79), .C1 (n_69_77), .C2 (n_75_74) );
AOI211_X1 g_56_82 (.ZN (n_56_82), .A (n_60_80), .B (n_63_80), .C1 (n_67_78), .C2 (n_73_75) );
AOI211_X1 g_54_83 (.ZN (n_54_83), .A (n_58_81), .B (n_64_78), .C1 (n_65_79), .C2 (n_71_76) );
AOI211_X1 g_55_81 (.ZN (n_55_81), .A (n_56_82), .B (n_62_79), .C1 (n_63_80), .C2 (n_69_77) );
AOI211_X1 g_53_82 (.ZN (n_53_82), .A (n_54_83), .B (n_60_80), .C1 (n_64_78), .C2 (n_67_78) );
AOI211_X1 g_51_83 (.ZN (n_51_83), .A (n_55_81), .B (n_58_81), .C1 (n_62_79), .C2 (n_65_79) );
AOI211_X1 g_49_84 (.ZN (n_49_84), .A (n_53_82), .B (n_56_82), .C1 (n_60_80), .C2 (n_63_80) );
AOI211_X1 g_47_85 (.ZN (n_47_85), .A (n_51_83), .B (n_54_83), .C1 (n_58_81), .C2 (n_64_78) );
AOI211_X1 g_45_86 (.ZN (n_45_86), .A (n_49_84), .B (n_55_81), .C1 (n_56_82), .C2 (n_62_79) );
AOI211_X1 g_43_85 (.ZN (n_43_85), .A (n_47_85), .B (n_53_82), .C1 (n_54_83), .C2 (n_60_80) );
AOI211_X1 g_41_86 (.ZN (n_41_86), .A (n_45_86), .B (n_51_83), .C1 (n_55_81), .C2 (n_58_81) );
AOI211_X1 g_39_87 (.ZN (n_39_87), .A (n_43_85), .B (n_49_84), .C1 (n_53_82), .C2 (n_56_82) );
AOI211_X1 g_37_88 (.ZN (n_37_88), .A (n_41_86), .B (n_47_85), .C1 (n_51_83), .C2 (n_54_83) );
AOI211_X1 g_35_89 (.ZN (n_35_89), .A (n_39_87), .B (n_45_86), .C1 (n_49_84), .C2 (n_55_81) );
AOI211_X1 g_33_90 (.ZN (n_33_90), .A (n_37_88), .B (n_43_85), .C1 (n_47_85), .C2 (n_53_82) );
AOI211_X1 g_31_91 (.ZN (n_31_91), .A (n_35_89), .B (n_41_86), .C1 (n_45_86), .C2 (n_51_83) );
AOI211_X1 g_33_92 (.ZN (n_33_92), .A (n_33_90), .B (n_39_87), .C1 (n_43_85), .C2 (n_49_84) );
AOI211_X1 g_35_91 (.ZN (n_35_91), .A (n_31_91), .B (n_37_88), .C1 (n_41_86), .C2 (n_47_85) );
AOI211_X1 g_37_90 (.ZN (n_37_90), .A (n_33_92), .B (n_35_89), .C1 (n_39_87), .C2 (n_45_86) );
AOI211_X1 g_39_89 (.ZN (n_39_89), .A (n_35_91), .B (n_33_90), .C1 (n_37_88), .C2 (n_43_85) );
AOI211_X1 g_41_88 (.ZN (n_41_88), .A (n_37_90), .B (n_31_91), .C1 (n_35_89), .C2 (n_41_86) );
AOI211_X1 g_43_87 (.ZN (n_43_87), .A (n_39_89), .B (n_33_92), .C1 (n_33_90), .C2 (n_39_87) );
AOI211_X1 g_42_89 (.ZN (n_42_89), .A (n_41_88), .B (n_35_91), .C1 (n_31_91), .C2 (n_37_88) );
AOI211_X1 g_41_87 (.ZN (n_41_87), .A (n_43_87), .B (n_37_90), .C1 (n_33_92), .C2 (n_35_89) );
AOI211_X1 g_43_86 (.ZN (n_43_86), .A (n_42_89), .B (n_39_89), .C1 (n_35_91), .C2 (n_33_90) );
AOI211_X1 g_45_85 (.ZN (n_45_85), .A (n_41_87), .B (n_41_88), .C1 (n_37_90), .C2 (n_31_91) );
AOI211_X1 g_47_84 (.ZN (n_47_84), .A (n_43_86), .B (n_43_87), .C1 (n_39_89), .C2 (n_33_92) );
AOI211_X1 g_46_86 (.ZN (n_46_86), .A (n_45_85), .B (n_42_89), .C1 (n_41_88), .C2 (n_35_91) );
AOI211_X1 g_48_85 (.ZN (n_48_85), .A (n_47_84), .B (n_41_87), .C1 (n_43_87), .C2 (n_37_90) );
AOI211_X1 g_50_84 (.ZN (n_50_84), .A (n_46_86), .B (n_43_86), .C1 (n_42_89), .C2 (n_39_89) );
AOI211_X1 g_52_83 (.ZN (n_52_83), .A (n_48_85), .B (n_45_85), .C1 (n_41_87), .C2 (n_41_88) );
AOI211_X1 g_54_82 (.ZN (n_54_82), .A (n_50_84), .B (n_47_84), .C1 (n_43_86), .C2 (n_43_87) );
AOI211_X1 g_56_81 (.ZN (n_56_81), .A (n_52_83), .B (n_46_86), .C1 (n_45_85), .C2 (n_42_89) );
AOI211_X1 g_55_83 (.ZN (n_55_83), .A (n_54_82), .B (n_48_85), .C1 (n_47_84), .C2 (n_41_87) );
AOI211_X1 g_57_82 (.ZN (n_57_82), .A (n_56_81), .B (n_50_84), .C1 (n_46_86), .C2 (n_43_86) );
AOI211_X1 g_56_84 (.ZN (n_56_84), .A (n_55_83), .B (n_52_83), .C1 (n_48_85), .C2 (n_45_85) );
AOI211_X1 g_58_83 (.ZN (n_58_83), .A (n_57_82), .B (n_54_82), .C1 (n_50_84), .C2 (n_47_84) );
AOI211_X1 g_60_82 (.ZN (n_60_82), .A (n_56_84), .B (n_56_81), .C1 (n_52_83), .C2 (n_46_86) );
AOI211_X1 g_61_80 (.ZN (n_61_80), .A (n_58_83), .B (n_55_83), .C1 (n_54_82), .C2 (n_48_85) );
AOI211_X1 g_63_79 (.ZN (n_63_79), .A (n_60_82), .B (n_57_82), .C1 (n_56_81), .C2 (n_50_84) );
AOI211_X1 g_65_78 (.ZN (n_65_78), .A (n_61_80), .B (n_56_84), .C1 (n_55_83), .C2 (n_52_83) );
AOI211_X1 g_67_77 (.ZN (n_67_77), .A (n_63_79), .B (n_58_83), .C1 (n_57_82), .C2 (n_54_82) );
AOI211_X1 g_69_76 (.ZN (n_69_76), .A (n_65_78), .B (n_60_82), .C1 (n_56_84), .C2 (n_56_81) );
AOI211_X1 g_71_75 (.ZN (n_71_75), .A (n_67_77), .B (n_61_80), .C1 (n_58_83), .C2 (n_55_83) );
AOI211_X1 g_70_77 (.ZN (n_70_77), .A (n_69_76), .B (n_63_79), .C1 (n_60_82), .C2 (n_57_82) );
AOI211_X1 g_72_76 (.ZN (n_72_76), .A (n_71_75), .B (n_65_78), .C1 (n_61_80), .C2 (n_56_84) );
AOI211_X1 g_74_75 (.ZN (n_74_75), .A (n_70_77), .B (n_67_77), .C1 (n_63_79), .C2 (n_58_83) );
AOI211_X1 g_76_74 (.ZN (n_76_74), .A (n_72_76), .B (n_69_76), .C1 (n_65_78), .C2 (n_60_82) );
AOI211_X1 g_78_73 (.ZN (n_78_73), .A (n_74_75), .B (n_71_75), .C1 (n_67_77), .C2 (n_61_80) );
AOI211_X1 g_80_72 (.ZN (n_80_72), .A (n_76_74), .B (n_70_77), .C1 (n_69_76), .C2 (n_63_79) );
AOI211_X1 g_82_71 (.ZN (n_82_71), .A (n_78_73), .B (n_72_76), .C1 (n_71_75), .C2 (n_65_78) );
AOI211_X1 g_84_70 (.ZN (n_84_70), .A (n_80_72), .B (n_74_75), .C1 (n_70_77), .C2 (n_67_77) );
AOI211_X1 g_86_69 (.ZN (n_86_69), .A (n_82_71), .B (n_76_74), .C1 (n_72_76), .C2 (n_69_76) );
AOI211_X1 g_88_68 (.ZN (n_88_68), .A (n_84_70), .B (n_78_73), .C1 (n_74_75), .C2 (n_71_75) );
AOI211_X1 g_90_67 (.ZN (n_90_67), .A (n_86_69), .B (n_80_72), .C1 (n_76_74), .C2 (n_70_77) );
AOI211_X1 g_92_68 (.ZN (n_92_68), .A (n_88_68), .B (n_82_71), .C1 (n_78_73), .C2 (n_72_76) );
AOI211_X1 g_90_69 (.ZN (n_90_69), .A (n_90_67), .B (n_84_70), .C1 (n_80_72), .C2 (n_74_75) );
AOI211_X1 g_88_70 (.ZN (n_88_70), .A (n_92_68), .B (n_86_69), .C1 (n_82_71), .C2 (n_76_74) );
AOI211_X1 g_89_68 (.ZN (n_89_68), .A (n_90_69), .B (n_88_68), .C1 (n_84_70), .C2 (n_78_73) );
AOI211_X1 g_87_69 (.ZN (n_87_69), .A (n_88_70), .B (n_90_67), .C1 (n_86_69), .C2 (n_80_72) );
AOI211_X1 g_86_71 (.ZN (n_86_71), .A (n_89_68), .B (n_92_68), .C1 (n_88_68), .C2 (n_82_71) );
AOI211_X1 g_84_72 (.ZN (n_84_72), .A (n_87_69), .B (n_90_69), .C1 (n_90_67), .C2 (n_84_70) );
AOI211_X1 g_85_70 (.ZN (n_85_70), .A (n_86_71), .B (n_88_70), .C1 (n_92_68), .C2 (n_86_69) );
AOI211_X1 g_86_68 (.ZN (n_86_68), .A (n_84_72), .B (n_89_68), .C1 (n_90_69), .C2 (n_88_68) );
AOI211_X1 g_84_69 (.ZN (n_84_69), .A (n_85_70), .B (n_87_69), .C1 (n_88_70), .C2 (n_90_67) );
AOI211_X1 g_82_70 (.ZN (n_82_70), .A (n_86_68), .B (n_86_71), .C1 (n_89_68), .C2 (n_92_68) );
AOI211_X1 g_80_71 (.ZN (n_80_71), .A (n_84_69), .B (n_84_72), .C1 (n_87_69), .C2 (n_90_69) );
AOI211_X1 g_78_72 (.ZN (n_78_72), .A (n_82_70), .B (n_85_70), .C1 (n_86_71), .C2 (n_88_70) );
AOI211_X1 g_76_73 (.ZN (n_76_73), .A (n_80_71), .B (n_86_68), .C1 (n_84_72), .C2 (n_89_68) );
AOI211_X1 g_75_75 (.ZN (n_75_75), .A (n_78_72), .B (n_84_69), .C1 (n_85_70), .C2 (n_87_69) );
AOI211_X1 g_77_74 (.ZN (n_77_74), .A (n_76_73), .B (n_82_70), .C1 (n_86_68), .C2 (n_86_71) );
AOI211_X1 g_79_73 (.ZN (n_79_73), .A (n_75_75), .B (n_80_71), .C1 (n_84_69), .C2 (n_84_72) );
AOI211_X1 g_81_72 (.ZN (n_81_72), .A (n_77_74), .B (n_78_72), .C1 (n_82_70), .C2 (n_85_70) );
AOI211_X1 g_83_71 (.ZN (n_83_71), .A (n_79_73), .B (n_76_73), .C1 (n_80_71), .C2 (n_86_68) );
AOI211_X1 g_82_73 (.ZN (n_82_73), .A (n_81_72), .B (n_75_75), .C1 (n_78_72), .C2 (n_84_69) );
AOI211_X1 g_80_74 (.ZN (n_80_74), .A (n_83_71), .B (n_77_74), .C1 (n_76_73), .C2 (n_82_70) );
AOI211_X1 g_78_75 (.ZN (n_78_75), .A (n_82_73), .B (n_79_73), .C1 (n_75_75), .C2 (n_80_71) );
AOI211_X1 g_76_76 (.ZN (n_76_76), .A (n_80_74), .B (n_81_72), .C1 (n_77_74), .C2 (n_78_72) );
AOI211_X1 g_74_77 (.ZN (n_74_77), .A (n_78_75), .B (n_83_71), .C1 (n_79_73), .C2 (n_76_73) );
AOI211_X1 g_72_78 (.ZN (n_72_78), .A (n_76_76), .B (n_82_73), .C1 (n_81_72), .C2 (n_75_75) );
AOI211_X1 g_73_76 (.ZN (n_73_76), .A (n_74_77), .B (n_80_74), .C1 (n_83_71), .C2 (n_77_74) );
AOI211_X1 g_71_77 (.ZN (n_71_77), .A (n_72_78), .B (n_78_75), .C1 (n_82_73), .C2 (n_79_73) );
AOI211_X1 g_72_75 (.ZN (n_72_75), .A (n_73_76), .B (n_76_76), .C1 (n_80_74), .C2 (n_81_72) );
AOI211_X1 g_73_77 (.ZN (n_73_77), .A (n_71_77), .B (n_74_77), .C1 (n_78_75), .C2 (n_83_71) );
AOI211_X1 g_75_76 (.ZN (n_75_76), .A (n_72_75), .B (n_72_78), .C1 (n_76_76), .C2 (n_82_73) );
AOI211_X1 g_77_75 (.ZN (n_77_75), .A (n_73_77), .B (n_73_76), .C1 (n_74_77), .C2 (n_80_74) );
AOI211_X1 g_79_74 (.ZN (n_79_74), .A (n_75_76), .B (n_71_77), .C1 (n_72_78), .C2 (n_78_75) );
AOI211_X1 g_81_73 (.ZN (n_81_73), .A (n_77_75), .B (n_72_75), .C1 (n_73_76), .C2 (n_76_76) );
AOI211_X1 g_83_72 (.ZN (n_83_72), .A (n_79_74), .B (n_73_77), .C1 (n_71_77), .C2 (n_74_77) );
AOI211_X1 g_85_71 (.ZN (n_85_71), .A (n_81_73), .B (n_75_76), .C1 (n_72_75), .C2 (n_72_78) );
AOI211_X1 g_87_70 (.ZN (n_87_70), .A (n_83_72), .B (n_77_75), .C1 (n_73_77), .C2 (n_73_76) );
AOI211_X1 g_89_69 (.ZN (n_89_69), .A (n_85_71), .B (n_79_74), .C1 (n_75_76), .C2 (n_71_77) );
AOI211_X1 g_91_70 (.ZN (n_91_70), .A (n_87_70), .B (n_81_73), .C1 (n_77_75), .C2 (n_72_75) );
AOI211_X1 g_93_71 (.ZN (n_93_71), .A (n_89_69), .B (n_83_72), .C1 (n_79_74), .C2 (n_73_77) );
AOI211_X1 g_95_72 (.ZN (n_95_72), .A (n_91_70), .B (n_85_71), .C1 (n_81_73), .C2 (n_75_76) );
AOI211_X1 g_97_73 (.ZN (n_97_73), .A (n_93_71), .B (n_87_70), .C1 (n_83_72), .C2 (n_77_75) );
AOI211_X1 g_96_75 (.ZN (n_96_75), .A (n_95_72), .B (n_89_69), .C1 (n_85_71), .C2 (n_79_74) );
AOI211_X1 g_94_74 (.ZN (n_94_74), .A (n_97_73), .B (n_91_70), .C1 (n_87_70), .C2 (n_81_73) );
AOI211_X1 g_92_73 (.ZN (n_92_73), .A (n_96_75), .B (n_93_71), .C1 (n_89_69), .C2 (n_83_72) );
AOI211_X1 g_94_72 (.ZN (n_94_72), .A (n_94_74), .B (n_95_72), .C1 (n_91_70), .C2 (n_85_71) );
AOI211_X1 g_93_70 (.ZN (n_93_70), .A (n_92_73), .B (n_97_73), .C1 (n_93_71), .C2 (n_87_70) );
AOI211_X1 g_91_69 (.ZN (n_91_69), .A (n_94_72), .B (n_96_75), .C1 (n_95_72), .C2 (n_89_69) );
AOI211_X1 g_89_70 (.ZN (n_89_70), .A (n_93_70), .B (n_94_74), .C1 (n_97_73), .C2 (n_91_70) );
AOI211_X1 g_91_71 (.ZN (n_91_71), .A (n_91_69), .B (n_92_73), .C1 (n_96_75), .C2 (n_93_71) );
AOI211_X1 g_89_72 (.ZN (n_89_72), .A (n_89_70), .B (n_94_72), .C1 (n_94_74), .C2 (n_95_72) );
AOI211_X1 g_90_70 (.ZN (n_90_70), .A (n_91_71), .B (n_93_70), .C1 (n_92_73), .C2 (n_97_73) );
AOI211_X1 g_88_69 (.ZN (n_88_69), .A (n_89_72), .B (n_91_69), .C1 (n_94_72), .C2 (n_96_75) );
AOI211_X1 g_87_71 (.ZN (n_87_71), .A (n_90_70), .B (n_89_70), .C1 (n_93_70), .C2 (n_94_74) );
AOI211_X1 g_85_72 (.ZN (n_85_72), .A (n_88_69), .B (n_91_71), .C1 (n_91_69), .C2 (n_92_73) );
AOI211_X1 g_86_70 (.ZN (n_86_70), .A (n_87_71), .B (n_89_72), .C1 (n_89_70), .C2 (n_94_72) );
AOI211_X1 g_84_71 (.ZN (n_84_71), .A (n_85_72), .B (n_90_70), .C1 (n_91_71), .C2 (n_93_70) );
AOI211_X1 g_82_72 (.ZN (n_82_72), .A (n_86_70), .B (n_88_69), .C1 (n_89_72), .C2 (n_91_69) );
AOI211_X1 g_80_73 (.ZN (n_80_73), .A (n_84_71), .B (n_87_71), .C1 (n_90_70), .C2 (n_89_70) );
AOI211_X1 g_78_74 (.ZN (n_78_74), .A (n_82_72), .B (n_85_72), .C1 (n_88_69), .C2 (n_91_71) );
AOI211_X1 g_76_75 (.ZN (n_76_75), .A (n_80_73), .B (n_86_70), .C1 (n_87_71), .C2 (n_89_72) );
AOI211_X1 g_74_76 (.ZN (n_74_76), .A (n_78_74), .B (n_84_71), .C1 (n_85_72), .C2 (n_90_70) );
AOI211_X1 g_72_77 (.ZN (n_72_77), .A (n_76_75), .B (n_82_72), .C1 (n_86_70), .C2 (n_88_69) );
AOI211_X1 g_70_78 (.ZN (n_70_78), .A (n_74_76), .B (n_80_73), .C1 (n_84_71), .C2 (n_87_71) );
AOI211_X1 g_68_79 (.ZN (n_68_79), .A (n_72_77), .B (n_78_74), .C1 (n_82_72), .C2 (n_85_72) );
AOI211_X1 g_66_80 (.ZN (n_66_80), .A (n_70_78), .B (n_76_75), .C1 (n_80_73), .C2 (n_86_70) );
AOI211_X1 g_64_79 (.ZN (n_64_79), .A (n_68_79), .B (n_74_76), .C1 (n_78_74), .C2 (n_84_71) );
AOI211_X1 g_62_80 (.ZN (n_62_80), .A (n_66_80), .B (n_72_77), .C1 (n_76_75), .C2 (n_82_72) );
AOI211_X1 g_60_81 (.ZN (n_60_81), .A (n_64_79), .B (n_70_78), .C1 (n_74_76), .C2 (n_80_73) );
AOI211_X1 g_58_82 (.ZN (n_58_82), .A (n_62_80), .B (n_68_79), .C1 (n_72_77), .C2 (n_78_74) );
AOI211_X1 g_56_83 (.ZN (n_56_83), .A (n_60_81), .B (n_66_80), .C1 (n_70_78), .C2 (n_76_75) );
AOI211_X1 g_54_84 (.ZN (n_54_84), .A (n_58_82), .B (n_64_79), .C1 (n_68_79), .C2 (n_74_76) );
AOI211_X1 g_52_85 (.ZN (n_52_85), .A (n_56_83), .B (n_62_80), .C1 (n_66_80), .C2 (n_72_77) );
AOI211_X1 g_53_83 (.ZN (n_53_83), .A (n_54_84), .B (n_60_81), .C1 (n_64_79), .C2 (n_70_78) );
AOI211_X1 g_51_84 (.ZN (n_51_84), .A (n_52_85), .B (n_58_82), .C1 (n_62_80), .C2 (n_68_79) );
AOI211_X1 g_49_85 (.ZN (n_49_85), .A (n_53_83), .B (n_56_83), .C1 (n_60_81), .C2 (n_66_80) );
AOI211_X1 g_47_86 (.ZN (n_47_86), .A (n_51_84), .B (n_54_84), .C1 (n_58_82), .C2 (n_64_79) );
AOI211_X1 g_45_87 (.ZN (n_45_87), .A (n_49_85), .B (n_52_85), .C1 (n_56_83), .C2 (n_62_80) );
AOI211_X1 g_43_88 (.ZN (n_43_88), .A (n_47_86), .B (n_53_83), .C1 (n_54_84), .C2 (n_60_81) );
AOI211_X1 g_44_86 (.ZN (n_44_86), .A (n_45_87), .B (n_51_84), .C1 (n_52_85), .C2 (n_58_82) );
AOI211_X1 g_42_87 (.ZN (n_42_87), .A (n_43_88), .B (n_49_85), .C1 (n_53_83), .C2 (n_56_83) );
AOI211_X1 g_40_88 (.ZN (n_40_88), .A (n_44_86), .B (n_47_86), .C1 (n_51_84), .C2 (n_54_84) );
AOI211_X1 g_38_89 (.ZN (n_38_89), .A (n_42_87), .B (n_45_87), .C1 (n_49_85), .C2 (n_52_85) );
AOI211_X1 g_36_90 (.ZN (n_36_90), .A (n_40_88), .B (n_43_88), .C1 (n_47_86), .C2 (n_53_83) );
AOI211_X1 g_34_91 (.ZN (n_34_91), .A (n_38_89), .B (n_44_86), .C1 (n_45_87), .C2 (n_51_84) );
AOI211_X1 g_33_89 (.ZN (n_33_89), .A (n_36_90), .B (n_42_87), .C1 (n_43_88), .C2 (n_49_85) );
AOI211_X1 g_31_90 (.ZN (n_31_90), .A (n_34_91), .B (n_40_88), .C1 (n_44_86), .C2 (n_47_86) );
AOI211_X1 g_29_91 (.ZN (n_29_91), .A (n_33_89), .B (n_38_89), .C1 (n_42_87), .C2 (n_45_87) );
AOI211_X1 g_27_92 (.ZN (n_27_92), .A (n_31_90), .B (n_36_90), .C1 (n_40_88), .C2 (n_43_88) );
AOI211_X1 g_25_93 (.ZN (n_25_93), .A (n_29_91), .B (n_34_91), .C1 (n_38_89), .C2 (n_44_86) );
AOI211_X1 g_23_94 (.ZN (n_23_94), .A (n_27_92), .B (n_33_89), .C1 (n_36_90), .C2 (n_42_87) );
AOI211_X1 g_22_96 (.ZN (n_22_96), .A (n_25_93), .B (n_31_90), .C1 (n_34_91), .C2 (n_40_88) );
AOI211_X1 g_23_98 (.ZN (n_23_98), .A (n_23_94), .B (n_29_91), .C1 (n_33_89), .C2 (n_38_89) );
AOI211_X1 g_24_100 (.ZN (n_24_100), .A (n_22_96), .B (n_27_92), .C1 (n_31_90), .C2 (n_36_90) );
AOI211_X1 g_22_99 (.ZN (n_22_99), .A (n_23_98), .B (n_25_93), .C1 (n_29_91), .C2 (n_34_91) );
AOI211_X1 g_20_98 (.ZN (n_20_98), .A (n_24_100), .B (n_23_94), .C1 (n_27_92), .C2 (n_33_89) );
AOI211_X1 g_18_97 (.ZN (n_18_97), .A (n_22_99), .B (n_22_96), .C1 (n_25_93), .C2 (n_31_90) );
AOI211_X1 g_16_96 (.ZN (n_16_96), .A (n_20_98), .B (n_23_98), .C1 (n_23_94), .C2 (n_29_91) );
AOI211_X1 g_18_95 (.ZN (n_18_95), .A (n_18_97), .B (n_24_100), .C1 (n_22_96), .C2 (n_27_92) );
AOI211_X1 g_20_96 (.ZN (n_20_96), .A (n_16_96), .B (n_22_99), .C1 (n_23_98), .C2 (n_25_93) );
AOI211_X1 g_21_98 (.ZN (n_21_98), .A (n_18_95), .B (n_20_98), .C1 (n_24_100), .C2 (n_23_94) );
AOI211_X1 g_19_97 (.ZN (n_19_97), .A (n_20_96), .B (n_18_97), .C1 (n_22_99), .C2 (n_22_96) );
AOI211_X1 g_17_98 (.ZN (n_17_98), .A (n_21_98), .B (n_16_96), .C1 (n_20_98), .C2 (n_23_98) );
AOI211_X1 g_19_99 (.ZN (n_19_99), .A (n_19_97), .B (n_18_95), .C1 (n_18_97), .C2 (n_24_100) );
AOI211_X1 g_21_100 (.ZN (n_21_100), .A (n_17_98), .B (n_20_96), .C1 (n_16_96), .C2 (n_22_99) );
AOI211_X1 g_22_98 (.ZN (n_22_98), .A (n_19_99), .B (n_21_98), .C1 (n_18_95), .C2 (n_20_98) );
AOI211_X1 g_21_96 (.ZN (n_21_96), .A (n_21_100), .B (n_19_97), .C1 (n_20_96), .C2 (n_18_97) );
AOI211_X1 g_23_95 (.ZN (n_23_95), .A (n_22_98), .B (n_17_98), .C1 (n_21_98), .C2 (n_16_96) );
AOI211_X1 g_22_97 (.ZN (n_22_97), .A (n_21_96), .B (n_19_99), .C1 (n_19_97), .C2 (n_18_95) );
AOI211_X1 g_24_96 (.ZN (n_24_96), .A (n_23_95), .B (n_21_100), .C1 (n_17_98), .C2 (n_20_96) );
AOI211_X1 g_26_95 (.ZN (n_26_95), .A (n_22_97), .B (n_22_98), .C1 (n_19_99), .C2 (n_21_98) );
AOI211_X1 g_28_94 (.ZN (n_28_94), .A (n_24_96), .B (n_21_96), .C1 (n_21_100), .C2 (n_19_97) );
AOI211_X1 g_30_93 (.ZN (n_30_93), .A (n_26_95), .B (n_23_95), .C1 (n_22_98), .C2 (n_17_98) );
AOI211_X1 g_32_92 (.ZN (n_32_92), .A (n_28_94), .B (n_22_97), .C1 (n_21_96), .C2 (n_19_99) );
AOI211_X1 g_34_93 (.ZN (n_34_93), .A (n_30_93), .B (n_24_96), .C1 (n_23_95), .C2 (n_21_100) );
AOI211_X1 g_33_91 (.ZN (n_33_91), .A (n_32_92), .B (n_26_95), .C1 (n_22_97), .C2 (n_22_98) );
AOI211_X1 g_35_90 (.ZN (n_35_90), .A (n_34_93), .B (n_28_94), .C1 (n_24_96), .C2 (n_21_96) );
AOI211_X1 g_37_89 (.ZN (n_37_89), .A (n_33_91), .B (n_30_93), .C1 (n_26_95), .C2 (n_23_95) );
AOI211_X1 g_39_88 (.ZN (n_39_88), .A (n_35_90), .B (n_32_92), .C1 (n_28_94), .C2 (n_22_97) );
AOI211_X1 g_40_90 (.ZN (n_40_90), .A (n_37_89), .B (n_34_93), .C1 (n_30_93), .C2 (n_24_96) );
AOI211_X1 g_38_91 (.ZN (n_38_91), .A (n_39_88), .B (n_33_91), .C1 (n_32_92), .C2 (n_26_95) );
AOI211_X1 g_36_92 (.ZN (n_36_92), .A (n_40_90), .B (n_35_90), .C1 (n_34_93), .C2 (n_28_94) );
AOI211_X1 g_35_94 (.ZN (n_35_94), .A (n_38_91), .B (n_37_89), .C1 (n_33_91), .C2 (n_30_93) );
AOI211_X1 g_34_92 (.ZN (n_34_92), .A (n_36_92), .B (n_39_88), .C1 (n_35_90), .C2 (n_32_92) );
AOI211_X1 g_32_91 (.ZN (n_32_91), .A (n_35_94), .B (n_40_90), .C1 (n_37_89), .C2 (n_34_93) );
AOI211_X1 g_30_92 (.ZN (n_30_92), .A (n_34_92), .B (n_38_91), .C1 (n_39_88), .C2 (n_33_91) );
AOI211_X1 g_28_93 (.ZN (n_28_93), .A (n_32_91), .B (n_36_92), .C1 (n_40_90), .C2 (n_35_90) );
AOI211_X1 g_26_94 (.ZN (n_26_94), .A (n_30_92), .B (n_35_94), .C1 (n_38_91), .C2 (n_37_89) );
AOI211_X1 g_24_95 (.ZN (n_24_95), .A (n_28_93), .B (n_34_92), .C1 (n_36_92), .C2 (n_39_88) );
AOI211_X1 g_23_97 (.ZN (n_23_97), .A (n_26_94), .B (n_32_91), .C1 (n_35_94), .C2 (n_40_90) );
AOI211_X1 g_25_96 (.ZN (n_25_96), .A (n_24_95), .B (n_30_92), .C1 (n_34_92), .C2 (n_38_91) );
AOI211_X1 g_27_95 (.ZN (n_27_95), .A (n_23_97), .B (n_28_93), .C1 (n_32_91), .C2 (n_36_92) );
AOI211_X1 g_29_94 (.ZN (n_29_94), .A (n_25_96), .B (n_26_94), .C1 (n_30_92), .C2 (n_35_94) );
AOI211_X1 g_31_93 (.ZN (n_31_93), .A (n_27_95), .B (n_24_95), .C1 (n_28_93), .C2 (n_34_92) );
AOI211_X1 g_33_94 (.ZN (n_33_94), .A (n_29_94), .B (n_23_97), .C1 (n_26_94), .C2 (n_32_91) );
AOI211_X1 g_35_93 (.ZN (n_35_93), .A (n_31_93), .B (n_25_96), .C1 (n_24_95), .C2 (n_30_92) );
AOI211_X1 g_36_91 (.ZN (n_36_91), .A (n_33_94), .B (n_27_95), .C1 (n_23_97), .C2 (n_28_93) );
AOI211_X1 g_38_90 (.ZN (n_38_90), .A (n_35_93), .B (n_29_94), .C1 (n_25_96), .C2 (n_26_94) );
AOI211_X1 g_40_89 (.ZN (n_40_89), .A (n_36_91), .B (n_31_93), .C1 (n_27_95), .C2 (n_24_95) );
AOI211_X1 g_42_88 (.ZN (n_42_88), .A (n_38_90), .B (n_33_94), .C1 (n_29_94), .C2 (n_23_97) );
AOI211_X1 g_44_87 (.ZN (n_44_87), .A (n_40_89), .B (n_35_93), .C1 (n_31_93), .C2 (n_25_96) );
AOI211_X1 g_43_89 (.ZN (n_43_89), .A (n_42_88), .B (n_36_91), .C1 (n_33_94), .C2 (n_27_95) );
AOI211_X1 g_45_88 (.ZN (n_45_88), .A (n_44_87), .B (n_38_90), .C1 (n_35_93), .C2 (n_29_94) );
AOI211_X1 g_47_87 (.ZN (n_47_87), .A (n_43_89), .B (n_40_89), .C1 (n_36_91), .C2 (n_31_93) );
AOI211_X1 g_49_86 (.ZN (n_49_86), .A (n_45_88), .B (n_42_88), .C1 (n_38_90), .C2 (n_33_94) );
AOI211_X1 g_51_85 (.ZN (n_51_85), .A (n_47_87), .B (n_44_87), .C1 (n_40_89), .C2 (n_35_93) );
AOI211_X1 g_53_84 (.ZN (n_53_84), .A (n_49_86), .B (n_43_89), .C1 (n_42_88), .C2 (n_36_91) );
AOI211_X1 g_55_85 (.ZN (n_55_85), .A (n_51_85), .B (n_45_88), .C1 (n_44_87), .C2 (n_38_90) );
AOI211_X1 g_57_84 (.ZN (n_57_84), .A (n_53_84), .B (n_47_87), .C1 (n_43_89), .C2 (n_40_89) );
AOI211_X1 g_59_83 (.ZN (n_59_83), .A (n_55_85), .B (n_49_86), .C1 (n_45_88), .C2 (n_42_88) );
AOI211_X1 g_61_82 (.ZN (n_61_82), .A (n_57_84), .B (n_51_85), .C1 (n_47_87), .C2 (n_44_87) );
AOI211_X1 g_63_81 (.ZN (n_63_81), .A (n_59_83), .B (n_53_84), .C1 (n_49_86), .C2 (n_43_89) );
AOI211_X1 g_65_80 (.ZN (n_65_80), .A (n_61_82), .B (n_55_85), .C1 (n_51_85), .C2 (n_45_88) );
AOI211_X1 g_64_82 (.ZN (n_64_82), .A (n_63_81), .B (n_57_84), .C1 (n_53_84), .C2 (n_47_87) );
AOI211_X1 g_62_81 (.ZN (n_62_81), .A (n_65_80), .B (n_59_83), .C1 (n_55_85), .C2 (n_49_86) );
AOI211_X1 g_64_80 (.ZN (n_64_80), .A (n_64_82), .B (n_61_82), .C1 (n_57_84), .C2 (n_51_85) );
AOI211_X1 g_66_79 (.ZN (n_66_79), .A (n_62_81), .B (n_63_81), .C1 (n_59_83), .C2 (n_53_84) );
AOI211_X1 g_68_78 (.ZN (n_68_78), .A (n_64_80), .B (n_65_80), .C1 (n_61_82), .C2 (n_55_85) );
AOI211_X1 g_70_79 (.ZN (n_70_79), .A (n_66_79), .B (n_64_82), .C1 (n_63_81), .C2 (n_57_84) );
AOI211_X1 g_68_80 (.ZN (n_68_80), .A (n_68_78), .B (n_62_81), .C1 (n_65_80), .C2 (n_59_83) );
AOI211_X1 g_69_78 (.ZN (n_69_78), .A (n_70_79), .B (n_64_80), .C1 (n_64_82), .C2 (n_61_82) );
AOI211_X1 g_71_79 (.ZN (n_71_79), .A (n_68_80), .B (n_66_79), .C1 (n_62_81), .C2 (n_63_81) );
AOI211_X1 g_73_78 (.ZN (n_73_78), .A (n_69_78), .B (n_68_78), .C1 (n_64_80), .C2 (n_65_80) );
AOI211_X1 g_75_77 (.ZN (n_75_77), .A (n_71_79), .B (n_70_79), .C1 (n_66_79), .C2 (n_64_82) );
AOI211_X1 g_77_76 (.ZN (n_77_76), .A (n_73_78), .B (n_68_80), .C1 (n_68_78), .C2 (n_62_81) );
AOI211_X1 g_79_75 (.ZN (n_79_75), .A (n_75_77), .B (n_69_78), .C1 (n_70_79), .C2 (n_64_80) );
AOI211_X1 g_81_74 (.ZN (n_81_74), .A (n_77_76), .B (n_71_79), .C1 (n_68_80), .C2 (n_66_79) );
AOI211_X1 g_83_73 (.ZN (n_83_73), .A (n_79_75), .B (n_73_78), .C1 (n_69_78), .C2 (n_68_78) );
AOI211_X1 g_82_75 (.ZN (n_82_75), .A (n_81_74), .B (n_75_77), .C1 (n_71_79), .C2 (n_70_79) );
AOI211_X1 g_84_74 (.ZN (n_84_74), .A (n_83_73), .B (n_77_76), .C1 (n_73_78), .C2 (n_68_80) );
AOI211_X1 g_86_73 (.ZN (n_86_73), .A (n_82_75), .B (n_79_75), .C1 (n_75_77), .C2 (n_69_78) );
AOI211_X1 g_88_72 (.ZN (n_88_72), .A (n_84_74), .B (n_81_74), .C1 (n_77_76), .C2 (n_71_79) );
AOI211_X1 g_90_71 (.ZN (n_90_71), .A (n_86_73), .B (n_83_73), .C1 (n_79_75), .C2 (n_73_78) );
AOI211_X1 g_92_72 (.ZN (n_92_72), .A (n_88_72), .B (n_82_75), .C1 (n_81_74), .C2 (n_75_77) );
AOI211_X1 g_94_73 (.ZN (n_94_73), .A (n_90_71), .B (n_84_74), .C1 (n_83_73), .C2 (n_77_76) );
AOI211_X1 g_96_74 (.ZN (n_96_74), .A (n_92_72), .B (n_86_73), .C1 (n_82_75), .C2 (n_79_75) );
AOI211_X1 g_98_75 (.ZN (n_98_75), .A (n_94_73), .B (n_88_72), .C1 (n_84_74), .C2 (n_81_74) );
AOI211_X1 g_97_77 (.ZN (n_97_77), .A (n_96_74), .B (n_90_71), .C1 (n_86_73), .C2 (n_83_73) );
AOI211_X1 g_95_76 (.ZN (n_95_76), .A (n_98_75), .B (n_92_72), .C1 (n_88_72), .C2 (n_82_75) );
AOI211_X1 g_97_75 (.ZN (n_97_75), .A (n_97_77), .B (n_94_73), .C1 (n_90_71), .C2 (n_84_74) );
AOI211_X1 g_95_74 (.ZN (n_95_74), .A (n_95_76), .B (n_96_74), .C1 (n_92_72), .C2 (n_86_73) );
AOI211_X1 g_93_75 (.ZN (n_93_75), .A (n_97_75), .B (n_98_75), .C1 (n_94_73), .C2 (n_88_72) );
AOI211_X1 g_91_74 (.ZN (n_91_74), .A (n_95_74), .B (n_97_77), .C1 (n_96_74), .C2 (n_90_71) );
AOI211_X1 g_93_73 (.ZN (n_93_73), .A (n_93_75), .B (n_95_76), .C1 (n_98_75), .C2 (n_92_72) );
AOI211_X1 g_92_71 (.ZN (n_92_71), .A (n_91_74), .B (n_97_75), .C1 (n_97_77), .C2 (n_94_73) );
AOI211_X1 g_90_72 (.ZN (n_90_72), .A (n_93_73), .B (n_95_74), .C1 (n_95_76), .C2 (n_96_74) );
AOI211_X1 g_88_71 (.ZN (n_88_71), .A (n_92_71), .B (n_93_75), .C1 (n_97_75), .C2 (n_98_75) );
AOI211_X1 g_86_72 (.ZN (n_86_72), .A (n_90_72), .B (n_91_74), .C1 (n_95_74), .C2 (n_97_77) );
AOI211_X1 g_84_73 (.ZN (n_84_73), .A (n_88_71), .B (n_93_73), .C1 (n_93_75), .C2 (n_95_76) );
AOI211_X1 g_82_74 (.ZN (n_82_74), .A (n_86_72), .B (n_92_71), .C1 (n_91_74), .C2 (n_97_75) );
AOI211_X1 g_80_75 (.ZN (n_80_75), .A (n_84_73), .B (n_90_72), .C1 (n_93_73), .C2 (n_95_74) );
AOI211_X1 g_78_76 (.ZN (n_78_76), .A (n_82_74), .B (n_88_71), .C1 (n_92_71), .C2 (n_93_75) );
AOI211_X1 g_76_77 (.ZN (n_76_77), .A (n_80_75), .B (n_86_72), .C1 (n_90_72), .C2 (n_91_74) );
AOI211_X1 g_74_78 (.ZN (n_74_78), .A (n_78_76), .B (n_84_73), .C1 (n_88_71), .C2 (n_93_73) );
AOI211_X1 g_72_79 (.ZN (n_72_79), .A (n_76_77), .B (n_82_74), .C1 (n_86_72), .C2 (n_92_71) );
AOI211_X1 g_70_80 (.ZN (n_70_80), .A (n_74_78), .B (n_80_75), .C1 (n_84_73), .C2 (n_90_72) );
AOI211_X1 g_71_78 (.ZN (n_71_78), .A (n_72_79), .B (n_78_76), .C1 (n_82_74), .C2 (n_88_71) );
AOI211_X1 g_69_79 (.ZN (n_69_79), .A (n_70_80), .B (n_76_77), .C1 (n_80_75), .C2 (n_86_72) );
AOI211_X1 g_67_80 (.ZN (n_67_80), .A (n_71_78), .B (n_74_78), .C1 (n_78_76), .C2 (n_84_73) );
AOI211_X1 g_65_81 (.ZN (n_65_81), .A (n_69_79), .B (n_72_79), .C1 (n_76_77), .C2 (n_82_74) );
AOI211_X1 g_63_82 (.ZN (n_63_82), .A (n_67_80), .B (n_70_80), .C1 (n_74_78), .C2 (n_80_75) );
AOI211_X1 g_61_81 (.ZN (n_61_81), .A (n_65_81), .B (n_71_78), .C1 (n_72_79), .C2 (n_78_76) );
AOI211_X1 g_59_82 (.ZN (n_59_82), .A (n_63_82), .B (n_69_79), .C1 (n_70_80), .C2 (n_76_77) );
AOI211_X1 g_57_83 (.ZN (n_57_83), .A (n_61_81), .B (n_67_80), .C1 (n_71_78), .C2 (n_74_78) );
AOI211_X1 g_55_84 (.ZN (n_55_84), .A (n_59_82), .B (n_65_81), .C1 (n_69_79), .C2 (n_72_79) );
AOI211_X1 g_53_85 (.ZN (n_53_85), .A (n_57_83), .B (n_63_82), .C1 (n_67_80), .C2 (n_70_80) );
AOI211_X1 g_51_86 (.ZN (n_51_86), .A (n_55_84), .B (n_61_81), .C1 (n_65_81), .C2 (n_71_78) );
AOI211_X1 g_52_84 (.ZN (n_52_84), .A (n_53_85), .B (n_59_82), .C1 (n_63_82), .C2 (n_69_79) );
AOI211_X1 g_50_85 (.ZN (n_50_85), .A (n_51_86), .B (n_57_83), .C1 (n_61_81), .C2 (n_67_80) );
AOI211_X1 g_48_86 (.ZN (n_48_86), .A (n_52_84), .B (n_55_84), .C1 (n_59_82), .C2 (n_65_81) );
AOI211_X1 g_46_87 (.ZN (n_46_87), .A (n_50_85), .B (n_53_85), .C1 (n_57_83), .C2 (n_63_82) );
AOI211_X1 g_44_88 (.ZN (n_44_88), .A (n_48_86), .B (n_51_86), .C1 (n_55_84), .C2 (n_61_81) );
AOI211_X1 g_46_89 (.ZN (n_46_89), .A (n_46_87), .B (n_52_84), .C1 (n_53_85), .C2 (n_59_82) );
AOI211_X1 g_48_88 (.ZN (n_48_88), .A (n_44_88), .B (n_50_85), .C1 (n_51_86), .C2 (n_57_83) );
AOI211_X1 g_50_87 (.ZN (n_50_87), .A (n_46_89), .B (n_48_86), .C1 (n_52_84), .C2 (n_55_84) );
AOI211_X1 g_52_86 (.ZN (n_52_86), .A (n_48_88), .B (n_46_87), .C1 (n_50_85), .C2 (n_53_85) );
AOI211_X1 g_54_85 (.ZN (n_54_85), .A (n_50_87), .B (n_44_88), .C1 (n_48_86), .C2 (n_51_86) );
AOI211_X1 g_53_87 (.ZN (n_53_87), .A (n_52_86), .B (n_46_89), .C1 (n_46_87), .C2 (n_52_84) );
AOI211_X1 g_55_86 (.ZN (n_55_86), .A (n_54_85), .B (n_48_88), .C1 (n_44_88), .C2 (n_50_85) );
AOI211_X1 g_57_85 (.ZN (n_57_85), .A (n_53_87), .B (n_50_87), .C1 (n_46_89), .C2 (n_48_86) );
AOI211_X1 g_59_84 (.ZN (n_59_84), .A (n_55_86), .B (n_52_86), .C1 (n_48_88), .C2 (n_46_87) );
AOI211_X1 g_61_83 (.ZN (n_61_83), .A (n_57_85), .B (n_54_85), .C1 (n_50_87), .C2 (n_44_88) );
AOI211_X1 g_60_85 (.ZN (n_60_85), .A (n_59_84), .B (n_53_87), .C1 (n_52_86), .C2 (n_46_89) );
AOI211_X1 g_58_84 (.ZN (n_58_84), .A (n_61_83), .B (n_55_86), .C1 (n_54_85), .C2 (n_48_88) );
AOI211_X1 g_60_83 (.ZN (n_60_83), .A (n_60_85), .B (n_57_85), .C1 (n_53_87), .C2 (n_50_87) );
AOI211_X1 g_62_82 (.ZN (n_62_82), .A (n_58_84), .B (n_59_84), .C1 (n_55_86), .C2 (n_52_86) );
AOI211_X1 g_64_81 (.ZN (n_64_81), .A (n_60_83), .B (n_61_83), .C1 (n_57_85), .C2 (n_54_85) );
AOI211_X1 g_63_83 (.ZN (n_63_83), .A (n_62_82), .B (n_60_85), .C1 (n_59_84), .C2 (n_53_87) );
AOI211_X1 g_65_82 (.ZN (n_65_82), .A (n_64_81), .B (n_58_84), .C1 (n_61_83), .C2 (n_55_86) );
AOI211_X1 g_67_81 (.ZN (n_67_81), .A (n_63_83), .B (n_60_83), .C1 (n_60_85), .C2 (n_57_85) );
AOI211_X1 g_69_80 (.ZN (n_69_80), .A (n_65_82), .B (n_62_82), .C1 (n_58_84), .C2 (n_59_84) );
AOI211_X1 g_71_81 (.ZN (n_71_81), .A (n_67_81), .B (n_64_81), .C1 (n_60_83), .C2 (n_61_83) );
AOI211_X1 g_73_80 (.ZN (n_73_80), .A (n_69_80), .B (n_63_83), .C1 (n_62_82), .C2 (n_60_85) );
AOI211_X1 g_75_79 (.ZN (n_75_79), .A (n_71_81), .B (n_65_82), .C1 (n_64_81), .C2 (n_58_84) );
AOI211_X1 g_77_78 (.ZN (n_77_78), .A (n_73_80), .B (n_67_81), .C1 (n_63_83), .C2 (n_60_83) );
AOI211_X1 g_79_77 (.ZN (n_79_77), .A (n_75_79), .B (n_69_80), .C1 (n_65_82), .C2 (n_62_82) );
AOI211_X1 g_81_76 (.ZN (n_81_76), .A (n_77_78), .B (n_71_81), .C1 (n_67_81), .C2 (n_64_81) );
AOI211_X1 g_83_75 (.ZN (n_83_75), .A (n_79_77), .B (n_73_80), .C1 (n_69_80), .C2 (n_63_83) );
AOI211_X1 g_85_74 (.ZN (n_85_74), .A (n_81_76), .B (n_75_79), .C1 (n_71_81), .C2 (n_65_82) );
AOI211_X1 g_87_73 (.ZN (n_87_73), .A (n_83_75), .B (n_77_78), .C1 (n_73_80), .C2 (n_67_81) );
AOI211_X1 g_89_74 (.ZN (n_89_74), .A (n_85_74), .B (n_79_77), .C1 (n_75_79), .C2 (n_69_80) );
AOI211_X1 g_91_73 (.ZN (n_91_73), .A (n_87_73), .B (n_81_76), .C1 (n_77_78), .C2 (n_71_81) );
AOI211_X1 g_93_74 (.ZN (n_93_74), .A (n_89_74), .B (n_83_75), .C1 (n_79_77), .C2 (n_73_80) );
AOI211_X1 g_95_75 (.ZN (n_95_75), .A (n_91_73), .B (n_85_74), .C1 (n_81_76), .C2 (n_75_79) );
AOI211_X1 g_97_76 (.ZN (n_97_76), .A (n_93_74), .B (n_87_73), .C1 (n_83_75), .C2 (n_77_78) );
AOI211_X1 g_99_77 (.ZN (n_99_77), .A (n_95_75), .B (n_89_74), .C1 (n_85_74), .C2 (n_79_77) );
AOI211_X1 g_100_79 (.ZN (n_100_79), .A (n_97_76), .B (n_91_73), .C1 (n_87_73), .C2 (n_81_76) );
AOI211_X1 g_98_78 (.ZN (n_98_78), .A (n_99_77), .B (n_93_74), .C1 (n_89_74), .C2 (n_83_75) );
AOI211_X1 g_96_77 (.ZN (n_96_77), .A (n_100_79), .B (n_95_75), .C1 (n_91_73), .C2 (n_85_74) );
AOI211_X1 g_94_76 (.ZN (n_94_76), .A (n_98_78), .B (n_97_76), .C1 (n_93_74), .C2 (n_87_73) );
AOI211_X1 g_92_75 (.ZN (n_92_75), .A (n_96_77), .B (n_99_77), .C1 (n_95_75), .C2 (n_89_74) );
AOI211_X1 g_90_74 (.ZN (n_90_74), .A (n_94_76), .B (n_100_79), .C1 (n_97_76), .C2 (n_91_73) );
AOI211_X1 g_91_72 (.ZN (n_91_72), .A (n_92_75), .B (n_98_78), .C1 (n_99_77), .C2 (n_93_74) );
AOI211_X1 g_89_71 (.ZN (n_89_71), .A (n_90_74), .B (n_96_77), .C1 (n_100_79), .C2 (n_95_75) );
AOI211_X1 g_88_73 (.ZN (n_88_73), .A (n_91_72), .B (n_94_76), .C1 (n_98_78), .C2 (n_97_76) );
AOI211_X1 g_87_75 (.ZN (n_87_75), .A (n_89_71), .B (n_92_75), .C1 (n_96_77), .C2 (n_99_77) );
AOI211_X1 g_85_76 (.ZN (n_85_76), .A (n_88_73), .B (n_90_74), .C1 (n_94_76), .C2 (n_100_79) );
AOI211_X1 g_86_74 (.ZN (n_86_74), .A (n_87_75), .B (n_91_72), .C1 (n_92_75), .C2 (n_98_78) );
AOI211_X1 g_87_72 (.ZN (n_87_72), .A (n_85_76), .B (n_89_71), .C1 (n_90_74), .C2 (n_96_77) );
AOI211_X1 g_89_73 (.ZN (n_89_73), .A (n_86_74), .B (n_88_73), .C1 (n_91_72), .C2 (n_94_76) );
AOI211_X1 g_88_75 (.ZN (n_88_75), .A (n_87_72), .B (n_87_75), .C1 (n_89_71), .C2 (n_92_75) );
AOI211_X1 g_90_76 (.ZN (n_90_76), .A (n_89_73), .B (n_85_76), .C1 (n_88_73), .C2 (n_90_74) );
AOI211_X1 g_92_77 (.ZN (n_92_77), .A (n_88_75), .B (n_86_74), .C1 (n_87_75), .C2 (n_91_72) );
AOI211_X1 g_91_75 (.ZN (n_91_75), .A (n_90_76), .B (n_87_72), .C1 (n_85_76), .C2 (n_89_71) );
AOI211_X1 g_90_73 (.ZN (n_90_73), .A (n_92_77), .B (n_89_73), .C1 (n_86_74), .C2 (n_88_73) );
AOI211_X1 g_88_74 (.ZN (n_88_74), .A (n_91_75), .B (n_88_75), .C1 (n_87_72), .C2 (n_87_75) );
AOI211_X1 g_89_76 (.ZN (n_89_76), .A (n_90_73), .B (n_90_76), .C1 (n_89_73), .C2 (n_85_76) );
AOI211_X1 g_87_77 (.ZN (n_87_77), .A (n_88_74), .B (n_92_77), .C1 (n_88_75), .C2 (n_86_74) );
AOI211_X1 g_86_75 (.ZN (n_86_75), .A (n_89_76), .B (n_91_75), .C1 (n_90_76), .C2 (n_87_72) );
AOI211_X1 g_85_73 (.ZN (n_85_73), .A (n_87_77), .B (n_90_73), .C1 (n_92_77), .C2 (n_89_73) );
AOI211_X1 g_83_74 (.ZN (n_83_74), .A (n_86_75), .B (n_88_74), .C1 (n_91_75), .C2 (n_88_75) );
AOI211_X1 g_81_75 (.ZN (n_81_75), .A (n_85_73), .B (n_89_76), .C1 (n_90_73), .C2 (n_90_76) );
AOI211_X1 g_79_76 (.ZN (n_79_76), .A (n_83_74), .B (n_87_77), .C1 (n_88_74), .C2 (n_92_77) );
AOI211_X1 g_77_77 (.ZN (n_77_77), .A (n_81_75), .B (n_86_75), .C1 (n_89_76), .C2 (n_91_75) );
AOI211_X1 g_75_78 (.ZN (n_75_78), .A (n_79_76), .B (n_85_73), .C1 (n_87_77), .C2 (n_90_73) );
AOI211_X1 g_73_79 (.ZN (n_73_79), .A (n_77_77), .B (n_83_74), .C1 (n_86_75), .C2 (n_88_74) );
AOI211_X1 g_71_80 (.ZN (n_71_80), .A (n_75_78), .B (n_81_75), .C1 (n_85_73), .C2 (n_89_76) );
AOI211_X1 g_69_81 (.ZN (n_69_81), .A (n_73_79), .B (n_79_76), .C1 (n_83_74), .C2 (n_87_77) );
AOI211_X1 g_67_82 (.ZN (n_67_82), .A (n_71_80), .B (n_77_77), .C1 (n_81_75), .C2 (n_86_75) );
AOI211_X1 g_65_83 (.ZN (n_65_83), .A (n_69_81), .B (n_75_78), .C1 (n_79_76), .C2 (n_85_73) );
AOI211_X1 g_66_81 (.ZN (n_66_81), .A (n_67_82), .B (n_73_79), .C1 (n_77_77), .C2 (n_83_74) );
AOI211_X1 g_68_82 (.ZN (n_68_82), .A (n_65_83), .B (n_71_80), .C1 (n_75_78), .C2 (n_81_75) );
AOI211_X1 g_70_81 (.ZN (n_70_81), .A (n_66_81), .B (n_69_81), .C1 (n_73_79), .C2 (n_79_76) );
AOI211_X1 g_72_80 (.ZN (n_72_80), .A (n_68_82), .B (n_67_82), .C1 (n_71_80), .C2 (n_77_77) );
AOI211_X1 g_74_79 (.ZN (n_74_79), .A (n_70_81), .B (n_65_83), .C1 (n_69_81), .C2 (n_75_78) );
AOI211_X1 g_76_78 (.ZN (n_76_78), .A (n_72_80), .B (n_66_81), .C1 (n_67_82), .C2 (n_73_79) );
AOI211_X1 g_78_77 (.ZN (n_78_77), .A (n_74_79), .B (n_68_82), .C1 (n_65_83), .C2 (n_71_80) );
AOI211_X1 g_80_76 (.ZN (n_80_76), .A (n_76_78), .B (n_70_81), .C1 (n_66_81), .C2 (n_69_81) );
AOI211_X1 g_79_78 (.ZN (n_79_78), .A (n_78_77), .B (n_72_80), .C1 (n_68_82), .C2 (n_67_82) );
AOI211_X1 g_81_77 (.ZN (n_81_77), .A (n_80_76), .B (n_74_79), .C1 (n_70_81), .C2 (n_65_83) );
AOI211_X1 g_83_76 (.ZN (n_83_76), .A (n_79_78), .B (n_76_78), .C1 (n_72_80), .C2 (n_66_81) );
AOI211_X1 g_85_75 (.ZN (n_85_75), .A (n_81_77), .B (n_78_77), .C1 (n_74_79), .C2 (n_68_82) );
AOI211_X1 g_87_74 (.ZN (n_87_74), .A (n_83_76), .B (n_80_76), .C1 (n_76_78), .C2 (n_70_81) );
AOI211_X1 g_89_75 (.ZN (n_89_75), .A (n_85_75), .B (n_79_78), .C1 (n_78_77), .C2 (n_72_80) );
AOI211_X1 g_87_76 (.ZN (n_87_76), .A (n_87_74), .B (n_81_77), .C1 (n_80_76), .C2 (n_74_79) );
AOI211_X1 g_85_77 (.ZN (n_85_77), .A (n_89_75), .B (n_83_76), .C1 (n_79_78), .C2 (n_76_78) );
AOI211_X1 g_84_75 (.ZN (n_84_75), .A (n_87_76), .B (n_85_75), .C1 (n_81_77), .C2 (n_78_77) );
AOI211_X1 g_82_76 (.ZN (n_82_76), .A (n_85_77), .B (n_87_74), .C1 (n_83_76), .C2 (n_80_76) );
AOI211_X1 g_80_77 (.ZN (n_80_77), .A (n_84_75), .B (n_89_75), .C1 (n_85_75), .C2 (n_79_78) );
AOI211_X1 g_78_78 (.ZN (n_78_78), .A (n_82_76), .B (n_87_76), .C1 (n_87_74), .C2 (n_81_77) );
AOI211_X1 g_76_79 (.ZN (n_76_79), .A (n_80_77), .B (n_85_77), .C1 (n_89_75), .C2 (n_83_76) );
AOI211_X1 g_74_80 (.ZN (n_74_80), .A (n_78_78), .B (n_84_75), .C1 (n_87_76), .C2 (n_85_75) );
AOI211_X1 g_72_81 (.ZN (n_72_81), .A (n_76_79), .B (n_82_76), .C1 (n_85_77), .C2 (n_87_74) );
AOI211_X1 g_70_82 (.ZN (n_70_82), .A (n_74_80), .B (n_80_77), .C1 (n_84_75), .C2 (n_89_75) );
AOI211_X1 g_68_81 (.ZN (n_68_81), .A (n_72_81), .B (n_78_78), .C1 (n_82_76), .C2 (n_87_76) );
AOI211_X1 g_66_82 (.ZN (n_66_82), .A (n_70_82), .B (n_76_79), .C1 (n_80_77), .C2 (n_85_77) );
AOI211_X1 g_64_83 (.ZN (n_64_83), .A (n_68_81), .B (n_74_80), .C1 (n_78_78), .C2 (n_84_75) );
AOI211_X1 g_62_84 (.ZN (n_62_84), .A (n_66_82), .B (n_72_81), .C1 (n_76_79), .C2 (n_82_76) );
AOI211_X1 g_64_85 (.ZN (n_64_85), .A (n_64_83), .B (n_70_82), .C1 (n_74_80), .C2 (n_80_77) );
AOI211_X1 g_66_84 (.ZN (n_66_84), .A (n_62_84), .B (n_68_81), .C1 (n_72_81), .C2 (n_78_78) );
AOI211_X1 g_68_83 (.ZN (n_68_83), .A (n_64_85), .B (n_66_82), .C1 (n_70_82), .C2 (n_76_79) );
AOI211_X1 g_67_85 (.ZN (n_67_85), .A (n_66_84), .B (n_64_83), .C1 (n_68_81), .C2 (n_74_80) );
AOI211_X1 g_66_83 (.ZN (n_66_83), .A (n_68_83), .B (n_62_84), .C1 (n_66_82), .C2 (n_72_81) );
AOI211_X1 g_64_84 (.ZN (n_64_84), .A (n_67_85), .B (n_64_85), .C1 (n_64_83), .C2 (n_70_82) );
AOI211_X1 g_62_83 (.ZN (n_62_83), .A (n_66_83), .B (n_66_84), .C1 (n_62_84), .C2 (n_68_81) );
AOI211_X1 g_60_84 (.ZN (n_60_84), .A (n_64_84), .B (n_68_83), .C1 (n_64_85), .C2 (n_66_82) );
AOI211_X1 g_58_85 (.ZN (n_58_85), .A (n_62_83), .B (n_67_85), .C1 (n_66_84), .C2 (n_64_83) );
AOI211_X1 g_56_86 (.ZN (n_56_86), .A (n_60_84), .B (n_66_83), .C1 (n_68_83), .C2 (n_62_84) );
AOI211_X1 g_54_87 (.ZN (n_54_87), .A (n_58_85), .B (n_64_84), .C1 (n_67_85), .C2 (n_64_85) );
AOI211_X1 g_52_88 (.ZN (n_52_88), .A (n_56_86), .B (n_62_83), .C1 (n_66_83), .C2 (n_66_84) );
AOI211_X1 g_53_86 (.ZN (n_53_86), .A (n_54_87), .B (n_60_84), .C1 (n_64_84), .C2 (n_68_83) );
AOI211_X1 g_51_87 (.ZN (n_51_87), .A (n_52_88), .B (n_58_85), .C1 (n_62_83), .C2 (n_67_85) );
AOI211_X1 g_49_88 (.ZN (n_49_88), .A (n_53_86), .B (n_56_86), .C1 (n_60_84), .C2 (n_66_83) );
AOI211_X1 g_50_86 (.ZN (n_50_86), .A (n_51_87), .B (n_54_87), .C1 (n_58_85), .C2 (n_64_84) );
AOI211_X1 g_48_87 (.ZN (n_48_87), .A (n_49_88), .B (n_52_88), .C1 (n_56_86), .C2 (n_62_83) );
AOI211_X1 g_46_88 (.ZN (n_46_88), .A (n_50_86), .B (n_53_86), .C1 (n_54_87), .C2 (n_60_84) );
AOI211_X1 g_44_89 (.ZN (n_44_89), .A (n_48_87), .B (n_51_87), .C1 (n_52_88), .C2 (n_58_85) );
AOI211_X1 g_42_90 (.ZN (n_42_90), .A (n_46_88), .B (n_49_88), .C1 (n_53_86), .C2 (n_56_86) );
AOI211_X1 g_40_91 (.ZN (n_40_91), .A (n_44_89), .B (n_50_86), .C1 (n_51_87), .C2 (n_54_87) );
AOI211_X1 g_41_89 (.ZN (n_41_89), .A (n_42_90), .B (n_48_87), .C1 (n_49_88), .C2 (n_52_88) );
AOI211_X1 g_39_90 (.ZN (n_39_90), .A (n_40_91), .B (n_46_88), .C1 (n_50_86), .C2 (n_53_86) );
AOI211_X1 g_37_91 (.ZN (n_37_91), .A (n_41_89), .B (n_44_89), .C1 (n_48_87), .C2 (n_51_87) );
AOI211_X1 g_35_92 (.ZN (n_35_92), .A (n_39_90), .B (n_42_90), .C1 (n_46_88), .C2 (n_49_88) );
AOI211_X1 g_33_93 (.ZN (n_33_93), .A (n_37_91), .B (n_40_91), .C1 (n_44_89), .C2 (n_50_86) );
AOI211_X1 g_31_92 (.ZN (n_31_92), .A (n_35_92), .B (n_41_89), .C1 (n_42_90), .C2 (n_48_87) );
AOI211_X1 g_29_93 (.ZN (n_29_93), .A (n_33_93), .B (n_39_90), .C1 (n_40_91), .C2 (n_46_88) );
AOI211_X1 g_27_94 (.ZN (n_27_94), .A (n_31_92), .B (n_37_91), .C1 (n_41_89), .C2 (n_44_89) );
AOI211_X1 g_25_95 (.ZN (n_25_95), .A (n_29_93), .B (n_35_92), .C1 (n_39_90), .C2 (n_42_90) );
AOI211_X1 g_23_96 (.ZN (n_23_96), .A (n_27_94), .B (n_33_93), .C1 (n_37_91), .C2 (n_40_91) );
AOI211_X1 g_24_98 (.ZN (n_24_98), .A (n_25_95), .B (n_31_92), .C1 (n_35_92), .C2 (n_41_89) );
AOI211_X1 g_26_97 (.ZN (n_26_97), .A (n_23_96), .B (n_29_93), .C1 (n_33_93), .C2 (n_39_90) );
AOI211_X1 g_28_96 (.ZN (n_28_96), .A (n_24_98), .B (n_27_94), .C1 (n_31_92), .C2 (n_37_91) );
AOI211_X1 g_30_95 (.ZN (n_30_95), .A (n_26_97), .B (n_25_95), .C1 (n_29_93), .C2 (n_35_92) );
AOI211_X1 g_32_94 (.ZN (n_32_94), .A (n_28_96), .B (n_23_96), .C1 (n_27_94), .C2 (n_33_93) );
AOI211_X1 g_34_95 (.ZN (n_34_95), .A (n_30_95), .B (n_24_98), .C1 (n_25_95), .C2 (n_31_92) );
AOI211_X1 g_36_94 (.ZN (n_36_94), .A (n_32_94), .B (n_26_97), .C1 (n_23_96), .C2 (n_29_93) );
AOI211_X1 g_37_92 (.ZN (n_37_92), .A (n_34_95), .B (n_28_96), .C1 (n_24_98), .C2 (n_27_94) );
AOI211_X1 g_39_91 (.ZN (n_39_91), .A (n_36_94), .B (n_30_95), .C1 (n_26_97), .C2 (n_25_95) );
AOI211_X1 g_41_90 (.ZN (n_41_90), .A (n_37_92), .B (n_32_94), .C1 (n_28_96), .C2 (n_23_96) );
AOI211_X1 g_40_92 (.ZN (n_40_92), .A (n_39_91), .B (n_34_95), .C1 (n_30_95), .C2 (n_24_98) );
AOI211_X1 g_38_93 (.ZN (n_38_93), .A (n_41_90), .B (n_36_94), .C1 (n_32_94), .C2 (n_26_97) );
AOI211_X1 g_37_95 (.ZN (n_37_95), .A (n_40_92), .B (n_37_92), .C1 (n_34_95), .C2 (n_28_96) );
AOI211_X1 g_36_93 (.ZN (n_36_93), .A (n_38_93), .B (n_39_91), .C1 (n_36_94), .C2 (n_30_95) );
AOI211_X1 g_38_92 (.ZN (n_38_92), .A (n_37_95), .B (n_41_90), .C1 (n_37_92), .C2 (n_32_94) );
AOI211_X1 g_37_94 (.ZN (n_37_94), .A (n_36_93), .B (n_40_92), .C1 (n_39_91), .C2 (n_34_95) );
AOI211_X1 g_39_93 (.ZN (n_39_93), .A (n_38_92), .B (n_38_93), .C1 (n_41_90), .C2 (n_36_94) );
AOI211_X1 g_41_92 (.ZN (n_41_92), .A (n_37_94), .B (n_37_95), .C1 (n_40_92), .C2 (n_37_92) );
AOI211_X1 g_43_91 (.ZN (n_43_91), .A (n_39_93), .B (n_36_93), .C1 (n_38_93), .C2 (n_39_91) );
AOI211_X1 g_45_90 (.ZN (n_45_90), .A (n_41_92), .B (n_38_92), .C1 (n_37_95), .C2 (n_41_90) );
AOI211_X1 g_47_89 (.ZN (n_47_89), .A (n_43_91), .B (n_37_94), .C1 (n_36_93), .C2 (n_40_92) );
AOI211_X1 g_49_90 (.ZN (n_49_90), .A (n_45_90), .B (n_39_93), .C1 (n_38_92), .C2 (n_38_93) );
AOI211_X1 g_50_88 (.ZN (n_50_88), .A (n_47_89), .B (n_41_92), .C1 (n_37_94), .C2 (n_37_95) );
AOI211_X1 g_52_87 (.ZN (n_52_87), .A (n_49_90), .B (n_43_91), .C1 (n_39_93), .C2 (n_36_93) );
AOI211_X1 g_54_86 (.ZN (n_54_86), .A (n_50_88), .B (n_45_90), .C1 (n_41_92), .C2 (n_38_92) );
AOI211_X1 g_56_85 (.ZN (n_56_85), .A (n_52_87), .B (n_47_89), .C1 (n_43_91), .C2 (n_37_94) );
AOI211_X1 g_58_86 (.ZN (n_58_86), .A (n_54_86), .B (n_49_90), .C1 (n_45_90), .C2 (n_39_93) );
AOI211_X1 g_56_87 (.ZN (n_56_87), .A (n_56_85), .B (n_50_88), .C1 (n_47_89), .C2 (n_41_92) );
AOI211_X1 g_54_88 (.ZN (n_54_88), .A (n_58_86), .B (n_52_87), .C1 (n_49_90), .C2 (n_43_91) );
AOI211_X1 g_52_89 (.ZN (n_52_89), .A (n_56_87), .B (n_54_86), .C1 (n_50_88), .C2 (n_45_90) );
AOI211_X1 g_50_90 (.ZN (n_50_90), .A (n_54_88), .B (n_56_85), .C1 (n_52_87), .C2 (n_47_89) );
AOI211_X1 g_51_88 (.ZN (n_51_88), .A (n_52_89), .B (n_58_86), .C1 (n_54_86), .C2 (n_49_90) );
AOI211_X1 g_49_87 (.ZN (n_49_87), .A (n_50_90), .B (n_56_87), .C1 (n_56_85), .C2 (n_50_88) );
AOI211_X1 g_48_89 (.ZN (n_48_89), .A (n_51_88), .B (n_54_88), .C1 (n_58_86), .C2 (n_52_87) );
AOI211_X1 g_47_91 (.ZN (n_47_91), .A (n_49_87), .B (n_52_89), .C1 (n_56_87), .C2 (n_54_86) );
AOI211_X1 g_45_92 (.ZN (n_45_92), .A (n_48_89), .B (n_50_90), .C1 (n_54_88), .C2 (n_56_85) );
AOI211_X1 g_44_90 (.ZN (n_44_90), .A (n_47_91), .B (n_51_88), .C1 (n_52_89), .C2 (n_58_86) );
AOI211_X1 g_42_91 (.ZN (n_42_91), .A (n_45_92), .B (n_49_87), .C1 (n_50_90), .C2 (n_56_87) );
AOI211_X1 g_43_93 (.ZN (n_43_93), .A (n_44_90), .B (n_48_89), .C1 (n_51_88), .C2 (n_54_88) );
AOI211_X1 g_44_91 (.ZN (n_44_91), .A (n_42_91), .B (n_47_91), .C1 (n_49_87), .C2 (n_52_89) );
AOI211_X1 g_46_90 (.ZN (n_46_90), .A (n_43_93), .B (n_45_92), .C1 (n_48_89), .C2 (n_50_90) );
AOI211_X1 g_47_88 (.ZN (n_47_88), .A (n_44_91), .B (n_44_90), .C1 (n_47_91), .C2 (n_51_88) );
AOI211_X1 g_45_89 (.ZN (n_45_89), .A (n_46_90), .B (n_42_91), .C1 (n_45_92), .C2 (n_49_87) );
AOI211_X1 g_43_90 (.ZN (n_43_90), .A (n_47_88), .B (n_43_93), .C1 (n_44_90), .C2 (n_48_89) );
AOI211_X1 g_41_91 (.ZN (n_41_91), .A (n_45_89), .B (n_44_91), .C1 (n_42_91), .C2 (n_47_91) );
AOI211_X1 g_39_92 (.ZN (n_39_92), .A (n_43_90), .B (n_46_90), .C1 (n_43_93), .C2 (n_45_92) );
AOI211_X1 g_37_93 (.ZN (n_37_93), .A (n_41_91), .B (n_47_88), .C1 (n_44_91), .C2 (n_44_90) );
AOI211_X1 g_39_94 (.ZN (n_39_94), .A (n_39_92), .B (n_45_89), .C1 (n_46_90), .C2 (n_42_91) );
AOI211_X1 g_41_93 (.ZN (n_41_93), .A (n_37_93), .B (n_43_90), .C1 (n_47_88), .C2 (n_43_93) );
AOI211_X1 g_43_92 (.ZN (n_43_92), .A (n_39_94), .B (n_41_91), .C1 (n_45_89), .C2 (n_44_91) );
AOI211_X1 g_45_91 (.ZN (n_45_91), .A (n_41_93), .B (n_39_92), .C1 (n_43_90), .C2 (n_46_90) );
AOI211_X1 g_47_90 (.ZN (n_47_90), .A (n_43_92), .B (n_37_93), .C1 (n_41_91), .C2 (n_47_88) );
AOI211_X1 g_49_89 (.ZN (n_49_89), .A (n_45_91), .B (n_39_94), .C1 (n_39_92), .C2 (n_45_89) );
AOI211_X1 g_48_91 (.ZN (n_48_91), .A (n_47_90), .B (n_41_93), .C1 (n_37_93), .C2 (n_43_90) );
AOI211_X1 g_46_92 (.ZN (n_46_92), .A (n_49_89), .B (n_43_92), .C1 (n_39_94), .C2 (n_41_91) );
AOI211_X1 g_44_93 (.ZN (n_44_93), .A (n_48_91), .B (n_45_91), .C1 (n_41_93), .C2 (n_39_92) );
AOI211_X1 g_42_92 (.ZN (n_42_92), .A (n_46_92), .B (n_47_90), .C1 (n_43_92), .C2 (n_37_93) );
AOI211_X1 g_40_93 (.ZN (n_40_93), .A (n_44_93), .B (n_49_89), .C1 (n_45_91), .C2 (n_39_94) );
AOI211_X1 g_38_94 (.ZN (n_38_94), .A (n_42_92), .B (n_48_91), .C1 (n_47_90), .C2 (n_41_93) );
AOI211_X1 g_36_95 (.ZN (n_36_95), .A (n_40_93), .B (n_46_92), .C1 (n_49_89), .C2 (n_43_92) );
AOI211_X1 g_34_94 (.ZN (n_34_94), .A (n_38_94), .B (n_44_93), .C1 (n_48_91), .C2 (n_45_91) );
AOI211_X1 g_32_93 (.ZN (n_32_93), .A (n_36_95), .B (n_42_92), .C1 (n_46_92), .C2 (n_47_90) );
AOI211_X1 g_30_94 (.ZN (n_30_94), .A (n_34_94), .B (n_40_93), .C1 (n_44_93), .C2 (n_49_89) );
AOI211_X1 g_28_95 (.ZN (n_28_95), .A (n_32_93), .B (n_38_94), .C1 (n_42_92), .C2 (n_48_91) );
AOI211_X1 g_26_96 (.ZN (n_26_96), .A (n_30_94), .B (n_36_95), .C1 (n_40_93), .C2 (n_46_92) );
AOI211_X1 g_24_97 (.ZN (n_24_97), .A (n_28_95), .B (n_34_94), .C1 (n_38_94), .C2 (n_44_93) );
AOI211_X1 g_23_99 (.ZN (n_23_99), .A (n_26_96), .B (n_32_93), .C1 (n_36_95), .C2 (n_42_92) );
AOI211_X1 g_25_98 (.ZN (n_25_98), .A (n_24_97), .B (n_30_94), .C1 (n_34_94), .C2 (n_40_93) );
AOI211_X1 g_27_97 (.ZN (n_27_97), .A (n_23_99), .B (n_28_95), .C1 (n_32_93), .C2 (n_38_94) );
AOI211_X1 g_26_99 (.ZN (n_26_99), .A (n_25_98), .B (n_26_96), .C1 (n_30_94), .C2 (n_36_95) );
AOI211_X1 g_25_97 (.ZN (n_25_97), .A (n_27_97), .B (n_24_97), .C1 (n_28_95), .C2 (n_34_94) );
AOI211_X1 g_27_98 (.ZN (n_27_98), .A (n_26_99), .B (n_23_99), .C1 (n_26_96), .C2 (n_32_93) );
AOI211_X1 g_28_100 (.ZN (n_28_100), .A (n_25_97), .B (n_25_98), .C1 (n_24_97), .C2 (n_30_94) );
AOI211_X1 g_29_98 (.ZN (n_29_98), .A (n_27_98), .B (n_27_97), .C1 (n_23_99), .C2 (n_28_95) );
AOI211_X1 g_27_99 (.ZN (n_27_99), .A (n_28_100), .B (n_26_99), .C1 (n_25_98), .C2 (n_26_96) );
AOI211_X1 g_25_100 (.ZN (n_25_100), .A (n_29_98), .B (n_25_97), .C1 (n_27_97), .C2 (n_24_97) );
AOI211_X1 g_26_98 (.ZN (n_26_98), .A (n_27_99), .B (n_27_98), .C1 (n_26_99), .C2 (n_23_99) );
AOI211_X1 g_28_97 (.ZN (n_28_97), .A (n_25_100), .B (n_28_100), .C1 (n_25_97), .C2 (n_25_98) );
AOI211_X1 g_30_96 (.ZN (n_30_96), .A (n_26_98), .B (n_29_98), .C1 (n_27_98), .C2 (n_27_97) );
AOI211_X1 g_32_95 (.ZN (n_32_95), .A (n_28_97), .B (n_27_99), .C1 (n_28_100), .C2 (n_26_99) );
AOI211_X1 g_31_97 (.ZN (n_31_97), .A (n_30_96), .B (n_25_100), .C1 (n_29_98), .C2 (n_25_97) );
AOI211_X1 g_29_96 (.ZN (n_29_96), .A (n_32_95), .B (n_26_98), .C1 (n_27_99), .C2 (n_27_98) );
AOI211_X1 g_31_95 (.ZN (n_31_95), .A (n_31_97), .B (n_28_97), .C1 (n_25_100), .C2 (n_28_100) );
AOI211_X1 g_33_96 (.ZN (n_33_96), .A (n_29_96), .B (n_30_96), .C1 (n_26_98), .C2 (n_29_98) );
AOI211_X1 g_35_95 (.ZN (n_35_95), .A (n_31_95), .B (n_32_95), .C1 (n_28_97), .C2 (n_27_99) );
AOI211_X1 g_36_97 (.ZN (n_36_97), .A (n_33_96), .B (n_31_97), .C1 (n_30_96), .C2 (n_25_100) );
AOI211_X1 g_34_96 (.ZN (n_34_96), .A (n_35_95), .B (n_29_96), .C1 (n_32_95), .C2 (n_26_98) );
AOI211_X1 g_32_97 (.ZN (n_32_97), .A (n_36_97), .B (n_31_95), .C1 (n_31_97), .C2 (n_28_97) );
AOI211_X1 g_30_98 (.ZN (n_30_98), .A (n_34_96), .B (n_33_96), .C1 (n_29_96), .C2 (n_30_96) );
AOI211_X1 g_29_100 (.ZN (n_29_100), .A (n_32_97), .B (n_35_95), .C1 (n_31_95), .C2 (n_32_95) );
AOI211_X1 g_31_99 (.ZN (n_31_99), .A (n_30_98), .B (n_36_97), .C1 (n_33_96), .C2 (n_31_97) );
AOI211_X1 g_33_100 (.ZN (n_33_100), .A (n_29_100), .B (n_34_96), .C1 (n_35_95), .C2 (n_29_96) );
AOI211_X1 g_34_98 (.ZN (n_34_98), .A (n_31_99), .B (n_32_97), .C1 (n_36_97), .C2 (n_31_95) );
AOI211_X1 g_35_96 (.ZN (n_35_96), .A (n_33_100), .B (n_30_98), .C1 (n_34_96), .C2 (n_33_96) );
AOI211_X1 g_33_95 (.ZN (n_33_95), .A (n_34_98), .B (n_29_100), .C1 (n_32_97), .C2 (n_35_95) );
AOI211_X1 g_31_94 (.ZN (n_31_94), .A (n_35_96), .B (n_31_99), .C1 (n_30_98), .C2 (n_36_97) );
AOI211_X1 g_29_95 (.ZN (n_29_95), .A (n_33_95), .B (n_33_100), .C1 (n_29_100), .C2 (n_34_96) );
AOI211_X1 g_27_96 (.ZN (n_27_96), .A (n_31_94), .B (n_34_98), .C1 (n_31_99), .C2 (n_32_97) );
AOI211_X1 g_28_98 (.ZN (n_28_98), .A (n_29_95), .B (n_35_96), .C1 (n_33_100), .C2 (n_30_98) );
AOI211_X1 g_30_97 (.ZN (n_30_97), .A (n_27_96), .B (n_33_95), .C1 (n_34_98), .C2 (n_29_100) );
AOI211_X1 g_32_96 (.ZN (n_32_96), .A (n_28_98), .B (n_31_94), .C1 (n_35_96), .C2 (n_31_99) );
AOI211_X1 g_31_98 (.ZN (n_31_98), .A (n_30_97), .B (n_29_95), .C1 (n_33_95), .C2 (n_33_100) );
AOI211_X1 g_29_97 (.ZN (n_29_97), .A (n_32_96), .B (n_27_96), .C1 (n_31_94), .C2 (n_34_98) );
AOI211_X1 g_31_96 (.ZN (n_31_96), .A (n_31_98), .B (n_28_98), .C1 (n_29_95), .C2 (n_35_96) );
AOI211_X1 g_33_97 (.ZN (n_33_97), .A (n_29_97), .B (n_30_97), .C1 (n_27_96), .C2 (n_33_95) );
AOI211_X1 g_35_98 (.ZN (n_35_98), .A (n_31_96), .B (n_32_96), .C1 (n_28_98), .C2 (n_31_94) );
AOI211_X1 g_36_100 (.ZN (n_36_100), .A (n_33_97), .B (n_31_98), .C1 (n_30_97), .C2 (n_29_95) );
AOI211_X1 g_34_99 (.ZN (n_34_99), .A (n_35_98), .B (n_29_97), .C1 (n_32_96), .C2 (n_27_96) );
AOI211_X1 g_32_98 (.ZN (n_32_98), .A (n_36_100), .B (n_31_96), .C1 (n_31_98), .C2 (n_28_98) );
AOI211_X1 g_30_99 (.ZN (n_30_99), .A (n_34_99), .B (n_33_97), .C1 (n_29_97), .C2 (n_30_97) );
AOI211_X1 g_32_100 (.ZN (n_32_100), .A (n_32_98), .B (n_35_98), .C1 (n_31_96), .C2 (n_32_96) );
AOI211_X1 g_33_98 (.ZN (n_33_98), .A (n_30_99), .B (n_36_100), .C1 (n_33_97), .C2 (n_31_98) );
AOI211_X1 g_35_97 (.ZN (n_35_97), .A (n_32_100), .B (n_34_99), .C1 (n_35_98), .C2 (n_29_97) );
AOI211_X1 g_37_96 (.ZN (n_37_96), .A (n_33_98), .B (n_32_98), .C1 (n_36_100), .C2 (n_31_96) );
AOI211_X1 g_38_98 (.ZN (n_38_98), .A (n_35_97), .B (n_30_99), .C1 (n_34_99), .C2 (n_33_97) );
AOI211_X1 g_37_100 (.ZN (n_37_100), .A (n_37_96), .B (n_32_100), .C1 (n_32_98), .C2 (n_35_98) );
AOI211_X1 g_35_99 (.ZN (n_35_99), .A (n_38_98), .B (n_33_98), .C1 (n_30_99), .C2 (n_36_100) );
AOI211_X1 g_34_97 (.ZN (n_34_97), .A (n_37_100), .B (n_35_97), .C1 (n_32_100), .C2 (n_34_99) );
AOI211_X1 g_36_98 (.ZN (n_36_98), .A (n_35_99), .B (n_37_96), .C1 (n_33_98), .C2 (n_32_98) );
AOI211_X1 g_38_99 (.ZN (n_38_99), .A (n_34_97), .B (n_38_98), .C1 (n_35_97), .C2 (n_30_99) );
AOI211_X1 g_37_97 (.ZN (n_37_97), .A (n_36_98), .B (n_37_100), .C1 (n_37_96), .C2 (n_32_100) );
AOI211_X1 g_39_96 (.ZN (n_39_96), .A (n_38_99), .B (n_35_99), .C1 (n_38_98), .C2 (n_33_98) );
AOI211_X1 g_40_94 (.ZN (n_40_94), .A (n_37_97), .B (n_34_97), .C1 (n_37_100), .C2 (n_35_97) );
AOI211_X1 g_38_95 (.ZN (n_38_95), .A (n_39_96), .B (n_36_98), .C1 (n_35_99), .C2 (n_37_96) );
AOI211_X1 g_36_96 (.ZN (n_36_96), .A (n_40_94), .B (n_38_99), .C1 (n_34_97), .C2 (n_38_98) );
AOI211_X1 g_37_98 (.ZN (n_37_98), .A (n_38_95), .B (n_37_97), .C1 (n_36_98), .C2 (n_37_100) );
AOI211_X1 g_39_97 (.ZN (n_39_97), .A (n_36_96), .B (n_39_96), .C1 (n_38_99), .C2 (n_35_99) );
AOI211_X1 g_40_95 (.ZN (n_40_95), .A (n_37_98), .B (n_40_94), .C1 (n_37_97), .C2 (n_34_97) );
AOI211_X1 g_38_96 (.ZN (n_38_96), .A (n_39_97), .B (n_38_95), .C1 (n_39_96), .C2 (n_36_98) );
AOI211_X1 g_39_98 (.ZN (n_39_98), .A (n_40_95), .B (n_36_96), .C1 (n_40_94), .C2 (n_38_99) );
AOI211_X1 g_40_100 (.ZN (n_40_100), .A (n_38_96), .B (n_37_98), .C1 (n_38_95), .C2 (n_37_97) );
AOI211_X1 g_42_99 (.ZN (n_42_99), .A (n_39_98), .B (n_39_97), .C1 (n_36_96), .C2 (n_39_96) );
AOI211_X1 g_41_97 (.ZN (n_41_97), .A (n_40_100), .B (n_40_95), .C1 (n_37_98), .C2 (n_40_94) );
AOI211_X1 g_42_95 (.ZN (n_42_95), .A (n_42_99), .B (n_38_96), .C1 (n_39_97), .C2 (n_38_95) );
AOI211_X1 g_40_96 (.ZN (n_40_96), .A (n_41_97), .B (n_39_98), .C1 (n_40_95), .C2 (n_36_96) );
AOI211_X1 g_41_94 (.ZN (n_41_94), .A (n_42_95), .B (n_40_100), .C1 (n_38_96), .C2 (n_37_98) );
AOI211_X1 g_39_95 (.ZN (n_39_95), .A (n_40_96), .B (n_42_99), .C1 (n_39_98), .C2 (n_39_97) );
AOI211_X1 g_38_97 (.ZN (n_38_97), .A (n_41_94), .B (n_41_97), .C1 (n_40_100), .C2 (n_40_95) );
AOI211_X1 g_39_99 (.ZN (n_39_99), .A (n_39_95), .B (n_42_95), .C1 (n_42_99), .C2 (n_38_96) );
AOI211_X1 g_41_98 (.ZN (n_41_98), .A (n_38_97), .B (n_40_96), .C1 (n_41_97), .C2 (n_39_98) );
AOI211_X1 g_43_97 (.ZN (n_43_97), .A (n_39_99), .B (n_41_94), .C1 (n_42_95), .C2 (n_40_100) );
AOI211_X1 g_41_96 (.ZN (n_41_96), .A (n_41_98), .B (n_39_95), .C1 (n_40_96), .C2 (n_42_99) );
AOI211_X1 g_42_94 (.ZN (n_42_94), .A (n_43_97), .B (n_38_97), .C1 (n_41_94), .C2 (n_41_97) );
AOI211_X1 g_44_95 (.ZN (n_44_95), .A (n_41_96), .B (n_39_99), .C1 (n_39_95), .C2 (n_42_95) );
AOI211_X1 g_42_96 (.ZN (n_42_96), .A (n_42_94), .B (n_41_98), .C1 (n_38_97), .C2 (n_40_96) );
AOI211_X1 g_40_97 (.ZN (n_40_97), .A (n_44_95), .B (n_43_97), .C1 (n_39_99), .C2 (n_41_94) );
AOI211_X1 g_42_98 (.ZN (n_42_98), .A (n_42_96), .B (n_41_96), .C1 (n_41_98), .C2 (n_39_95) );
AOI211_X1 g_41_100 (.ZN (n_41_100), .A (n_40_97), .B (n_42_94), .C1 (n_43_97), .C2 (n_38_97) );
AOI211_X1 g_40_98 (.ZN (n_40_98), .A (n_42_98), .B (n_44_95), .C1 (n_41_96), .C2 (n_39_99) );
AOI211_X1 g_42_97 (.ZN (n_42_97), .A (n_41_100), .B (n_42_96), .C1 (n_42_94), .C2 (n_41_98) );
AOI211_X1 g_41_95 (.ZN (n_41_95), .A (n_40_98), .B (n_40_97), .C1 (n_44_95), .C2 (n_43_97) );
AOI211_X1 g_42_93 (.ZN (n_42_93), .A (n_42_97), .B (n_42_98), .C1 (n_42_96), .C2 (n_41_96) );
AOI211_X1 g_43_95 (.ZN (n_43_95), .A (n_41_95), .B (n_41_100), .C1 (n_40_97), .C2 (n_42_94) );
AOI211_X1 g_44_97 (.ZN (n_44_97), .A (n_42_93), .B (n_40_98), .C1 (n_42_98), .C2 (n_44_95) );
AOI211_X1 g_43_99 (.ZN (n_43_99), .A (n_43_95), .B (n_42_97), .C1 (n_41_100), .C2 (n_42_96) );
AOI211_X1 g_45_100 (.ZN (n_45_100), .A (n_44_97), .B (n_41_95), .C1 (n_40_98), .C2 (n_40_97) );
AOI211_X1 g_46_98 (.ZN (n_46_98), .A (n_43_99), .B (n_42_93), .C1 (n_42_97), .C2 (n_42_98) );
AOI211_X1 g_45_96 (.ZN (n_45_96), .A (n_45_100), .B (n_43_95), .C1 (n_41_95), .C2 (n_41_100) );
AOI211_X1 g_44_94 (.ZN (n_44_94), .A (n_46_98), .B (n_44_97), .C1 (n_42_93), .C2 (n_40_98) );
AOI211_X1 g_43_96 (.ZN (n_43_96), .A (n_45_96), .B (n_43_99), .C1 (n_43_95), .C2 (n_42_97) );
AOI211_X1 g_44_98 (.ZN (n_44_98), .A (n_44_94), .B (n_45_100), .C1 (n_44_97), .C2 (n_41_95) );
AOI211_X1 g_46_99 (.ZN (n_46_99), .A (n_43_96), .B (n_46_98), .C1 (n_43_99), .C2 (n_42_93) );
AOI211_X1 g_44_100 (.ZN (n_44_100), .A (n_44_98), .B (n_45_96), .C1 (n_45_100), .C2 (n_43_95) );
AOI211_X1 g_43_98 (.ZN (n_43_98), .A (n_46_99), .B (n_44_94), .C1 (n_46_98), .C2 (n_44_97) );
AOI211_X1 g_45_97 (.ZN (n_45_97), .A (n_44_100), .B (n_43_96), .C1 (n_45_96), .C2 (n_43_99) );
AOI211_X1 g_47_98 (.ZN (n_47_98), .A (n_43_98), .B (n_44_98), .C1 (n_44_94), .C2 (n_45_100) );
AOI211_X1 g_48_100 (.ZN (n_48_100), .A (n_45_97), .B (n_46_99), .C1 (n_43_96), .C2 (n_46_98) );
AOI211_X1 g_50_99 (.ZN (n_50_99), .A (n_47_98), .B (n_44_100), .C1 (n_44_98), .C2 (n_45_96) );
AOI211_X1 g_52_100 (.ZN (n_52_100), .A (n_48_100), .B (n_43_98), .C1 (n_46_99), .C2 (n_44_94) );
AOI211_X1 g_51_98 (.ZN (n_51_98), .A (n_50_99), .B (n_45_97), .C1 (n_44_100), .C2 (n_43_96) );
AOI211_X1 g_49_97 (.ZN (n_49_97), .A (n_52_100), .B (n_47_98), .C1 (n_43_98), .C2 (n_44_98) );
AOI211_X1 g_47_96 (.ZN (n_47_96), .A (n_51_98), .B (n_48_100), .C1 (n_45_97), .C2 (n_46_99) );
AOI211_X1 g_46_94 (.ZN (n_46_94), .A (n_49_97), .B (n_50_99), .C1 (n_47_98), .C2 (n_44_100) );
AOI211_X1 g_48_93 (.ZN (n_48_93), .A (n_47_96), .B (n_52_100), .C1 (n_48_100), .C2 (n_43_98) );
AOI211_X1 g_50_92 (.ZN (n_50_92), .A (n_46_94), .B (n_51_98), .C1 (n_50_99), .C2 (n_45_97) );
AOI211_X1 g_51_90 (.ZN (n_51_90), .A (n_48_93), .B (n_49_97), .C1 (n_52_100), .C2 (n_47_98) );
AOI211_X1 g_53_89 (.ZN (n_53_89), .A (n_50_92), .B (n_47_96), .C1 (n_51_98), .C2 (n_48_100) );
AOI211_X1 g_55_88 (.ZN (n_55_88), .A (n_51_90), .B (n_46_94), .C1 (n_49_97), .C2 (n_50_99) );
AOI211_X1 g_57_87 (.ZN (n_57_87), .A (n_53_89), .B (n_48_93), .C1 (n_47_96), .C2 (n_52_100) );
AOI211_X1 g_59_86 (.ZN (n_59_86), .A (n_55_88), .B (n_50_92), .C1 (n_46_94), .C2 (n_51_98) );
AOI211_X1 g_61_85 (.ZN (n_61_85), .A (n_57_87), .B (n_51_90), .C1 (n_48_93), .C2 (n_49_97) );
AOI211_X1 g_63_84 (.ZN (n_63_84), .A (n_59_86), .B (n_53_89), .C1 (n_50_92), .C2 (n_47_96) );
AOI211_X1 g_62_86 (.ZN (n_62_86), .A (n_61_85), .B (n_55_88), .C1 (n_51_90), .C2 (n_46_94) );
AOI211_X1 g_61_84 (.ZN (n_61_84), .A (n_63_84), .B (n_57_87), .C1 (n_53_89), .C2 (n_48_93) );
AOI211_X1 g_59_85 (.ZN (n_59_85), .A (n_62_86), .B (n_59_86), .C1 (n_55_88), .C2 (n_50_92) );
AOI211_X1 g_57_86 (.ZN (n_57_86), .A (n_61_84), .B (n_61_85), .C1 (n_57_87), .C2 (n_51_90) );
AOI211_X1 g_55_87 (.ZN (n_55_87), .A (n_59_85), .B (n_63_84), .C1 (n_59_86), .C2 (n_53_89) );
AOI211_X1 g_53_88 (.ZN (n_53_88), .A (n_57_86), .B (n_62_86), .C1 (n_61_85), .C2 (n_55_88) );
AOI211_X1 g_51_89 (.ZN (n_51_89), .A (n_55_87), .B (n_61_84), .C1 (n_63_84), .C2 (n_57_87) );
AOI211_X1 g_52_91 (.ZN (n_52_91), .A (n_53_88), .B (n_59_85), .C1 (n_62_86), .C2 (n_59_86) );
AOI211_X1 g_54_90 (.ZN (n_54_90), .A (n_51_89), .B (n_57_86), .C1 (n_61_84), .C2 (n_61_85) );
AOI211_X1 g_56_89 (.ZN (n_56_89), .A (n_52_91), .B (n_55_87), .C1 (n_59_85), .C2 (n_63_84) );
AOI211_X1 g_58_88 (.ZN (n_58_88), .A (n_54_90), .B (n_53_88), .C1 (n_57_86), .C2 (n_62_86) );
AOI211_X1 g_60_87 (.ZN (n_60_87), .A (n_56_89), .B (n_51_89), .C1 (n_55_87), .C2 (n_61_84) );
AOI211_X1 g_59_89 (.ZN (n_59_89), .A (n_58_88), .B (n_52_91), .C1 (n_53_88), .C2 (n_59_85) );
AOI211_X1 g_58_87 (.ZN (n_58_87), .A (n_60_87), .B (n_54_90), .C1 (n_51_89), .C2 (n_57_86) );
AOI211_X1 g_60_86 (.ZN (n_60_86), .A (n_59_89), .B (n_56_89), .C1 (n_52_91), .C2 (n_55_87) );
AOI211_X1 g_62_85 (.ZN (n_62_85), .A (n_58_87), .B (n_58_88), .C1 (n_54_90), .C2 (n_53_88) );
AOI211_X1 g_61_87 (.ZN (n_61_87), .A (n_60_86), .B (n_60_87), .C1 (n_56_89), .C2 (n_51_89) );
AOI211_X1 g_63_86 (.ZN (n_63_86), .A (n_62_85), .B (n_59_89), .C1 (n_58_88), .C2 (n_52_91) );
AOI211_X1 g_65_85 (.ZN (n_65_85), .A (n_61_87), .B (n_58_87), .C1 (n_60_87), .C2 (n_54_90) );
AOI211_X1 g_67_84 (.ZN (n_67_84), .A (n_63_86), .B (n_60_86), .C1 (n_59_89), .C2 (n_56_89) );
AOI211_X1 g_69_83 (.ZN (n_69_83), .A (n_65_85), .B (n_62_85), .C1 (n_58_87), .C2 (n_58_88) );
AOI211_X1 g_71_82 (.ZN (n_71_82), .A (n_67_84), .B (n_61_87), .C1 (n_60_86), .C2 (n_60_87) );
AOI211_X1 g_73_81 (.ZN (n_73_81), .A (n_69_83), .B (n_63_86), .C1 (n_62_85), .C2 (n_59_89) );
AOI211_X1 g_75_80 (.ZN (n_75_80), .A (n_71_82), .B (n_65_85), .C1 (n_61_87), .C2 (n_58_87) );
AOI211_X1 g_77_79 (.ZN (n_77_79), .A (n_73_81), .B (n_67_84), .C1 (n_63_86), .C2 (n_60_86) );
AOI211_X1 g_76_81 (.ZN (n_76_81), .A (n_75_80), .B (n_69_83), .C1 (n_65_85), .C2 (n_62_85) );
AOI211_X1 g_78_80 (.ZN (n_78_80), .A (n_77_79), .B (n_71_82), .C1 (n_67_84), .C2 (n_61_87) );
AOI211_X1 g_80_79 (.ZN (n_80_79), .A (n_76_81), .B (n_73_81), .C1 (n_69_83), .C2 (n_63_86) );
AOI211_X1 g_82_78 (.ZN (n_82_78), .A (n_78_80), .B (n_75_80), .C1 (n_71_82), .C2 (n_65_85) );
AOI211_X1 g_84_77 (.ZN (n_84_77), .A (n_80_79), .B (n_77_79), .C1 (n_73_81), .C2 (n_67_84) );
AOI211_X1 g_86_76 (.ZN (n_86_76), .A (n_82_78), .B (n_76_81), .C1 (n_75_80), .C2 (n_69_83) );
AOI211_X1 g_88_77 (.ZN (n_88_77), .A (n_84_77), .B (n_78_80), .C1 (n_77_79), .C2 (n_71_82) );
AOI211_X1 g_86_78 (.ZN (n_86_78), .A (n_86_76), .B (n_80_79), .C1 (n_76_81), .C2 (n_73_81) );
AOI211_X1 g_84_79 (.ZN (n_84_79), .A (n_88_77), .B (n_82_78), .C1 (n_78_80), .C2 (n_75_80) );
AOI211_X1 g_83_77 (.ZN (n_83_77), .A (n_86_78), .B (n_84_77), .C1 (n_80_79), .C2 (n_77_79) );
AOI211_X1 g_81_78 (.ZN (n_81_78), .A (n_84_79), .B (n_86_76), .C1 (n_82_78), .C2 (n_76_81) );
AOI211_X1 g_79_79 (.ZN (n_79_79), .A (n_83_77), .B (n_88_77), .C1 (n_84_77), .C2 (n_78_80) );
AOI211_X1 g_77_80 (.ZN (n_77_80), .A (n_81_78), .B (n_86_78), .C1 (n_86_76), .C2 (n_80_79) );
AOI211_X1 g_75_81 (.ZN (n_75_81), .A (n_79_79), .B (n_84_79), .C1 (n_88_77), .C2 (n_82_78) );
AOI211_X1 g_73_82 (.ZN (n_73_82), .A (n_77_80), .B (n_83_77), .C1 (n_86_78), .C2 (n_84_77) );
AOI211_X1 g_71_83 (.ZN (n_71_83), .A (n_75_81), .B (n_81_78), .C1 (n_84_79), .C2 (n_86_76) );
AOI211_X1 g_69_82 (.ZN (n_69_82), .A (n_73_82), .B (n_79_79), .C1 (n_83_77), .C2 (n_88_77) );
AOI211_X1 g_67_83 (.ZN (n_67_83), .A (n_71_83), .B (n_77_80), .C1 (n_81_78), .C2 (n_86_78) );
AOI211_X1 g_65_84 (.ZN (n_65_84), .A (n_69_82), .B (n_75_81), .C1 (n_79_79), .C2 (n_84_79) );
AOI211_X1 g_63_85 (.ZN (n_63_85), .A (n_67_83), .B (n_73_82), .C1 (n_77_80), .C2 (n_83_77) );
AOI211_X1 g_61_86 (.ZN (n_61_86), .A (n_65_84), .B (n_71_83), .C1 (n_75_81), .C2 (n_81_78) );
AOI211_X1 g_59_87 (.ZN (n_59_87), .A (n_63_85), .B (n_69_82), .C1 (n_73_82), .C2 (n_79_79) );
AOI211_X1 g_57_88 (.ZN (n_57_88), .A (n_61_86), .B (n_67_83), .C1 (n_71_83), .C2 (n_77_80) );
AOI211_X1 g_55_89 (.ZN (n_55_89), .A (n_59_87), .B (n_65_84), .C1 (n_69_82), .C2 (n_75_81) );
AOI211_X1 g_53_90 (.ZN (n_53_90), .A (n_57_88), .B (n_63_85), .C1 (n_67_83), .C2 (n_73_82) );
AOI211_X1 g_51_91 (.ZN (n_51_91), .A (n_55_89), .B (n_61_86), .C1 (n_65_84), .C2 (n_71_83) );
AOI211_X1 g_50_89 (.ZN (n_50_89), .A (n_53_90), .B (n_59_87), .C1 (n_63_85), .C2 (n_69_82) );
AOI211_X1 g_49_91 (.ZN (n_49_91), .A (n_51_91), .B (n_57_88), .C1 (n_61_86), .C2 (n_67_83) );
AOI211_X1 g_47_92 (.ZN (n_47_92), .A (n_50_89), .B (n_55_89), .C1 (n_59_87), .C2 (n_65_84) );
AOI211_X1 g_48_90 (.ZN (n_48_90), .A (n_49_91), .B (n_53_90), .C1 (n_57_88), .C2 (n_63_85) );
AOI211_X1 g_46_91 (.ZN (n_46_91), .A (n_47_92), .B (n_51_91), .C1 (n_55_89), .C2 (n_61_86) );
AOI211_X1 g_44_92 (.ZN (n_44_92), .A (n_48_90), .B (n_50_89), .C1 (n_53_90), .C2 (n_59_87) );
AOI211_X1 g_43_94 (.ZN (n_43_94), .A (n_46_91), .B (n_49_91), .C1 (n_51_91), .C2 (n_57_88) );
AOI211_X1 g_45_93 (.ZN (n_45_93), .A (n_44_92), .B (n_47_92), .C1 (n_50_89), .C2 (n_55_89) );
AOI211_X1 g_46_95 (.ZN (n_46_95), .A (n_43_94), .B (n_48_90), .C1 (n_49_91), .C2 (n_53_90) );
AOI211_X1 g_44_96 (.ZN (n_44_96), .A (n_45_93), .B (n_46_91), .C1 (n_47_92), .C2 (n_51_91) );
AOI211_X1 g_45_94 (.ZN (n_45_94), .A (n_46_95), .B (n_44_92), .C1 (n_48_90), .C2 (n_50_89) );
AOI211_X1 g_47_93 (.ZN (n_47_93), .A (n_44_96), .B (n_43_94), .C1 (n_46_91), .C2 (n_49_91) );
AOI211_X1 g_49_92 (.ZN (n_49_92), .A (n_45_94), .B (n_45_93), .C1 (n_44_92), .C2 (n_47_92) );
AOI211_X1 g_48_94 (.ZN (n_48_94), .A (n_47_93), .B (n_46_95), .C1 (n_43_94), .C2 (n_48_90) );
AOI211_X1 g_46_93 (.ZN (n_46_93), .A (n_49_92), .B (n_44_96), .C1 (n_45_93), .C2 (n_46_91) );
AOI211_X1 g_45_95 (.ZN (n_45_95), .A (n_48_94), .B (n_45_94), .C1 (n_46_95), .C2 (n_44_92) );
AOI211_X1 g_46_97 (.ZN (n_46_97), .A (n_46_93), .B (n_47_93), .C1 (n_44_96), .C2 (n_43_94) );
AOI211_X1 g_47_95 (.ZN (n_47_95), .A (n_45_95), .B (n_49_92), .C1 (n_45_94), .C2 (n_45_93) );
AOI211_X1 g_49_94 (.ZN (n_49_94), .A (n_46_97), .B (n_48_94), .C1 (n_47_93), .C2 (n_46_95) );
AOI211_X1 g_48_92 (.ZN (n_48_92), .A (n_47_95), .B (n_46_93), .C1 (n_49_92), .C2 (n_44_96) );
AOI211_X1 g_50_91 (.ZN (n_50_91), .A (n_49_94), .B (n_45_95), .C1 (n_48_94), .C2 (n_45_94) );
AOI211_X1 g_52_90 (.ZN (n_52_90), .A (n_48_92), .B (n_46_97), .C1 (n_46_93), .C2 (n_47_93) );
AOI211_X1 g_54_89 (.ZN (n_54_89), .A (n_50_91), .B (n_47_95), .C1 (n_45_95), .C2 (n_49_92) );
AOI211_X1 g_56_88 (.ZN (n_56_88), .A (n_52_90), .B (n_49_94), .C1 (n_46_97), .C2 (n_48_94) );
AOI211_X1 g_57_90 (.ZN (n_57_90), .A (n_54_89), .B (n_48_92), .C1 (n_47_95), .C2 (n_46_93) );
AOI211_X1 g_55_91 (.ZN (n_55_91), .A (n_56_88), .B (n_50_91), .C1 (n_49_94), .C2 (n_45_95) );
AOI211_X1 g_53_92 (.ZN (n_53_92), .A (n_57_90), .B (n_52_90), .C1 (n_48_92), .C2 (n_46_97) );
AOI211_X1 g_51_93 (.ZN (n_51_93), .A (n_55_91), .B (n_54_89), .C1 (n_50_91), .C2 (n_47_95) );
AOI211_X1 g_50_95 (.ZN (n_50_95), .A (n_53_92), .B (n_56_88), .C1 (n_52_90), .C2 (n_49_94) );
AOI211_X1 g_48_96 (.ZN (n_48_96), .A (n_51_93), .B (n_57_90), .C1 (n_54_89), .C2 (n_48_92) );
AOI211_X1 g_47_94 (.ZN (n_47_94), .A (n_50_95), .B (n_55_91), .C1 (n_56_88), .C2 (n_50_91) );
AOI211_X1 g_49_93 (.ZN (n_49_93), .A (n_48_96), .B (n_53_92), .C1 (n_57_90), .C2 (n_52_90) );
AOI211_X1 g_51_92 (.ZN (n_51_92), .A (n_47_94), .B (n_51_93), .C1 (n_55_91), .C2 (n_54_89) );
AOI211_X1 g_53_91 (.ZN (n_53_91), .A (n_49_93), .B (n_50_95), .C1 (n_53_92), .C2 (n_56_88) );
AOI211_X1 g_55_90 (.ZN (n_55_90), .A (n_51_92), .B (n_48_96), .C1 (n_51_93), .C2 (n_57_90) );
AOI211_X1 g_57_89 (.ZN (n_57_89), .A (n_53_91), .B (n_47_94), .C1 (n_50_95), .C2 (n_55_91) );
AOI211_X1 g_59_88 (.ZN (n_59_88), .A (n_55_90), .B (n_49_93), .C1 (n_48_96), .C2 (n_53_92) );
AOI211_X1 g_58_90 (.ZN (n_58_90), .A (n_57_89), .B (n_51_92), .C1 (n_47_94), .C2 (n_51_93) );
AOI211_X1 g_60_89 (.ZN (n_60_89), .A (n_59_88), .B (n_53_91), .C1 (n_49_93), .C2 (n_50_95) );
AOI211_X1 g_62_88 (.ZN (n_62_88), .A (n_58_90), .B (n_55_90), .C1 (n_51_92), .C2 (n_48_96) );
AOI211_X1 g_64_87 (.ZN (n_64_87), .A (n_60_89), .B (n_57_89), .C1 (n_53_91), .C2 (n_47_94) );
AOI211_X1 g_66_86 (.ZN (n_66_86), .A (n_62_88), .B (n_59_88), .C1 (n_55_90), .C2 (n_49_93) );
AOI211_X1 g_68_85 (.ZN (n_68_85), .A (n_64_87), .B (n_58_90), .C1 (n_57_89), .C2 (n_51_92) );
AOI211_X1 g_70_84 (.ZN (n_70_84), .A (n_66_86), .B (n_60_89), .C1 (n_59_88), .C2 (n_53_91) );
AOI211_X1 g_72_83 (.ZN (n_72_83), .A (n_68_85), .B (n_62_88), .C1 (n_58_90), .C2 (n_55_90) );
AOI211_X1 g_74_82 (.ZN (n_74_82), .A (n_70_84), .B (n_64_87), .C1 (n_60_89), .C2 (n_57_89) );
AOI211_X1 g_73_84 (.ZN (n_73_84), .A (n_72_83), .B (n_66_86), .C1 (n_62_88), .C2 (n_59_88) );
AOI211_X1 g_72_82 (.ZN (n_72_82), .A (n_74_82), .B (n_68_85), .C1 (n_64_87), .C2 (n_58_90) );
AOI211_X1 g_74_81 (.ZN (n_74_81), .A (n_73_84), .B (n_70_84), .C1 (n_66_86), .C2 (n_60_89) );
AOI211_X1 g_76_80 (.ZN (n_76_80), .A (n_72_82), .B (n_72_83), .C1 (n_68_85), .C2 (n_62_88) );
AOI211_X1 g_78_79 (.ZN (n_78_79), .A (n_74_81), .B (n_74_82), .C1 (n_70_84), .C2 (n_64_87) );
AOI211_X1 g_80_78 (.ZN (n_80_78), .A (n_76_80), .B (n_73_84), .C1 (n_72_83), .C2 (n_66_86) );
AOI211_X1 g_82_77 (.ZN (n_82_77), .A (n_78_79), .B (n_72_82), .C1 (n_74_82), .C2 (n_68_85) );
AOI211_X1 g_84_76 (.ZN (n_84_76), .A (n_80_78), .B (n_74_81), .C1 (n_73_84), .C2 (n_70_84) );
AOI211_X1 g_83_78 (.ZN (n_83_78), .A (n_82_77), .B (n_76_80), .C1 (n_72_82), .C2 (n_72_83) );
AOI211_X1 g_81_79 (.ZN (n_81_79), .A (n_84_76), .B (n_78_79), .C1 (n_74_81), .C2 (n_74_82) );
AOI211_X1 g_79_80 (.ZN (n_79_80), .A (n_83_78), .B (n_80_78), .C1 (n_76_80), .C2 (n_73_84) );
AOI211_X1 g_77_81 (.ZN (n_77_81), .A (n_81_79), .B (n_82_77), .C1 (n_78_79), .C2 (n_72_82) );
AOI211_X1 g_75_82 (.ZN (n_75_82), .A (n_79_80), .B (n_84_76), .C1 (n_80_78), .C2 (n_74_81) );
AOI211_X1 g_73_83 (.ZN (n_73_83), .A (n_77_81), .B (n_83_78), .C1 (n_82_77), .C2 (n_76_80) );
AOI211_X1 g_71_84 (.ZN (n_71_84), .A (n_75_82), .B (n_81_79), .C1 (n_84_76), .C2 (n_78_79) );
AOI211_X1 g_69_85 (.ZN (n_69_85), .A (n_73_83), .B (n_79_80), .C1 (n_83_78), .C2 (n_80_78) );
AOI211_X1 g_70_83 (.ZN (n_70_83), .A (n_71_84), .B (n_77_81), .C1 (n_81_79), .C2 (n_82_77) );
AOI211_X1 g_68_84 (.ZN (n_68_84), .A (n_69_85), .B (n_75_82), .C1 (n_79_80), .C2 (n_84_76) );
AOI211_X1 g_66_85 (.ZN (n_66_85), .A (n_70_83), .B (n_73_83), .C1 (n_77_81), .C2 (n_83_78) );
AOI211_X1 g_64_86 (.ZN (n_64_86), .A (n_68_84), .B (n_71_84), .C1 (n_75_82), .C2 (n_81_79) );
AOI211_X1 g_62_87 (.ZN (n_62_87), .A (n_66_85), .B (n_69_85), .C1 (n_73_83), .C2 (n_79_80) );
AOI211_X1 g_60_88 (.ZN (n_60_88), .A (n_64_86), .B (n_70_83), .C1 (n_71_84), .C2 (n_77_81) );
AOI211_X1 g_58_89 (.ZN (n_58_89), .A (n_62_87), .B (n_68_84), .C1 (n_69_85), .C2 (n_75_82) );
AOI211_X1 g_56_90 (.ZN (n_56_90), .A (n_60_88), .B (n_66_85), .C1 (n_70_83), .C2 (n_73_83) );
AOI211_X1 g_54_91 (.ZN (n_54_91), .A (n_58_89), .B (n_64_86), .C1 (n_68_84), .C2 (n_71_84) );
AOI211_X1 g_52_92 (.ZN (n_52_92), .A (n_56_90), .B (n_62_87), .C1 (n_66_85), .C2 (n_69_85) );
AOI211_X1 g_50_93 (.ZN (n_50_93), .A (n_54_91), .B (n_60_88), .C1 (n_64_86), .C2 (n_70_83) );
AOI211_X1 g_49_95 (.ZN (n_49_95), .A (n_52_92), .B (n_58_89), .C1 (n_62_87), .C2 (n_68_84) );
AOI211_X1 g_51_94 (.ZN (n_51_94), .A (n_50_93), .B (n_56_90), .C1 (n_60_88), .C2 (n_66_85) );
AOI211_X1 g_53_93 (.ZN (n_53_93), .A (n_49_95), .B (n_54_91), .C1 (n_58_89), .C2 (n_64_86) );
AOI211_X1 g_55_92 (.ZN (n_55_92), .A (n_51_94), .B (n_52_92), .C1 (n_56_90), .C2 (n_62_87) );
AOI211_X1 g_57_91 (.ZN (n_57_91), .A (n_53_93), .B (n_50_93), .C1 (n_54_91), .C2 (n_60_88) );
AOI211_X1 g_59_90 (.ZN (n_59_90), .A (n_55_92), .B (n_49_95), .C1 (n_52_92), .C2 (n_58_89) );
AOI211_X1 g_61_89 (.ZN (n_61_89), .A (n_57_91), .B (n_51_94), .C1 (n_50_93), .C2 (n_56_90) );
AOI211_X1 g_63_88 (.ZN (n_63_88), .A (n_59_90), .B (n_53_93), .C1 (n_49_95), .C2 (n_54_91) );
AOI211_X1 g_65_87 (.ZN (n_65_87), .A (n_61_89), .B (n_55_92), .C1 (n_51_94), .C2 (n_52_92) );
AOI211_X1 g_67_86 (.ZN (n_67_86), .A (n_63_88), .B (n_57_91), .C1 (n_53_93), .C2 (n_50_93) );
AOI211_X1 g_66_88 (.ZN (n_66_88), .A (n_65_87), .B (n_59_90), .C1 (n_55_92), .C2 (n_49_95) );
AOI211_X1 g_65_86 (.ZN (n_65_86), .A (n_67_86), .B (n_61_89), .C1 (n_57_91), .C2 (n_51_94) );
AOI211_X1 g_63_87 (.ZN (n_63_87), .A (n_66_88), .B (n_63_88), .C1 (n_59_90), .C2 (n_53_93) );
AOI211_X1 g_61_88 (.ZN (n_61_88), .A (n_65_86), .B (n_65_87), .C1 (n_61_89), .C2 (n_55_92) );
AOI211_X1 g_60_90 (.ZN (n_60_90), .A (n_63_87), .B (n_67_86), .C1 (n_63_88), .C2 (n_57_91) );
AOI211_X1 g_62_89 (.ZN (n_62_89), .A (n_61_88), .B (n_66_88), .C1 (n_65_87), .C2 (n_59_90) );
AOI211_X1 g_64_88 (.ZN (n_64_88), .A (n_60_90), .B (n_65_86), .C1 (n_67_86), .C2 (n_61_89) );
AOI211_X1 g_66_87 (.ZN (n_66_87), .A (n_62_89), .B (n_63_87), .C1 (n_66_88), .C2 (n_63_88) );
AOI211_X1 g_68_86 (.ZN (n_68_86), .A (n_64_88), .B (n_61_88), .C1 (n_65_86), .C2 (n_65_87) );
AOI211_X1 g_69_84 (.ZN (n_69_84), .A (n_66_87), .B (n_60_90), .C1 (n_63_87), .C2 (n_67_86) );
AOI211_X1 g_71_85 (.ZN (n_71_85), .A (n_68_86), .B (n_62_89), .C1 (n_61_88), .C2 (n_66_88) );
AOI211_X1 g_69_86 (.ZN (n_69_86), .A (n_69_84), .B (n_64_88), .C1 (n_60_90), .C2 (n_65_86) );
AOI211_X1 g_67_87 (.ZN (n_67_87), .A (n_71_85), .B (n_66_87), .C1 (n_62_89), .C2 (n_63_87) );
AOI211_X1 g_65_88 (.ZN (n_65_88), .A (n_69_86), .B (n_68_86), .C1 (n_64_88), .C2 (n_61_88) );
AOI211_X1 g_63_89 (.ZN (n_63_89), .A (n_67_87), .B (n_69_84), .C1 (n_66_87), .C2 (n_60_90) );
AOI211_X1 g_61_90 (.ZN (n_61_90), .A (n_65_88), .B (n_71_85), .C1 (n_68_86), .C2 (n_62_89) );
AOI211_X1 g_59_91 (.ZN (n_59_91), .A (n_63_89), .B (n_69_86), .C1 (n_69_84), .C2 (n_64_88) );
AOI211_X1 g_57_92 (.ZN (n_57_92), .A (n_61_90), .B (n_67_87), .C1 (n_71_85), .C2 (n_66_87) );
AOI211_X1 g_55_93 (.ZN (n_55_93), .A (n_59_91), .B (n_65_88), .C1 (n_69_86), .C2 (n_68_86) );
AOI211_X1 g_56_91 (.ZN (n_56_91), .A (n_57_92), .B (n_63_89), .C1 (n_67_87), .C2 (n_69_84) );
AOI211_X1 g_54_92 (.ZN (n_54_92), .A (n_55_93), .B (n_61_90), .C1 (n_65_88), .C2 (n_71_85) );
AOI211_X1 g_52_93 (.ZN (n_52_93), .A (n_56_91), .B (n_59_91), .C1 (n_63_89), .C2 (n_69_86) );
AOI211_X1 g_50_94 (.ZN (n_50_94), .A (n_54_92), .B (n_57_92), .C1 (n_61_90), .C2 (n_67_87) );
AOI211_X1 g_48_95 (.ZN (n_48_95), .A (n_52_93), .B (n_55_93), .C1 (n_59_91), .C2 (n_65_88) );
AOI211_X1 g_46_96 (.ZN (n_46_96), .A (n_50_94), .B (n_56_91), .C1 (n_57_92), .C2 (n_63_89) );
AOI211_X1 g_45_98 (.ZN (n_45_98), .A (n_48_95), .B (n_54_92), .C1 (n_55_93), .C2 (n_61_90) );
AOI211_X1 g_47_97 (.ZN (n_47_97), .A (n_46_96), .B (n_52_93), .C1 (n_56_91), .C2 (n_59_91) );
AOI211_X1 g_49_96 (.ZN (n_49_96), .A (n_45_98), .B (n_50_94), .C1 (n_54_92), .C2 (n_57_92) );
AOI211_X1 g_48_98 (.ZN (n_48_98), .A (n_47_97), .B (n_48_95), .C1 (n_52_93), .C2 (n_55_93) );
AOI211_X1 g_49_100 (.ZN (n_49_100), .A (n_49_96), .B (n_46_96), .C1 (n_50_94), .C2 (n_56_91) );
AOI211_X1 g_47_99 (.ZN (n_47_99), .A (n_48_98), .B (n_45_98), .C1 (n_48_95), .C2 (n_54_92) );
AOI211_X1 g_48_97 (.ZN (n_48_97), .A (n_49_100), .B (n_47_97), .C1 (n_46_96), .C2 (n_52_93) );
AOI211_X1 g_50_98 (.ZN (n_50_98), .A (n_47_99), .B (n_49_96), .C1 (n_45_98), .C2 (n_50_94) );
AOI211_X1 g_51_96 (.ZN (n_51_96), .A (n_48_97), .B (n_48_98), .C1 (n_47_97), .C2 (n_48_95) );
AOI211_X1 g_52_94 (.ZN (n_52_94), .A (n_50_98), .B (n_49_100), .C1 (n_49_96), .C2 (n_46_96) );
AOI211_X1 g_54_93 (.ZN (n_54_93), .A (n_51_96), .B (n_47_99), .C1 (n_48_98), .C2 (n_45_98) );
AOI211_X1 g_56_92 (.ZN (n_56_92), .A (n_52_94), .B (n_48_97), .C1 (n_49_100), .C2 (n_47_97) );
AOI211_X1 g_58_91 (.ZN (n_58_91), .A (n_54_93), .B (n_50_98), .C1 (n_47_99), .C2 (n_49_96) );
AOI211_X1 g_57_93 (.ZN (n_57_93), .A (n_56_92), .B (n_51_96), .C1 (n_48_97), .C2 (n_48_98) );
AOI211_X1 g_59_92 (.ZN (n_59_92), .A (n_58_91), .B (n_52_94), .C1 (n_50_98), .C2 (n_49_100) );
AOI211_X1 g_61_91 (.ZN (n_61_91), .A (n_57_93), .B (n_54_93), .C1 (n_51_96), .C2 (n_47_99) );
AOI211_X1 g_63_90 (.ZN (n_63_90), .A (n_59_92), .B (n_56_92), .C1 (n_52_94), .C2 (n_48_97) );
AOI211_X1 g_65_89 (.ZN (n_65_89), .A (n_61_91), .B (n_58_91), .C1 (n_54_93), .C2 (n_50_98) );
AOI211_X1 g_67_88 (.ZN (n_67_88), .A (n_63_90), .B (n_57_93), .C1 (n_56_92), .C2 (n_51_96) );
AOI211_X1 g_69_87 (.ZN (n_69_87), .A (n_65_89), .B (n_59_92), .C1 (n_58_91), .C2 (n_52_94) );
AOI211_X1 g_70_85 (.ZN (n_70_85), .A (n_67_88), .B (n_61_91), .C1 (n_57_93), .C2 (n_54_93) );
AOI211_X1 g_72_84 (.ZN (n_72_84), .A (n_69_87), .B (n_63_90), .C1 (n_59_92), .C2 (n_56_92) );
AOI211_X1 g_74_83 (.ZN (n_74_83), .A (n_70_85), .B (n_65_89), .C1 (n_61_91), .C2 (n_58_91) );
AOI211_X1 g_76_82 (.ZN (n_76_82), .A (n_72_84), .B (n_67_88), .C1 (n_63_90), .C2 (n_57_93) );
AOI211_X1 g_78_81 (.ZN (n_78_81), .A (n_74_83), .B (n_69_87), .C1 (n_65_89), .C2 (n_59_92) );
AOI211_X1 g_80_80 (.ZN (n_80_80), .A (n_76_82), .B (n_70_85), .C1 (n_67_88), .C2 (n_61_91) );
AOI211_X1 g_82_79 (.ZN (n_82_79), .A (n_78_81), .B (n_72_84), .C1 (n_69_87), .C2 (n_63_90) );
AOI211_X1 g_84_78 (.ZN (n_84_78), .A (n_80_80), .B (n_74_83), .C1 (n_70_85), .C2 (n_65_89) );
AOI211_X1 g_86_77 (.ZN (n_86_77), .A (n_82_79), .B (n_76_82), .C1 (n_72_84), .C2 (n_67_88) );
AOI211_X1 g_88_76 (.ZN (n_88_76), .A (n_84_78), .B (n_78_81), .C1 (n_74_83), .C2 (n_69_87) );
AOI211_X1 g_90_75 (.ZN (n_90_75), .A (n_86_77), .B (n_80_80), .C1 (n_76_82), .C2 (n_70_85) );
AOI211_X1 g_92_74 (.ZN (n_92_74), .A (n_88_76), .B (n_82_79), .C1 (n_78_81), .C2 (n_72_84) );
AOI211_X1 g_91_76 (.ZN (n_91_76), .A (n_90_75), .B (n_84_78), .C1 (n_80_80), .C2 (n_74_83) );
AOI211_X1 g_89_77 (.ZN (n_89_77), .A (n_92_74), .B (n_86_77), .C1 (n_82_79), .C2 (n_76_82) );
AOI211_X1 g_87_78 (.ZN (n_87_78), .A (n_91_76), .B (n_88_76), .C1 (n_84_78), .C2 (n_78_81) );
AOI211_X1 g_85_79 (.ZN (n_85_79), .A (n_89_77), .B (n_90_75), .C1 (n_86_77), .C2 (n_80_80) );
AOI211_X1 g_83_80 (.ZN (n_83_80), .A (n_87_78), .B (n_92_74), .C1 (n_88_76), .C2 (n_82_79) );
AOI211_X1 g_81_81 (.ZN (n_81_81), .A (n_85_79), .B (n_91_76), .C1 (n_90_75), .C2 (n_84_78) );
AOI211_X1 g_79_82 (.ZN (n_79_82), .A (n_83_80), .B (n_89_77), .C1 (n_92_74), .C2 (n_86_77) );
AOI211_X1 g_77_83 (.ZN (n_77_83), .A (n_81_81), .B (n_87_78), .C1 (n_91_76), .C2 (n_88_76) );
AOI211_X1 g_75_84 (.ZN (n_75_84), .A (n_79_82), .B (n_85_79), .C1 (n_89_77), .C2 (n_90_75) );
AOI211_X1 g_73_85 (.ZN (n_73_85), .A (n_77_83), .B (n_83_80), .C1 (n_87_78), .C2 (n_92_74) );
AOI211_X1 g_71_86 (.ZN (n_71_86), .A (n_75_84), .B (n_81_81), .C1 (n_85_79), .C2 (n_91_76) );
AOI211_X1 g_70_88 (.ZN (n_70_88), .A (n_73_85), .B (n_79_82), .C1 (n_83_80), .C2 (n_89_77) );
AOI211_X1 g_68_87 (.ZN (n_68_87), .A (n_71_86), .B (n_77_83), .C1 (n_81_81), .C2 (n_87_78) );
AOI211_X1 g_70_86 (.ZN (n_70_86), .A (n_70_88), .B (n_75_84), .C1 (n_79_82), .C2 (n_85_79) );
AOI211_X1 g_72_85 (.ZN (n_72_85), .A (n_68_87), .B (n_73_85), .C1 (n_77_83), .C2 (n_83_80) );
AOI211_X1 g_74_84 (.ZN (n_74_84), .A (n_70_86), .B (n_71_86), .C1 (n_75_84), .C2 (n_81_81) );
AOI211_X1 g_76_83 (.ZN (n_76_83), .A (n_72_85), .B (n_70_88), .C1 (n_73_85), .C2 (n_79_82) );
AOI211_X1 g_78_82 (.ZN (n_78_82), .A (n_74_84), .B (n_68_87), .C1 (n_71_86), .C2 (n_77_83) );
AOI211_X1 g_80_81 (.ZN (n_80_81), .A (n_76_83), .B (n_70_86), .C1 (n_70_88), .C2 (n_75_84) );
AOI211_X1 g_82_80 (.ZN (n_82_80), .A (n_78_82), .B (n_72_85), .C1 (n_68_87), .C2 (n_73_85) );
AOI211_X1 g_81_82 (.ZN (n_81_82), .A (n_80_81), .B (n_74_84), .C1 (n_70_86), .C2 (n_71_86) );
AOI211_X1 g_79_81 (.ZN (n_79_81), .A (n_82_80), .B (n_76_83), .C1 (n_72_85), .C2 (n_70_88) );
AOI211_X1 g_81_80 (.ZN (n_81_80), .A (n_81_82), .B (n_78_82), .C1 (n_74_84), .C2 (n_68_87) );
AOI211_X1 g_83_79 (.ZN (n_83_79), .A (n_79_81), .B (n_80_81), .C1 (n_76_83), .C2 (n_70_86) );
AOI211_X1 g_85_78 (.ZN (n_85_78), .A (n_81_80), .B (n_82_80), .C1 (n_78_82), .C2 (n_72_85) );
AOI211_X1 g_84_80 (.ZN (n_84_80), .A (n_83_79), .B (n_81_82), .C1 (n_80_81), .C2 (n_74_84) );
AOI211_X1 g_86_79 (.ZN (n_86_79), .A (n_85_78), .B (n_79_81), .C1 (n_82_80), .C2 (n_76_83) );
AOI211_X1 g_88_78 (.ZN (n_88_78), .A (n_84_80), .B (n_81_80), .C1 (n_81_82), .C2 (n_78_82) );
AOI211_X1 g_90_77 (.ZN (n_90_77), .A (n_86_79), .B (n_83_79), .C1 (n_79_81), .C2 (n_80_81) );
AOI211_X1 g_92_76 (.ZN (n_92_76), .A (n_88_78), .B (n_85_78), .C1 (n_81_80), .C2 (n_82_80) );
AOI211_X1 g_94_75 (.ZN (n_94_75), .A (n_90_77), .B (n_84_80), .C1 (n_83_79), .C2 (n_81_82) );
AOI211_X1 g_93_77 (.ZN (n_93_77), .A (n_92_76), .B (n_86_79), .C1 (n_85_78), .C2 (n_79_81) );
AOI211_X1 g_91_78 (.ZN (n_91_78), .A (n_94_75), .B (n_88_78), .C1 (n_84_80), .C2 (n_81_80) );
AOI211_X1 g_89_79 (.ZN (n_89_79), .A (n_93_77), .B (n_90_77), .C1 (n_86_79), .C2 (n_83_79) );
AOI211_X1 g_87_80 (.ZN (n_87_80), .A (n_91_78), .B (n_92_76), .C1 (n_88_78), .C2 (n_85_78) );
AOI211_X1 g_85_81 (.ZN (n_85_81), .A (n_89_79), .B (n_94_75), .C1 (n_90_77), .C2 (n_84_80) );
AOI211_X1 g_83_82 (.ZN (n_83_82), .A (n_87_80), .B (n_93_77), .C1 (n_92_76), .C2 (n_86_79) );
AOI211_X1 g_81_83 (.ZN (n_81_83), .A (n_85_81), .B (n_91_78), .C1 (n_94_75), .C2 (n_88_78) );
AOI211_X1 g_82_81 (.ZN (n_82_81), .A (n_83_82), .B (n_89_79), .C1 (n_93_77), .C2 (n_90_77) );
AOI211_X1 g_80_82 (.ZN (n_80_82), .A (n_81_83), .B (n_87_80), .C1 (n_91_78), .C2 (n_92_76) );
AOI211_X1 g_78_83 (.ZN (n_78_83), .A (n_82_81), .B (n_85_81), .C1 (n_89_79), .C2 (n_94_75) );
AOI211_X1 g_76_84 (.ZN (n_76_84), .A (n_80_82), .B (n_83_82), .C1 (n_87_80), .C2 (n_93_77) );
AOI211_X1 g_77_82 (.ZN (n_77_82), .A (n_78_83), .B (n_81_83), .C1 (n_85_81), .C2 (n_91_78) );
AOI211_X1 g_75_83 (.ZN (n_75_83), .A (n_76_84), .B (n_82_81), .C1 (n_83_82), .C2 (n_89_79) );
AOI211_X1 g_74_85 (.ZN (n_74_85), .A (n_77_82), .B (n_80_82), .C1 (n_81_83), .C2 (n_87_80) );
AOI211_X1 g_72_86 (.ZN (n_72_86), .A (n_75_83), .B (n_78_83), .C1 (n_82_81), .C2 (n_85_81) );
AOI211_X1 g_70_87 (.ZN (n_70_87), .A (n_74_85), .B (n_76_84), .C1 (n_80_82), .C2 (n_83_82) );
AOI211_X1 g_68_88 (.ZN (n_68_88), .A (n_72_86), .B (n_77_82), .C1 (n_78_83), .C2 (n_81_83) );
AOI211_X1 g_66_89 (.ZN (n_66_89), .A (n_70_87), .B (n_75_83), .C1 (n_76_84), .C2 (n_82_81) );
AOI211_X1 g_64_90 (.ZN (n_64_90), .A (n_68_88), .B (n_74_85), .C1 (n_77_82), .C2 (n_80_82) );
AOI211_X1 g_62_91 (.ZN (n_62_91), .A (n_66_89), .B (n_72_86), .C1 (n_75_83), .C2 (n_78_83) );
AOI211_X1 g_60_92 (.ZN (n_60_92), .A (n_64_90), .B (n_70_87), .C1 (n_74_85), .C2 (n_76_84) );
AOI211_X1 g_58_93 (.ZN (n_58_93), .A (n_62_91), .B (n_68_88), .C1 (n_72_86), .C2 (n_77_82) );
AOI211_X1 g_56_94 (.ZN (n_56_94), .A (n_60_92), .B (n_66_89), .C1 (n_70_87), .C2 (n_75_83) );
AOI211_X1 g_54_95 (.ZN (n_54_95), .A (n_58_93), .B (n_64_90), .C1 (n_68_88), .C2 (n_74_85) );
AOI211_X1 g_52_96 (.ZN (n_52_96), .A (n_56_94), .B (n_62_91), .C1 (n_66_89), .C2 (n_72_86) );
AOI211_X1 g_53_94 (.ZN (n_53_94), .A (n_54_95), .B (n_60_92), .C1 (n_64_90), .C2 (n_70_87) );
AOI211_X1 g_51_95 (.ZN (n_51_95), .A (n_52_96), .B (n_58_93), .C1 (n_62_91), .C2 (n_68_88) );
AOI211_X1 g_50_97 (.ZN (n_50_97), .A (n_53_94), .B (n_56_94), .C1 (n_60_92), .C2 (n_66_89) );
AOI211_X1 g_51_99 (.ZN (n_51_99), .A (n_51_95), .B (n_54_95), .C1 (n_58_93), .C2 (n_64_90) );
AOI211_X1 g_49_98 (.ZN (n_49_98), .A (n_50_97), .B (n_52_96), .C1 (n_56_94), .C2 (n_62_91) );
AOI211_X1 g_50_96 (.ZN (n_50_96), .A (n_51_99), .B (n_53_94), .C1 (n_54_95), .C2 (n_60_92) );
AOI211_X1 g_52_97 (.ZN (n_52_97), .A (n_49_98), .B (n_51_95), .C1 (n_52_96), .C2 (n_58_93) );
AOI211_X1 g_53_95 (.ZN (n_53_95), .A (n_50_96), .B (n_50_97), .C1 (n_53_94), .C2 (n_56_94) );
AOI211_X1 g_55_94 (.ZN (n_55_94), .A (n_52_97), .B (n_51_99), .C1 (n_51_95), .C2 (n_54_95) );
AOI211_X1 g_54_96 (.ZN (n_54_96), .A (n_53_95), .B (n_49_98), .C1 (n_50_97), .C2 (n_52_96) );
AOI211_X1 g_52_95 (.ZN (n_52_95), .A (n_55_94), .B (n_50_96), .C1 (n_51_99), .C2 (n_53_94) );
AOI211_X1 g_51_97 (.ZN (n_51_97), .A (n_54_96), .B (n_52_97), .C1 (n_49_98), .C2 (n_51_95) );
AOI211_X1 g_53_98 (.ZN (n_53_98), .A (n_52_95), .B (n_53_95), .C1 (n_50_96), .C2 (n_50_97) );
AOI211_X1 g_55_97 (.ZN (n_55_97), .A (n_51_97), .B (n_55_94), .C1 (n_52_97), .C2 (n_51_99) );
AOI211_X1 g_56_95 (.ZN (n_56_95), .A (n_53_98), .B (n_54_96), .C1 (n_53_95), .C2 (n_49_98) );
AOI211_X1 g_54_94 (.ZN (n_54_94), .A (n_55_97), .B (n_52_95), .C1 (n_55_94), .C2 (n_50_96) );
AOI211_X1 g_53_96 (.ZN (n_53_96), .A (n_56_95), .B (n_51_97), .C1 (n_54_96), .C2 (n_52_97) );
AOI211_X1 g_52_98 (.ZN (n_52_98), .A (n_54_94), .B (n_53_98), .C1 (n_52_95), .C2 (n_53_95) );
AOI211_X1 g_53_100 (.ZN (n_53_100), .A (n_53_96), .B (n_55_97), .C1 (n_51_97), .C2 (n_55_94) );
AOI211_X1 g_54_98 (.ZN (n_54_98), .A (n_52_98), .B (n_56_95), .C1 (n_53_98), .C2 (n_54_96) );
AOI211_X1 g_55_96 (.ZN (n_55_96), .A (n_53_100), .B (n_54_94), .C1 (n_55_97), .C2 (n_52_95) );
AOI211_X1 g_53_97 (.ZN (n_53_97), .A (n_54_98), .B (n_53_96), .C1 (n_56_95), .C2 (n_51_97) );
AOI211_X1 g_54_99 (.ZN (n_54_99), .A (n_55_96), .B (n_52_98), .C1 (n_54_94), .C2 (n_53_98) );
AOI211_X1 g_56_100 (.ZN (n_56_100), .A (n_53_97), .B (n_53_100), .C1 (n_53_96), .C2 (n_55_97) );
AOI211_X1 g_55_98 (.ZN (n_55_98), .A (n_54_99), .B (n_54_98), .C1 (n_52_98), .C2 (n_56_95) );
AOI211_X1 g_57_97 (.ZN (n_57_97), .A (n_56_100), .B (n_55_96), .C1 (n_53_100), .C2 (n_54_94) );
AOI211_X1 g_58_99 (.ZN (n_58_99), .A (n_55_98), .B (n_53_97), .C1 (n_54_98), .C2 (n_53_96) );
AOI211_X1 g_60_100 (.ZN (n_60_100), .A (n_57_97), .B (n_54_99), .C1 (n_55_96), .C2 (n_52_98) );
AOI211_X1 g_59_98 (.ZN (n_59_98), .A (n_58_99), .B (n_56_100), .C1 (n_53_97), .C2 (n_53_100) );
AOI211_X1 g_61_97 (.ZN (n_61_97), .A (n_60_100), .B (n_55_98), .C1 (n_54_99), .C2 (n_54_98) );
AOI211_X1 g_62_99 (.ZN (n_62_99), .A (n_59_98), .B (n_57_97), .C1 (n_56_100), .C2 (n_55_96) );
AOI211_X1 g_64_100 (.ZN (n_64_100), .A (n_61_97), .B (n_58_99), .C1 (n_55_98), .C2 (n_53_97) );
AOI211_X1 g_63_98 (.ZN (n_63_98), .A (n_62_99), .B (n_60_100), .C1 (n_57_97), .C2 (n_54_99) );
AOI211_X1 g_65_97 (.ZN (n_65_97), .A (n_64_100), .B (n_59_98), .C1 (n_58_99), .C2 (n_56_100) );
AOI211_X1 g_66_99 (.ZN (n_66_99), .A (n_63_98), .B (n_61_97), .C1 (n_60_100), .C2 (n_55_98) );
AOI211_X1 g_68_100 (.ZN (n_68_100), .A (n_65_97), .B (n_62_99), .C1 (n_59_98), .C2 (n_57_97) );
AOI211_X1 g_67_98 (.ZN (n_67_98), .A (n_66_99), .B (n_64_100), .C1 (n_61_97), .C2 (n_58_99) );
AOI211_X1 g_69_97 (.ZN (n_69_97), .A (n_68_100), .B (n_63_98), .C1 (n_62_99), .C2 (n_60_100) );
AOI211_X1 g_70_99 (.ZN (n_70_99), .A (n_67_98), .B (n_65_97), .C1 (n_64_100), .C2 (n_59_98) );
AOI211_X1 g_72_100 (.ZN (n_72_100), .A (n_69_97), .B (n_66_99), .C1 (n_63_98), .C2 (n_61_97) );
AOI211_X1 g_71_98 (.ZN (n_71_98), .A (n_70_99), .B (n_68_100), .C1 (n_65_97), .C2 (n_62_99) );
AOI211_X1 g_73_97 (.ZN (n_73_97), .A (n_72_100), .B (n_67_98), .C1 (n_66_99), .C2 (n_64_100) );
AOI211_X1 g_74_99 (.ZN (n_74_99), .A (n_71_98), .B (n_69_97), .C1 (n_68_100), .C2 (n_63_98) );
AOI211_X1 g_76_100 (.ZN (n_76_100), .A (n_73_97), .B (n_70_99), .C1 (n_67_98), .C2 (n_65_97) );
AOI211_X1 g_75_98 (.ZN (n_75_98), .A (n_74_99), .B (n_72_100), .C1 (n_69_97), .C2 (n_66_99) );
AOI211_X1 g_77_97 (.ZN (n_77_97), .A (n_76_100), .B (n_71_98), .C1 (n_70_99), .C2 (n_68_100) );
AOI211_X1 g_78_99 (.ZN (n_78_99), .A (n_75_98), .B (n_73_97), .C1 (n_72_100), .C2 (n_67_98) );
AOI211_X1 g_80_100 (.ZN (n_80_100), .A (n_77_97), .B (n_74_99), .C1 (n_71_98), .C2 (n_69_97) );
AOI211_X1 g_79_98 (.ZN (n_79_98), .A (n_78_99), .B (n_76_100), .C1 (n_73_97), .C2 (n_70_99) );
AOI211_X1 g_81_97 (.ZN (n_81_97), .A (n_80_100), .B (n_75_98), .C1 (n_74_99), .C2 (n_72_100) );
AOI211_X1 g_82_99 (.ZN (n_82_99), .A (n_79_98), .B (n_77_97), .C1 (n_76_100), .C2 (n_71_98) );
AOI211_X1 g_84_100 (.ZN (n_84_100), .A (n_81_97), .B (n_78_99), .C1 (n_75_98), .C2 (n_73_97) );
AOI211_X1 g_83_98 (.ZN (n_83_98), .A (n_82_99), .B (n_80_100), .C1 (n_77_97), .C2 (n_74_99) );
AOI211_X1 g_85_97 (.ZN (n_85_97), .A (n_84_100), .B (n_79_98), .C1 (n_78_99), .C2 (n_76_100) );
AOI211_X1 g_86_99 (.ZN (n_86_99), .A (n_83_98), .B (n_81_97), .C1 (n_80_100), .C2 (n_75_98) );
AOI211_X1 g_88_100 (.ZN (n_88_100), .A (n_85_97), .B (n_82_99), .C1 (n_79_98), .C2 (n_77_97) );
AOI211_X1 g_87_98 (.ZN (n_87_98), .A (n_86_99), .B (n_84_100), .C1 (n_81_97), .C2 (n_78_99) );
AOI211_X1 g_89_97 (.ZN (n_89_97), .A (n_88_100), .B (n_83_98), .C1 (n_82_99), .C2 (n_80_100) );
AOI211_X1 g_90_99 (.ZN (n_90_99), .A (n_87_98), .B (n_85_97), .C1 (n_84_100), .C2 (n_79_98) );
AOI211_X1 g_92_100 (.ZN (n_92_100), .A (n_89_97), .B (n_86_99), .C1 (n_83_98), .C2 (n_81_97) );
AOI211_X1 g_91_98 (.ZN (n_91_98), .A (n_90_99), .B (n_88_100), .C1 (n_85_97), .C2 (n_82_99) );
AOI211_X1 g_93_97 (.ZN (n_93_97), .A (n_92_100), .B (n_87_98), .C1 (n_86_99), .C2 (n_84_100) );
AOI211_X1 g_94_99 (.ZN (n_94_99), .A (n_91_98), .B (n_89_97), .C1 (n_88_100), .C2 (n_83_98) );
AOI211_X1 g_96_98 (.ZN (n_96_98), .A (n_93_97), .B (n_90_99), .C1 (n_87_98), .C2 (n_85_97) );
AOI211_X1 g_98_97 (.ZN (n_98_97), .A (n_94_99), .B (n_92_100), .C1 (n_89_97), .C2 (n_86_99) );
AOI211_X1 g_99_95 (.ZN (n_99_95), .A (n_96_98), .B (n_91_98), .C1 (n_90_99), .C2 (n_88_100) );
AOI211_X1 g_100_93 (.ZN (n_100_93), .A (n_98_97), .B (n_93_97), .C1 (n_92_100), .C2 (n_87_98) );
AOI211_X1 g_98_94 (.ZN (n_98_94), .A (n_99_95), .B (n_94_99), .C1 (n_91_98), .C2 (n_89_97) );
AOI211_X1 g_97_96 (.ZN (n_97_96), .A (n_100_93), .B (n_96_98), .C1 (n_93_97), .C2 (n_90_99) );
AOI211_X1 g_95_97 (.ZN (n_95_97), .A (n_98_94), .B (n_98_97), .C1 (n_94_99), .C2 (n_92_100) );
AOI211_X1 g_93_98 (.ZN (n_93_98), .A (n_97_96), .B (n_99_95), .C1 (n_96_98), .C2 (n_91_98) );
AOI211_X1 g_91_99 (.ZN (n_91_99), .A (n_95_97), .B (n_100_93), .C1 (n_98_97), .C2 (n_93_97) );
AOI211_X1 g_89_100 (.ZN (n_89_100), .A (n_93_98), .B (n_98_94), .C1 (n_99_95), .C2 (n_94_99) );
AOI211_X1 g_90_98 (.ZN (n_90_98), .A (n_91_99), .B (n_97_96), .C1 (n_100_93), .C2 (n_96_98) );
AOI211_X1 g_92_97 (.ZN (n_92_97), .A (n_89_100), .B (n_95_97), .C1 (n_98_94), .C2 (n_98_97) );
AOI211_X1 g_94_96 (.ZN (n_94_96), .A (n_90_98), .B (n_93_98), .C1 (n_97_96), .C2 (n_99_95) );
AOI211_X1 g_95_98 (.ZN (n_95_98), .A (n_92_97), .B (n_91_99), .C1 (n_95_97), .C2 (n_100_93) );
AOI211_X1 g_97_97 (.ZN (n_97_97), .A (n_94_96), .B (n_89_100), .C1 (n_93_98), .C2 (n_98_94) );
AOI211_X1 g_96_95 (.ZN (n_96_95), .A (n_95_98), .B (n_90_98), .C1 (n_91_99), .C2 (n_97_96) );
AOI211_X1 g_97_93 (.ZN (n_97_93), .A (n_97_97), .B (n_92_97), .C1 (n_89_100), .C2 (n_95_97) );
AOI211_X1 g_98_95 (.ZN (n_98_95), .A (n_96_95), .B (n_94_96), .C1 (n_90_98), .C2 (n_93_98) );
AOI211_X1 g_99_93 (.ZN (n_99_93), .A (n_97_93), .B (n_95_98), .C1 (n_92_97), .C2 (n_91_99) );
AOI211_X1 g_100_91 (.ZN (n_100_91), .A (n_98_95), .B (n_97_97), .C1 (n_94_96), .C2 (n_89_100) );
AOI211_X1 g_98_92 (.ZN (n_98_92), .A (n_99_93), .B (n_96_95), .C1 (n_95_98), .C2 (n_90_98) );
AOI211_X1 g_97_94 (.ZN (n_97_94), .A (n_100_91), .B (n_97_93), .C1 (n_97_97), .C2 (n_92_97) );
AOI211_X1 g_96_96 (.ZN (n_96_96), .A (n_98_92), .B (n_98_95), .C1 (n_96_95), .C2 (n_94_96) );
AOI211_X1 g_94_97 (.ZN (n_94_97), .A (n_97_94), .B (n_99_93), .C1 (n_97_93), .C2 (n_95_98) );
AOI211_X1 g_92_98 (.ZN (n_92_98), .A (n_96_96), .B (n_100_91), .C1 (n_98_95), .C2 (n_97_97) );
AOI211_X1 g_91_96 (.ZN (n_91_96), .A (n_94_97), .B (n_98_92), .C1 (n_99_93), .C2 (n_96_95) );
AOI211_X1 g_93_95 (.ZN (n_93_95), .A (n_92_98), .B (n_97_94), .C1 (n_100_91), .C2 (n_97_93) );
AOI211_X1 g_95_96 (.ZN (n_95_96), .A (n_91_96), .B (n_96_96), .C1 (n_98_92), .C2 (n_98_95) );
AOI211_X1 g_97_95 (.ZN (n_97_95), .A (n_93_95), .B (n_94_97), .C1 (n_97_94), .C2 (n_99_93) );
AOI211_X1 g_95_94 (.ZN (n_95_94), .A (n_95_96), .B (n_92_98), .C1 (n_96_96), .C2 (n_100_91) );
AOI211_X1 g_96_92 (.ZN (n_96_92), .A (n_97_95), .B (n_91_96), .C1 (n_94_97), .C2 (n_98_92) );
AOI211_X1 g_98_91 (.ZN (n_98_91), .A (n_95_94), .B (n_93_95), .C1 (n_92_98), .C2 (n_97_94) );
AOI211_X1 g_99_89 (.ZN (n_99_89), .A (n_96_92), .B (n_95_96), .C1 (n_91_96), .C2 (n_96_96) );
AOI211_X1 g_100_87 (.ZN (n_100_87), .A (n_98_91), .B (n_97_95), .C1 (n_93_95), .C2 (n_94_97) );
AOI211_X1 g_99_85 (.ZN (n_99_85), .A (n_99_89), .B (n_95_94), .C1 (n_95_96), .C2 (n_92_98) );
AOI211_X1 g_100_83 (.ZN (n_100_83), .A (n_100_87), .B (n_96_92), .C1 (n_97_95), .C2 (n_91_96) );
AOI211_X1 g_99_81 (.ZN (n_99_81), .A (n_99_85), .B (n_98_91), .C1 (n_95_94), .C2 (n_93_95) );
AOI211_X1 g_98_79 (.ZN (n_98_79), .A (n_100_83), .B (n_99_89), .C1 (n_96_92), .C2 (n_95_96) );
AOI211_X1 g_96_78 (.ZN (n_96_78), .A (n_99_81), .B (n_100_87), .C1 (n_98_91), .C2 (n_97_95) );
AOI211_X1 g_98_77 (.ZN (n_98_77), .A (n_98_79), .B (n_99_85), .C1 (n_99_89), .C2 (n_95_94) );
AOI211_X1 g_96_76 (.ZN (n_96_76), .A (n_96_78), .B (n_100_83), .C1 (n_100_87), .C2 (n_96_92) );
AOI211_X1 g_94_77 (.ZN (n_94_77), .A (n_98_77), .B (n_99_81), .C1 (n_99_85), .C2 (n_98_91) );
AOI211_X1 g_92_78 (.ZN (n_92_78), .A (n_96_76), .B (n_98_79), .C1 (n_100_83), .C2 (n_99_89) );
AOI211_X1 g_93_76 (.ZN (n_93_76), .A (n_94_77), .B (n_96_78), .C1 (n_99_81), .C2 (n_100_87) );
AOI211_X1 g_91_77 (.ZN (n_91_77), .A (n_92_78), .B (n_98_77), .C1 (n_98_79), .C2 (n_99_85) );
AOI211_X1 g_89_78 (.ZN (n_89_78), .A (n_93_76), .B (n_96_76), .C1 (n_96_78), .C2 (n_100_83) );
AOI211_X1 g_87_79 (.ZN (n_87_79), .A (n_91_77), .B (n_94_77), .C1 (n_98_77), .C2 (n_99_81) );
AOI211_X1 g_85_80 (.ZN (n_85_80), .A (n_89_78), .B (n_92_78), .C1 (n_96_76), .C2 (n_98_79) );
AOI211_X1 g_83_81 (.ZN (n_83_81), .A (n_87_79), .B (n_93_76), .C1 (n_94_77), .C2 (n_96_78) );
AOI211_X1 g_82_83 (.ZN (n_82_83), .A (n_85_80), .B (n_91_77), .C1 (n_92_78), .C2 (n_98_77) );
AOI211_X1 g_84_82 (.ZN (n_84_82), .A (n_83_81), .B (n_89_78), .C1 (n_93_76), .C2 (n_96_76) );
AOI211_X1 g_86_81 (.ZN (n_86_81), .A (n_82_83), .B (n_87_79), .C1 (n_91_77), .C2 (n_94_77) );
AOI211_X1 g_88_80 (.ZN (n_88_80), .A (n_84_82), .B (n_85_80), .C1 (n_89_78), .C2 (n_92_78) );
AOI211_X1 g_90_79 (.ZN (n_90_79), .A (n_86_81), .B (n_83_81), .C1 (n_87_79), .C2 (n_93_76) );
AOI211_X1 g_89_81 (.ZN (n_89_81), .A (n_88_80), .B (n_82_83), .C1 (n_85_80), .C2 (n_91_77) );
AOI211_X1 g_88_79 (.ZN (n_88_79), .A (n_90_79), .B (n_84_82), .C1 (n_83_81), .C2 (n_89_78) );
AOI211_X1 g_90_78 (.ZN (n_90_78), .A (n_89_81), .B (n_86_81), .C1 (n_82_83), .C2 (n_87_79) );
AOI211_X1 g_91_80 (.ZN (n_91_80), .A (n_88_79), .B (n_88_80), .C1 (n_84_82), .C2 (n_85_80) );
AOI211_X1 g_93_79 (.ZN (n_93_79), .A (n_90_78), .B (n_90_79), .C1 (n_86_81), .C2 (n_83_81) );
AOI211_X1 g_95_78 (.ZN (n_95_78), .A (n_91_80), .B (n_89_81), .C1 (n_88_80), .C2 (n_82_83) );
AOI211_X1 g_97_79 (.ZN (n_97_79), .A (n_93_79), .B (n_88_79), .C1 (n_90_79), .C2 (n_84_82) );
AOI211_X1 g_95_80 (.ZN (n_95_80), .A (n_95_78), .B (n_90_78), .C1 (n_89_81), .C2 (n_86_81) );
AOI211_X1 g_94_78 (.ZN (n_94_78), .A (n_97_79), .B (n_91_80), .C1 (n_88_79), .C2 (n_88_80) );
AOI211_X1 g_92_79 (.ZN (n_92_79), .A (n_95_80), .B (n_93_79), .C1 (n_90_78), .C2 (n_90_79) );
AOI211_X1 g_90_80 (.ZN (n_90_80), .A (n_94_78), .B (n_95_78), .C1 (n_91_80), .C2 (n_89_81) );
AOI211_X1 g_88_81 (.ZN (n_88_81), .A (n_92_79), .B (n_97_79), .C1 (n_93_79), .C2 (n_88_79) );
AOI211_X1 g_86_80 (.ZN (n_86_80), .A (n_90_80), .B (n_95_80), .C1 (n_95_78), .C2 (n_90_78) );
AOI211_X1 g_84_81 (.ZN (n_84_81), .A (n_88_81), .B (n_94_78), .C1 (n_97_79), .C2 (n_91_80) );
AOI211_X1 g_82_82 (.ZN (n_82_82), .A (n_86_80), .B (n_92_79), .C1 (n_95_80), .C2 (n_93_79) );
AOI211_X1 g_80_83 (.ZN (n_80_83), .A (n_84_81), .B (n_90_80), .C1 (n_94_78), .C2 (n_95_78) );
AOI211_X1 g_78_84 (.ZN (n_78_84), .A (n_82_82), .B (n_88_81), .C1 (n_92_79), .C2 (n_97_79) );
AOI211_X1 g_76_85 (.ZN (n_76_85), .A (n_80_83), .B (n_86_80), .C1 (n_90_80), .C2 (n_95_80) );
AOI211_X1 g_74_86 (.ZN (n_74_86), .A (n_78_84), .B (n_84_81), .C1 (n_88_81), .C2 (n_94_78) );
AOI211_X1 g_72_87 (.ZN (n_72_87), .A (n_76_85), .B (n_82_82), .C1 (n_86_80), .C2 (n_92_79) );
AOI211_X1 g_71_89 (.ZN (n_71_89), .A (n_74_86), .B (n_80_83), .C1 (n_84_81), .C2 (n_90_80) );
AOI211_X1 g_69_88 (.ZN (n_69_88), .A (n_72_87), .B (n_78_84), .C1 (n_82_82), .C2 (n_88_81) );
AOI211_X1 g_71_87 (.ZN (n_71_87), .A (n_71_89), .B (n_76_85), .C1 (n_80_83), .C2 (n_86_80) );
AOI211_X1 g_73_86 (.ZN (n_73_86), .A (n_69_88), .B (n_74_86), .C1 (n_78_84), .C2 (n_84_81) );
AOI211_X1 g_75_85 (.ZN (n_75_85), .A (n_71_87), .B (n_72_87), .C1 (n_76_85), .C2 (n_82_82) );
AOI211_X1 g_77_84 (.ZN (n_77_84), .A (n_73_86), .B (n_71_89), .C1 (n_74_86), .C2 (n_80_83) );
AOI211_X1 g_79_83 (.ZN (n_79_83), .A (n_75_85), .B (n_69_88), .C1 (n_72_87), .C2 (n_78_84) );
AOI211_X1 g_78_85 (.ZN (n_78_85), .A (n_77_84), .B (n_71_87), .C1 (n_71_89), .C2 (n_76_85) );
AOI211_X1 g_80_84 (.ZN (n_80_84), .A (n_79_83), .B (n_73_86), .C1 (n_69_88), .C2 (n_74_86) );
AOI211_X1 g_79_86 (.ZN (n_79_86), .A (n_78_85), .B (n_75_85), .C1 (n_71_87), .C2 (n_72_87) );
AOI211_X1 g_77_85 (.ZN (n_77_85), .A (n_80_84), .B (n_77_84), .C1 (n_73_86), .C2 (n_71_89) );
AOI211_X1 g_79_84 (.ZN (n_79_84), .A (n_79_86), .B (n_79_83), .C1 (n_75_85), .C2 (n_69_88) );
AOI211_X1 g_81_85 (.ZN (n_81_85), .A (n_77_85), .B (n_78_85), .C1 (n_77_84), .C2 (n_71_87) );
AOI211_X1 g_83_84 (.ZN (n_83_84), .A (n_79_84), .B (n_80_84), .C1 (n_79_83), .C2 (n_73_86) );
AOI211_X1 g_85_83 (.ZN (n_85_83), .A (n_81_85), .B (n_79_86), .C1 (n_78_85), .C2 (n_75_85) );
AOI211_X1 g_87_82 (.ZN (n_87_82), .A (n_83_84), .B (n_77_85), .C1 (n_80_84), .C2 (n_77_84) );
AOI211_X1 g_89_83 (.ZN (n_89_83), .A (n_85_83), .B (n_79_84), .C1 (n_79_86), .C2 (n_79_83) );
AOI211_X1 g_91_82 (.ZN (n_91_82), .A (n_87_82), .B (n_81_85), .C1 (n_77_85), .C2 (n_78_85) );
AOI211_X1 g_93_81 (.ZN (n_93_81), .A (n_89_83), .B (n_83_84), .C1 (n_79_84), .C2 (n_80_84) );
AOI211_X1 g_94_79 (.ZN (n_94_79), .A (n_91_82), .B (n_85_83), .C1 (n_81_85), .C2 (n_79_86) );
AOI211_X1 g_95_77 (.ZN (n_95_77), .A (n_93_81), .B (n_87_82), .C1 (n_83_84), .C2 (n_77_85) );
AOI211_X1 g_93_78 (.ZN (n_93_78), .A (n_94_79), .B (n_89_83), .C1 (n_85_83), .C2 (n_79_84) );
AOI211_X1 g_92_80 (.ZN (n_92_80), .A (n_95_77), .B (n_91_82), .C1 (n_87_82), .C2 (n_81_85) );
AOI211_X1 g_90_81 (.ZN (n_90_81), .A (n_93_78), .B (n_93_81), .C1 (n_89_83), .C2 (n_83_84) );
AOI211_X1 g_91_79 (.ZN (n_91_79), .A (n_92_80), .B (n_94_79), .C1 (n_91_82), .C2 (n_85_83) );
AOI211_X1 g_89_80 (.ZN (n_89_80), .A (n_90_81), .B (n_95_77), .C1 (n_93_81), .C2 (n_87_82) );
AOI211_X1 g_87_81 (.ZN (n_87_81), .A (n_91_79), .B (n_93_78), .C1 (n_94_79), .C2 (n_89_83) );
AOI211_X1 g_85_82 (.ZN (n_85_82), .A (n_89_80), .B (n_92_80), .C1 (n_95_77), .C2 (n_91_82) );
AOI211_X1 g_83_83 (.ZN (n_83_83), .A (n_87_81), .B (n_90_81), .C1 (n_93_78), .C2 (n_93_81) );
AOI211_X1 g_81_84 (.ZN (n_81_84), .A (n_85_82), .B (n_91_79), .C1 (n_92_80), .C2 (n_94_79) );
AOI211_X1 g_79_85 (.ZN (n_79_85), .A (n_83_83), .B (n_89_80), .C1 (n_90_81), .C2 (n_95_77) );
AOI211_X1 g_77_86 (.ZN (n_77_86), .A (n_81_84), .B (n_87_81), .C1 (n_91_79), .C2 (n_93_78) );
AOI211_X1 g_75_87 (.ZN (n_75_87), .A (n_79_85), .B (n_85_82), .C1 (n_89_80), .C2 (n_92_80) );
AOI211_X1 g_73_88 (.ZN (n_73_88), .A (n_77_86), .B (n_83_83), .C1 (n_87_81), .C2 (n_90_81) );
AOI211_X1 g_72_90 (.ZN (n_72_90), .A (n_75_87), .B (n_81_84), .C1 (n_85_82), .C2 (n_91_79) );
AOI211_X1 g_71_88 (.ZN (n_71_88), .A (n_73_88), .B (n_79_85), .C1 (n_83_83), .C2 (n_89_80) );
AOI211_X1 g_73_87 (.ZN (n_73_87), .A (n_72_90), .B (n_77_86), .C1 (n_81_84), .C2 (n_87_81) );
AOI211_X1 g_75_86 (.ZN (n_75_86), .A (n_71_88), .B (n_75_87), .C1 (n_79_85), .C2 (n_85_82) );
AOI211_X1 g_77_87 (.ZN (n_77_87), .A (n_73_87), .B (n_73_88), .C1 (n_77_86), .C2 (n_83_83) );
AOI211_X1 g_75_88 (.ZN (n_75_88), .A (n_75_86), .B (n_72_90), .C1 (n_75_87), .C2 (n_81_84) );
AOI211_X1 g_76_86 (.ZN (n_76_86), .A (n_77_87), .B (n_71_88), .C1 (n_73_88), .C2 (n_79_85) );
AOI211_X1 g_74_87 (.ZN (n_74_87), .A (n_75_88), .B (n_73_87), .C1 (n_72_90), .C2 (n_77_86) );
AOI211_X1 g_72_88 (.ZN (n_72_88), .A (n_76_86), .B (n_75_86), .C1 (n_71_88), .C2 (n_75_87) );
AOI211_X1 g_70_89 (.ZN (n_70_89), .A (n_74_87), .B (n_77_87), .C1 (n_73_87), .C2 (n_73_88) );
AOI211_X1 g_68_90 (.ZN (n_68_90), .A (n_72_88), .B (n_75_88), .C1 (n_75_86), .C2 (n_72_90) );
AOI211_X1 g_66_91 (.ZN (n_66_91), .A (n_70_89), .B (n_76_86), .C1 (n_77_87), .C2 (n_71_88) );
AOI211_X1 g_67_89 (.ZN (n_67_89), .A (n_68_90), .B (n_74_87), .C1 (n_75_88), .C2 (n_73_87) );
AOI211_X1 g_65_90 (.ZN (n_65_90), .A (n_66_91), .B (n_72_88), .C1 (n_76_86), .C2 (n_75_86) );
AOI211_X1 g_64_92 (.ZN (n_64_92), .A (n_67_89), .B (n_70_89), .C1 (n_74_87), .C2 (n_77_87) );
AOI211_X1 g_62_93 (.ZN (n_62_93), .A (n_65_90), .B (n_68_90), .C1 (n_72_88), .C2 (n_75_88) );
AOI211_X1 g_63_91 (.ZN (n_63_91), .A (n_64_92), .B (n_66_91), .C1 (n_70_89), .C2 (n_76_86) );
AOI211_X1 g_64_89 (.ZN (n_64_89), .A (n_62_93), .B (n_67_89), .C1 (n_68_90), .C2 (n_74_87) );
AOI211_X1 g_62_90 (.ZN (n_62_90), .A (n_63_91), .B (n_65_90), .C1 (n_66_91), .C2 (n_72_88) );
AOI211_X1 g_60_91 (.ZN (n_60_91), .A (n_64_89), .B (n_64_92), .C1 (n_67_89), .C2 (n_70_89) );
AOI211_X1 g_58_92 (.ZN (n_58_92), .A (n_62_90), .B (n_62_93), .C1 (n_65_90), .C2 (n_68_90) );
AOI211_X1 g_56_93 (.ZN (n_56_93), .A (n_60_91), .B (n_63_91), .C1 (n_64_92), .C2 (n_66_91) );
AOI211_X1 g_55_95 (.ZN (n_55_95), .A (n_58_92), .B (n_64_89), .C1 (n_62_93), .C2 (n_67_89) );
AOI211_X1 g_54_97 (.ZN (n_54_97), .A (n_56_93), .B (n_62_90), .C1 (n_63_91), .C2 (n_65_90) );
AOI211_X1 g_55_99 (.ZN (n_55_99), .A (n_55_95), .B (n_60_91), .C1 (n_64_89), .C2 (n_64_92) );
AOI211_X1 g_56_97 (.ZN (n_56_97), .A (n_54_97), .B (n_58_92), .C1 (n_62_90), .C2 (n_62_93) );
AOI211_X1 g_57_95 (.ZN (n_57_95), .A (n_55_99), .B (n_56_93), .C1 (n_60_91), .C2 (n_63_91) );
AOI211_X1 g_59_94 (.ZN (n_59_94), .A (n_56_97), .B (n_55_95), .C1 (n_58_92), .C2 (n_64_89) );
AOI211_X1 g_61_93 (.ZN (n_61_93), .A (n_57_95), .B (n_54_97), .C1 (n_56_93), .C2 (n_62_90) );
AOI211_X1 g_63_92 (.ZN (n_63_92), .A (n_59_94), .B (n_55_99), .C1 (n_55_95), .C2 (n_60_91) );
AOI211_X1 g_65_91 (.ZN (n_65_91), .A (n_61_93), .B (n_56_97), .C1 (n_54_97), .C2 (n_58_92) );
AOI211_X1 g_67_90 (.ZN (n_67_90), .A (n_63_92), .B (n_57_95), .C1 (n_55_99), .C2 (n_56_93) );
AOI211_X1 g_69_89 (.ZN (n_69_89), .A (n_65_91), .B (n_59_94), .C1 (n_56_97), .C2 (n_55_95) );
AOI211_X1 g_70_91 (.ZN (n_70_91), .A (n_67_90), .B (n_61_93), .C1 (n_57_95), .C2 (n_54_97) );
AOI211_X1 g_68_92 (.ZN (n_68_92), .A (n_69_89), .B (n_63_92), .C1 (n_59_94), .C2 (n_55_99) );
AOI211_X1 g_69_90 (.ZN (n_69_90), .A (n_70_91), .B (n_65_91), .C1 (n_61_93), .C2 (n_56_97) );
AOI211_X1 g_67_91 (.ZN (n_67_91), .A (n_68_92), .B (n_67_90), .C1 (n_63_92), .C2 (n_57_95) );
AOI211_X1 g_68_89 (.ZN (n_68_89), .A (n_69_90), .B (n_69_89), .C1 (n_65_91), .C2 (n_59_94) );
AOI211_X1 g_66_90 (.ZN (n_66_90), .A (n_67_91), .B (n_70_91), .C1 (n_67_90), .C2 (n_61_93) );
AOI211_X1 g_64_91 (.ZN (n_64_91), .A (n_68_89), .B (n_68_92), .C1 (n_69_89), .C2 (n_63_92) );
AOI211_X1 g_62_92 (.ZN (n_62_92), .A (n_66_90), .B (n_69_90), .C1 (n_70_91), .C2 (n_65_91) );
AOI211_X1 g_60_93 (.ZN (n_60_93), .A (n_64_91), .B (n_67_91), .C1 (n_68_92), .C2 (n_67_90) );
AOI211_X1 g_58_94 (.ZN (n_58_94), .A (n_62_92), .B (n_68_89), .C1 (n_69_90), .C2 (n_69_89) );
AOI211_X1 g_57_96 (.ZN (n_57_96), .A (n_60_93), .B (n_66_90), .C1 (n_67_91), .C2 (n_70_91) );
AOI211_X1 g_56_98 (.ZN (n_56_98), .A (n_58_94), .B (n_64_91), .C1 (n_68_89), .C2 (n_68_92) );
AOI211_X1 g_57_100 (.ZN (n_57_100), .A (n_57_96), .B (n_62_92), .C1 (n_66_90), .C2 (n_69_90) );
AOI211_X1 g_58_98 (.ZN (n_58_98), .A (n_56_98), .B (n_60_93), .C1 (n_64_91), .C2 (n_67_91) );
AOI211_X1 g_59_96 (.ZN (n_59_96), .A (n_57_100), .B (n_58_94), .C1 (n_62_92), .C2 (n_68_89) );
AOI211_X1 g_61_95 (.ZN (n_61_95), .A (n_58_98), .B (n_57_96), .C1 (n_60_93), .C2 (n_66_90) );
AOI211_X1 g_63_94 (.ZN (n_63_94), .A (n_59_96), .B (n_56_98), .C1 (n_58_94), .C2 (n_64_91) );
AOI211_X1 g_65_93 (.ZN (n_65_93), .A (n_61_95), .B (n_57_100), .C1 (n_57_96), .C2 (n_62_92) );
AOI211_X1 g_67_92 (.ZN (n_67_92), .A (n_63_94), .B (n_58_98), .C1 (n_56_98), .C2 (n_60_93) );
AOI211_X1 g_69_91 (.ZN (n_69_91), .A (n_65_93), .B (n_59_96), .C1 (n_57_100), .C2 (n_58_94) );
AOI211_X1 g_71_90 (.ZN (n_71_90), .A (n_67_92), .B (n_61_95), .C1 (n_58_98), .C2 (n_57_96) );
AOI211_X1 g_73_89 (.ZN (n_73_89), .A (n_69_91), .B (n_63_94), .C1 (n_59_96), .C2 (n_56_98) );
AOI211_X1 g_72_91 (.ZN (n_72_91), .A (n_71_90), .B (n_65_93), .C1 (n_61_95), .C2 (n_57_100) );
AOI211_X1 g_70_90 (.ZN (n_70_90), .A (n_73_89), .B (n_67_92), .C1 (n_63_94), .C2 (n_58_98) );
AOI211_X1 g_72_89 (.ZN (n_72_89), .A (n_72_91), .B (n_69_91), .C1 (n_65_93), .C2 (n_59_96) );
AOI211_X1 g_74_88 (.ZN (n_74_88), .A (n_70_90), .B (n_71_90), .C1 (n_67_92), .C2 (n_61_95) );
AOI211_X1 g_76_87 (.ZN (n_76_87), .A (n_72_89), .B (n_73_89), .C1 (n_69_91), .C2 (n_63_94) );
AOI211_X1 g_78_86 (.ZN (n_78_86), .A (n_74_88), .B (n_72_91), .C1 (n_71_90), .C2 (n_65_93) );
AOI211_X1 g_80_85 (.ZN (n_80_85), .A (n_76_87), .B (n_70_90), .C1 (n_73_89), .C2 (n_67_92) );
AOI211_X1 g_82_84 (.ZN (n_82_84), .A (n_78_86), .B (n_72_89), .C1 (n_72_91), .C2 (n_69_91) );
AOI211_X1 g_84_83 (.ZN (n_84_83), .A (n_80_85), .B (n_74_88), .C1 (n_70_90), .C2 (n_71_90) );
AOI211_X1 g_86_82 (.ZN (n_86_82), .A (n_82_84), .B (n_76_87), .C1 (n_72_89), .C2 (n_73_89) );
AOI211_X1 g_85_84 (.ZN (n_85_84), .A (n_84_83), .B (n_78_86), .C1 (n_74_88), .C2 (n_72_91) );
AOI211_X1 g_87_83 (.ZN (n_87_83), .A (n_86_82), .B (n_80_85), .C1 (n_76_87), .C2 (n_70_90) );
AOI211_X1 g_89_82 (.ZN (n_89_82), .A (n_85_84), .B (n_82_84), .C1 (n_78_86), .C2 (n_72_89) );
AOI211_X1 g_91_81 (.ZN (n_91_81), .A (n_87_83), .B (n_84_83), .C1 (n_80_85), .C2 (n_74_88) );
AOI211_X1 g_93_80 (.ZN (n_93_80), .A (n_89_82), .B (n_86_82), .C1 (n_82_84), .C2 (n_76_87) );
AOI211_X1 g_95_79 (.ZN (n_95_79), .A (n_91_81), .B (n_85_84), .C1 (n_84_83), .C2 (n_78_86) );
AOI211_X1 g_97_78 (.ZN (n_97_78), .A (n_93_80), .B (n_87_83), .C1 (n_86_82), .C2 (n_80_85) );
AOI211_X1 g_99_79 (.ZN (n_99_79), .A (n_95_79), .B (n_89_82), .C1 (n_85_84), .C2 (n_82_84) );
AOI211_X1 g_97_80 (.ZN (n_97_80), .A (n_97_78), .B (n_91_81), .C1 (n_87_83), .C2 (n_84_83) );
AOI211_X1 g_98_82 (.ZN (n_98_82), .A (n_99_79), .B (n_93_80), .C1 (n_89_82), .C2 (n_86_82) );
AOI211_X1 g_100_81 (.ZN (n_100_81), .A (n_97_80), .B (n_95_79), .C1 (n_91_81), .C2 (n_85_84) );
AOI211_X1 g_98_80 (.ZN (n_98_80), .A (n_98_82), .B (n_97_78), .C1 (n_93_80), .C2 (n_87_83) );
AOI211_X1 g_96_79 (.ZN (n_96_79), .A (n_100_81), .B (n_99_79), .C1 (n_95_79), .C2 (n_89_82) );
AOI211_X1 g_97_81 (.ZN (n_97_81), .A (n_98_80), .B (n_97_80), .C1 (n_97_78), .C2 (n_91_81) );
AOI211_X1 g_98_83 (.ZN (n_98_83), .A (n_96_79), .B (n_98_82), .C1 (n_99_79), .C2 (n_93_80) );
AOI211_X1 g_96_82 (.ZN (n_96_82), .A (n_97_81), .B (n_100_81), .C1 (n_97_80), .C2 (n_95_79) );
AOI211_X1 g_98_81 (.ZN (n_98_81), .A (n_98_83), .B (n_98_80), .C1 (n_98_82), .C2 (n_97_78) );
AOI211_X1 g_96_80 (.ZN (n_96_80), .A (n_96_82), .B (n_96_79), .C1 (n_100_81), .C2 (n_99_79) );
AOI211_X1 g_94_81 (.ZN (n_94_81), .A (n_98_81), .B (n_97_81), .C1 (n_98_80), .C2 (n_97_80) );
AOI211_X1 g_92_82 (.ZN (n_92_82), .A (n_96_80), .B (n_98_83), .C1 (n_96_79), .C2 (n_98_82) );
AOI211_X1 g_90_83 (.ZN (n_90_83), .A (n_94_81), .B (n_96_82), .C1 (n_97_81), .C2 (n_100_81) );
AOI211_X1 g_88_82 (.ZN (n_88_82), .A (n_92_82), .B (n_98_81), .C1 (n_98_83), .C2 (n_98_80) );
AOI211_X1 g_86_83 (.ZN (n_86_83), .A (n_90_83), .B (n_96_80), .C1 (n_96_82), .C2 (n_96_79) );
AOI211_X1 g_84_84 (.ZN (n_84_84), .A (n_88_82), .B (n_94_81), .C1 (n_98_81), .C2 (n_97_81) );
AOI211_X1 g_82_85 (.ZN (n_82_85), .A (n_86_83), .B (n_92_82), .C1 (n_96_80), .C2 (n_98_83) );
AOI211_X1 g_80_86 (.ZN (n_80_86), .A (n_84_84), .B (n_90_83), .C1 (n_94_81), .C2 (n_96_82) );
AOI211_X1 g_78_87 (.ZN (n_78_87), .A (n_82_85), .B (n_88_82), .C1 (n_92_82), .C2 (n_98_81) );
AOI211_X1 g_76_88 (.ZN (n_76_88), .A (n_80_86), .B (n_86_83), .C1 (n_90_83), .C2 (n_96_80) );
AOI211_X1 g_74_89 (.ZN (n_74_89), .A (n_78_87), .B (n_84_84), .C1 (n_88_82), .C2 (n_94_81) );
AOI211_X1 g_73_91 (.ZN (n_73_91), .A (n_76_88), .B (n_82_85), .C1 (n_86_83), .C2 (n_92_82) );
AOI211_X1 g_75_90 (.ZN (n_75_90), .A (n_74_89), .B (n_80_86), .C1 (n_84_84), .C2 (n_90_83) );
AOI211_X1 g_77_89 (.ZN (n_77_89), .A (n_73_91), .B (n_78_87), .C1 (n_82_85), .C2 (n_88_82) );
AOI211_X1 g_79_88 (.ZN (n_79_88), .A (n_75_90), .B (n_76_88), .C1 (n_80_86), .C2 (n_86_83) );
AOI211_X1 g_81_87 (.ZN (n_81_87), .A (n_77_89), .B (n_74_89), .C1 (n_78_87), .C2 (n_84_84) );
AOI211_X1 g_83_86 (.ZN (n_83_86), .A (n_79_88), .B (n_73_91), .C1 (n_76_88), .C2 (n_82_85) );
AOI211_X1 g_85_85 (.ZN (n_85_85), .A (n_81_87), .B (n_75_90), .C1 (n_74_89), .C2 (n_80_86) );
AOI211_X1 g_87_84 (.ZN (n_87_84), .A (n_83_86), .B (n_77_89), .C1 (n_73_91), .C2 (n_78_87) );
AOI211_X1 g_86_86 (.ZN (n_86_86), .A (n_85_85), .B (n_79_88), .C1 (n_75_90), .C2 (n_76_88) );
AOI211_X1 g_84_85 (.ZN (n_84_85), .A (n_87_84), .B (n_81_87), .C1 (n_77_89), .C2 (n_74_89) );
AOI211_X1 g_86_84 (.ZN (n_86_84), .A (n_86_86), .B (n_83_86), .C1 (n_79_88), .C2 (n_73_91) );
AOI211_X1 g_88_83 (.ZN (n_88_83), .A (n_84_85), .B (n_85_85), .C1 (n_81_87), .C2 (n_75_90) );
AOI211_X1 g_90_82 (.ZN (n_90_82), .A (n_86_84), .B (n_87_84), .C1 (n_83_86), .C2 (n_77_89) );
AOI211_X1 g_92_81 (.ZN (n_92_81), .A (n_88_83), .B (n_86_86), .C1 (n_85_85), .C2 (n_79_88) );
AOI211_X1 g_94_80 (.ZN (n_94_80), .A (n_90_82), .B (n_84_85), .C1 (n_87_84), .C2 (n_81_87) );
AOI211_X1 g_96_81 (.ZN (n_96_81), .A (n_92_81), .B (n_86_84), .C1 (n_86_86), .C2 (n_83_86) );
AOI211_X1 g_94_82 (.ZN (n_94_82), .A (n_94_80), .B (n_88_83), .C1 (n_84_85), .C2 (n_85_85) );
AOI211_X1 g_92_83 (.ZN (n_92_83), .A (n_96_81), .B (n_90_82), .C1 (n_86_84), .C2 (n_87_84) );
AOI211_X1 g_90_84 (.ZN (n_90_84), .A (n_94_82), .B (n_92_81), .C1 (n_88_83), .C2 (n_86_86) );
AOI211_X1 g_88_85 (.ZN (n_88_85), .A (n_92_83), .B (n_94_80), .C1 (n_90_82), .C2 (n_84_85) );
AOI211_X1 g_87_87 (.ZN (n_87_87), .A (n_90_84), .B (n_96_81), .C1 (n_92_81), .C2 (n_86_84) );
AOI211_X1 g_86_85 (.ZN (n_86_85), .A (n_88_85), .B (n_94_82), .C1 (n_94_80), .C2 (n_88_83) );
AOI211_X1 g_88_84 (.ZN (n_88_84), .A (n_87_87), .B (n_92_83), .C1 (n_96_81), .C2 (n_90_82) );
AOI211_X1 g_87_86 (.ZN (n_87_86), .A (n_86_85), .B (n_90_84), .C1 (n_94_82), .C2 (n_92_81) );
AOI211_X1 g_89_85 (.ZN (n_89_85), .A (n_88_84), .B (n_88_85), .C1 (n_92_83), .C2 (n_94_80) );
AOI211_X1 g_91_84 (.ZN (n_91_84), .A (n_87_86), .B (n_87_87), .C1 (n_90_84), .C2 (n_96_81) );
AOI211_X1 g_93_83 (.ZN (n_93_83), .A (n_89_85), .B (n_86_85), .C1 (n_88_85), .C2 (n_94_82) );
AOI211_X1 g_95_82 (.ZN (n_95_82), .A (n_91_84), .B (n_88_84), .C1 (n_87_87), .C2 (n_92_83) );
AOI211_X1 g_97_83 (.ZN (n_97_83), .A (n_93_83), .B (n_87_86), .C1 (n_86_85), .C2 (n_90_84) );
AOI211_X1 g_95_84 (.ZN (n_95_84), .A (n_95_82), .B (n_89_85), .C1 (n_88_84), .C2 (n_88_85) );
AOI211_X1 g_97_85 (.ZN (n_97_85), .A (n_97_83), .B (n_91_84), .C1 (n_87_86), .C2 (n_87_87) );
AOI211_X1 g_98_87 (.ZN (n_98_87), .A (n_95_84), .B (n_93_83), .C1 (n_89_85), .C2 (n_86_85) );
AOI211_X1 g_97_89 (.ZN (n_97_89), .A (n_97_85), .B (n_95_82), .C1 (n_91_84), .C2 (n_88_84) );
AOI211_X1 g_96_91 (.ZN (n_96_91), .A (n_98_87), .B (n_97_83), .C1 (n_93_83), .C2 (n_87_86) );
AOI211_X1 g_98_90 (.ZN (n_98_90), .A (n_97_89), .B (n_95_84), .C1 (n_95_82), .C2 (n_89_85) );
AOI211_X1 g_100_89 (.ZN (n_100_89), .A (n_96_91), .B (n_97_85), .C1 (n_97_83), .C2 (n_91_84) );
AOI211_X1 g_98_88 (.ZN (n_98_88), .A (n_98_90), .B (n_98_87), .C1 (n_95_84), .C2 (n_93_83) );
AOI211_X1 g_97_90 (.ZN (n_97_90), .A (n_100_89), .B (n_97_89), .C1 (n_97_85), .C2 (n_95_82) );
AOI211_X1 g_99_91 (.ZN (n_99_91), .A (n_98_88), .B (n_96_91), .C1 (n_98_87), .C2 (n_97_83) );
AOI211_X1 g_98_93 (.ZN (n_98_93), .A (n_97_90), .B (n_98_90), .C1 (n_97_89), .C2 (n_95_84) );
AOI211_X1 g_96_94 (.ZN (n_96_94), .A (n_99_91), .B (n_100_89), .C1 (n_96_91), .C2 (n_97_85) );
AOI211_X1 g_97_92 (.ZN (n_97_92), .A (n_98_93), .B (n_98_88), .C1 (n_98_90), .C2 (n_98_87) );
AOI211_X1 g_95_93 (.ZN (n_95_93), .A (n_96_94), .B (n_97_90), .C1 (n_100_89), .C2 (n_97_89) );
AOI211_X1 g_94_95 (.ZN (n_94_95), .A (n_97_92), .B (n_99_91), .C1 (n_98_88), .C2 (n_96_91) );
AOI211_X1 g_92_96 (.ZN (n_92_96), .A (n_95_93), .B (n_98_93), .C1 (n_97_90), .C2 (n_98_90) );
AOI211_X1 g_90_97 (.ZN (n_90_97), .A (n_94_95), .B (n_96_94), .C1 (n_99_91), .C2 (n_100_89) );
AOI211_X1 g_88_98 (.ZN (n_88_98), .A (n_92_96), .B (n_97_92), .C1 (n_98_93), .C2 (n_98_88) );
AOI211_X1 g_87_96 (.ZN (n_87_96), .A (n_90_97), .B (n_95_93), .C1 (n_96_94), .C2 (n_97_90) );
AOI211_X1 g_86_98 (.ZN (n_86_98), .A (n_88_98), .B (n_94_95), .C1 (n_97_92), .C2 (n_99_91) );
AOI211_X1 g_85_100 (.ZN (n_85_100), .A (n_87_96), .B (n_92_96), .C1 (n_95_93), .C2 (n_98_93) );
AOI211_X1 g_87_99 (.ZN (n_87_99), .A (n_86_98), .B (n_90_97), .C1 (n_94_95), .C2 (n_96_94) );
AOI211_X1 g_89_98 (.ZN (n_89_98), .A (n_85_100), .B (n_88_98), .C1 (n_92_96), .C2 (n_97_92) );
AOI211_X1 g_91_97 (.ZN (n_91_97), .A (n_87_99), .B (n_87_96), .C1 (n_90_97), .C2 (n_95_93) );
AOI211_X1 g_93_96 (.ZN (n_93_96), .A (n_89_98), .B (n_86_98), .C1 (n_88_98), .C2 (n_94_95) );
AOI211_X1 g_95_95 (.ZN (n_95_95), .A (n_91_97), .B (n_85_100), .C1 (n_87_96), .C2 (n_92_96) );
AOI211_X1 g_96_93 (.ZN (n_96_93), .A (n_93_96), .B (n_87_99), .C1 (n_86_98), .C2 (n_90_97) );
AOI211_X1 g_97_91 (.ZN (n_97_91), .A (n_95_95), .B (n_89_98), .C1 (n_85_100), .C2 (n_88_98) );
AOI211_X1 g_98_89 (.ZN (n_98_89), .A (n_96_93), .B (n_91_97), .C1 (n_87_99), .C2 (n_87_96) );
AOI211_X1 g_99_87 (.ZN (n_99_87), .A (n_97_91), .B (n_93_96), .C1 (n_89_98), .C2 (n_86_98) );
AOI211_X1 g_100_85 (.ZN (n_100_85), .A (n_98_89), .B (n_95_95), .C1 (n_91_97), .C2 (n_85_100) );
AOI211_X1 g_99_83 (.ZN (n_99_83), .A (n_99_87), .B (n_96_93), .C1 (n_93_96), .C2 (n_87_99) );
AOI211_X1 g_98_85 (.ZN (n_98_85), .A (n_100_85), .B (n_97_91), .C1 (n_95_95), .C2 (n_89_98) );
AOI211_X1 g_97_87 (.ZN (n_97_87), .A (n_99_83), .B (n_98_89), .C1 (n_96_93), .C2 (n_91_97) );
AOI211_X1 g_96_89 (.ZN (n_96_89), .A (n_98_85), .B (n_99_87), .C1 (n_97_91), .C2 (n_93_96) );
AOI211_X1 g_95_91 (.ZN (n_95_91), .A (n_97_87), .B (n_100_85), .C1 (n_98_89), .C2 (n_95_95) );
AOI211_X1 g_94_93 (.ZN (n_94_93), .A (n_96_89), .B (n_99_83), .C1 (n_99_87), .C2 (n_96_93) );
AOI211_X1 g_92_94 (.ZN (n_92_94), .A (n_95_91), .B (n_98_85), .C1 (n_100_85), .C2 (n_97_91) );
AOI211_X1 g_90_95 (.ZN (n_90_95), .A (n_94_93), .B (n_97_87), .C1 (n_99_83), .C2 (n_98_89) );
AOI211_X1 g_88_96 (.ZN (n_88_96), .A (n_92_94), .B (n_96_89), .C1 (n_98_85), .C2 (n_99_87) );
AOI211_X1 g_86_97 (.ZN (n_86_97), .A (n_90_95), .B (n_95_91), .C1 (n_97_87), .C2 (n_100_85) );
AOI211_X1 g_84_98 (.ZN (n_84_98), .A (n_88_96), .B (n_94_93), .C1 (n_96_89), .C2 (n_99_83) );
AOI211_X1 g_83_96 (.ZN (n_83_96), .A (n_86_97), .B (n_92_94), .C1 (n_95_91), .C2 (n_98_85) );
AOI211_X1 g_82_98 (.ZN (n_82_98), .A (n_84_98), .B (n_90_95), .C1 (n_94_93), .C2 (n_97_87) );
AOI211_X1 g_81_100 (.ZN (n_81_100), .A (n_83_96), .B (n_88_96), .C1 (n_92_94), .C2 (n_96_89) );
AOI211_X1 g_83_99 (.ZN (n_83_99), .A (n_82_98), .B (n_86_97), .C1 (n_90_95), .C2 (n_95_91) );
AOI211_X1 g_85_98 (.ZN (n_85_98), .A (n_81_100), .B (n_84_98), .C1 (n_88_96), .C2 (n_94_93) );
AOI211_X1 g_87_97 (.ZN (n_87_97), .A (n_83_99), .B (n_83_96), .C1 (n_86_97), .C2 (n_92_94) );
AOI211_X1 g_89_96 (.ZN (n_89_96), .A (n_85_98), .B (n_82_98), .C1 (n_84_98), .C2 (n_90_95) );
AOI211_X1 g_91_95 (.ZN (n_91_95), .A (n_87_97), .B (n_81_100), .C1 (n_83_96), .C2 (n_88_96) );
AOI211_X1 g_93_94 (.ZN (n_93_94), .A (n_89_96), .B (n_83_99), .C1 (n_82_98), .C2 (n_86_97) );
AOI211_X1 g_94_92 (.ZN (n_94_92), .A (n_91_95), .B (n_85_98), .C1 (n_81_100), .C2 (n_84_98) );
AOI211_X1 g_95_90 (.ZN (n_95_90), .A (n_93_94), .B (n_87_97), .C1 (n_83_99), .C2 (n_83_96) );
AOI211_X1 g_96_88 (.ZN (n_96_88), .A (n_94_92), .B (n_89_96), .C1 (n_85_98), .C2 (n_82_98) );
AOI211_X1 g_97_86 (.ZN (n_97_86), .A (n_95_90), .B (n_91_95), .C1 (n_87_97), .C2 (n_81_100) );
AOI211_X1 g_98_84 (.ZN (n_98_84), .A (n_96_88), .B (n_93_94), .C1 (n_89_96), .C2 (n_83_99) );
AOI211_X1 g_97_82 (.ZN (n_97_82), .A (n_97_86), .B (n_94_92), .C1 (n_91_95), .C2 (n_85_98) );
AOI211_X1 g_95_81 (.ZN (n_95_81), .A (n_98_84), .B (n_95_90), .C1 (n_93_94), .C2 (n_87_97) );
AOI211_X1 g_96_83 (.ZN (n_96_83), .A (n_97_82), .B (n_96_88), .C1 (n_94_92), .C2 (n_89_96) );
AOI211_X1 g_94_84 (.ZN (n_94_84), .A (n_95_81), .B (n_97_86), .C1 (n_95_90), .C2 (n_91_95) );
AOI211_X1 g_93_82 (.ZN (n_93_82), .A (n_96_83), .B (n_98_84), .C1 (n_96_88), .C2 (n_93_94) );
AOI211_X1 g_91_83 (.ZN (n_91_83), .A (n_94_84), .B (n_97_82), .C1 (n_97_86), .C2 (n_94_92) );
AOI211_X1 g_89_84 (.ZN (n_89_84), .A (n_93_82), .B (n_95_81), .C1 (n_98_84), .C2 (n_95_90) );
AOI211_X1 g_87_85 (.ZN (n_87_85), .A (n_91_83), .B (n_96_83), .C1 (n_97_82), .C2 (n_96_88) );
AOI211_X1 g_85_86 (.ZN (n_85_86), .A (n_89_84), .B (n_94_84), .C1 (n_95_81), .C2 (n_97_86) );
AOI211_X1 g_83_85 (.ZN (n_83_85), .A (n_87_85), .B (n_93_82), .C1 (n_96_83), .C2 (n_98_84) );
AOI211_X1 g_81_86 (.ZN (n_81_86), .A (n_85_86), .B (n_91_83), .C1 (n_94_84), .C2 (n_97_82) );
AOI211_X1 g_79_87 (.ZN (n_79_87), .A (n_83_85), .B (n_89_84), .C1 (n_93_82), .C2 (n_95_81) );
AOI211_X1 g_77_88 (.ZN (n_77_88), .A (n_81_86), .B (n_87_85), .C1 (n_91_83), .C2 (n_96_83) );
AOI211_X1 g_75_89 (.ZN (n_75_89), .A (n_79_87), .B (n_85_86), .C1 (n_89_84), .C2 (n_94_84) );
AOI211_X1 g_73_90 (.ZN (n_73_90), .A (n_77_88), .B (n_83_85), .C1 (n_87_85), .C2 (n_93_82) );
AOI211_X1 g_71_91 (.ZN (n_71_91), .A (n_75_89), .B (n_81_86), .C1 (n_85_86), .C2 (n_91_83) );
AOI211_X1 g_69_92 (.ZN (n_69_92), .A (n_73_90), .B (n_79_87), .C1 (n_83_85), .C2 (n_89_84) );
AOI211_X1 g_71_93 (.ZN (n_71_93), .A (n_71_91), .B (n_77_88), .C1 (n_81_86), .C2 (n_87_85) );
AOI211_X1 g_73_92 (.ZN (n_73_92), .A (n_69_92), .B (n_75_89), .C1 (n_79_87), .C2 (n_85_86) );
AOI211_X1 g_74_90 (.ZN (n_74_90), .A (n_71_93), .B (n_73_90), .C1 (n_77_88), .C2 (n_83_85) );
AOI211_X1 g_76_89 (.ZN (n_76_89), .A (n_73_92), .B (n_71_91), .C1 (n_75_89), .C2 (n_81_86) );
AOI211_X1 g_78_88 (.ZN (n_78_88), .A (n_74_90), .B (n_69_92), .C1 (n_73_90), .C2 (n_79_87) );
AOI211_X1 g_80_87 (.ZN (n_80_87), .A (n_76_89), .B (n_71_93), .C1 (n_71_91), .C2 (n_77_88) );
AOI211_X1 g_82_86 (.ZN (n_82_86), .A (n_78_88), .B (n_73_92), .C1 (n_69_92), .C2 (n_75_89) );
AOI211_X1 g_84_87 (.ZN (n_84_87), .A (n_80_87), .B (n_74_90), .C1 (n_71_93), .C2 (n_73_90) );
AOI211_X1 g_82_88 (.ZN (n_82_88), .A (n_82_86), .B (n_76_89), .C1 (n_73_92), .C2 (n_71_91) );
AOI211_X1 g_80_89 (.ZN (n_80_89), .A (n_84_87), .B (n_78_88), .C1 (n_74_90), .C2 (n_69_92) );
AOI211_X1 g_78_90 (.ZN (n_78_90), .A (n_82_88), .B (n_80_87), .C1 (n_76_89), .C2 (n_71_93) );
AOI211_X1 g_76_91 (.ZN (n_76_91), .A (n_80_89), .B (n_82_86), .C1 (n_78_88), .C2 (n_73_92) );
AOI211_X1 g_74_92 (.ZN (n_74_92), .A (n_78_90), .B (n_84_87), .C1 (n_80_87), .C2 (n_74_90) );
AOI211_X1 g_72_93 (.ZN (n_72_93), .A (n_76_91), .B (n_82_88), .C1 (n_82_86), .C2 (n_76_89) );
AOI211_X1 g_70_92 (.ZN (n_70_92), .A (n_74_92), .B (n_80_89), .C1 (n_84_87), .C2 (n_78_88) );
AOI211_X1 g_68_91 (.ZN (n_68_91), .A (n_72_93), .B (n_78_90), .C1 (n_82_88), .C2 (n_80_87) );
AOI211_X1 g_66_92 (.ZN (n_66_92), .A (n_70_92), .B (n_76_91), .C1 (n_80_89), .C2 (n_82_86) );
AOI211_X1 g_64_93 (.ZN (n_64_93), .A (n_68_91), .B (n_74_92), .C1 (n_78_90), .C2 (n_84_87) );
AOI211_X1 g_62_94 (.ZN (n_62_94), .A (n_66_92), .B (n_72_93), .C1 (n_76_91), .C2 (n_82_88) );
AOI211_X1 g_61_92 (.ZN (n_61_92), .A (n_64_93), .B (n_70_92), .C1 (n_74_92), .C2 (n_80_89) );
AOI211_X1 g_60_94 (.ZN (n_60_94), .A (n_62_94), .B (n_68_91), .C1 (n_72_93), .C2 (n_78_90) );
AOI211_X1 g_58_95 (.ZN (n_58_95), .A (n_61_92), .B (n_66_92), .C1 (n_70_92), .C2 (n_76_91) );
AOI211_X1 g_59_93 (.ZN (n_59_93), .A (n_60_94), .B (n_64_93), .C1 (n_68_91), .C2 (n_74_92) );
AOI211_X1 g_57_94 (.ZN (n_57_94), .A (n_58_95), .B (n_62_94), .C1 (n_66_92), .C2 (n_72_93) );
AOI211_X1 g_56_96 (.ZN (n_56_96), .A (n_59_93), .B (n_61_92), .C1 (n_64_93), .C2 (n_70_92) );
AOI211_X1 g_57_98 (.ZN (n_57_98), .A (n_57_94), .B (n_60_94), .C1 (n_62_94), .C2 (n_68_91) );
AOI211_X1 g_58_96 (.ZN (n_58_96), .A (n_56_96), .B (n_58_95), .C1 (n_61_92), .C2 (n_66_92) );
AOI211_X1 g_60_95 (.ZN (n_60_95), .A (n_57_98), .B (n_59_93), .C1 (n_60_94), .C2 (n_64_93) );
AOI211_X1 g_59_97 (.ZN (n_59_97), .A (n_58_96), .B (n_57_94), .C1 (n_58_95), .C2 (n_62_94) );
AOI211_X1 g_61_96 (.ZN (n_61_96), .A (n_60_95), .B (n_56_96), .C1 (n_59_93), .C2 (n_61_92) );
AOI211_X1 g_59_95 (.ZN (n_59_95), .A (n_59_97), .B (n_57_98), .C1 (n_57_94), .C2 (n_60_94) );
AOI211_X1 g_58_97 (.ZN (n_58_97), .A (n_61_96), .B (n_58_96), .C1 (n_56_96), .C2 (n_58_95) );
AOI211_X1 g_60_98 (.ZN (n_60_98), .A (n_59_95), .B (n_60_95), .C1 (n_57_98), .C2 (n_59_93) );
AOI211_X1 g_61_100 (.ZN (n_61_100), .A (n_58_97), .B (n_59_97), .C1 (n_58_96), .C2 (n_57_94) );
AOI211_X1 g_59_99 (.ZN (n_59_99), .A (n_60_98), .B (n_61_96), .C1 (n_60_95), .C2 (n_56_96) );
AOI211_X1 g_60_97 (.ZN (n_60_97), .A (n_61_100), .B (n_59_95), .C1 (n_59_97), .C2 (n_57_98) );
AOI211_X1 g_62_98 (.ZN (n_62_98), .A (n_59_99), .B (n_58_97), .C1 (n_61_96), .C2 (n_58_96) );
AOI211_X1 g_63_96 (.ZN (n_63_96), .A (n_60_97), .B (n_60_98), .C1 (n_59_95), .C2 (n_60_95) );
AOI211_X1 g_64_98 (.ZN (n_64_98), .A (n_62_98), .B (n_61_100), .C1 (n_58_97), .C2 (n_59_97) );
AOI211_X1 g_65_100 (.ZN (n_65_100), .A (n_63_96), .B (n_59_99), .C1 (n_60_98), .C2 (n_61_96) );
AOI211_X1 g_66_98 (.ZN (n_66_98), .A (n_64_98), .B (n_60_97), .C1 (n_61_100), .C2 (n_59_95) );
AOI211_X1 g_67_96 (.ZN (n_67_96), .A (n_65_100), .B (n_62_98), .C1 (n_59_99), .C2 (n_58_97) );
AOI211_X1 g_65_95 (.ZN (n_65_95), .A (n_66_98), .B (n_63_96), .C1 (n_60_97), .C2 (n_60_98) );
AOI211_X1 g_66_93 (.ZN (n_66_93), .A (n_67_96), .B (n_64_98), .C1 (n_62_98), .C2 (n_61_100) );
AOI211_X1 g_64_94 (.ZN (n_64_94), .A (n_65_95), .B (n_65_100), .C1 (n_63_96), .C2 (n_59_99) );
AOI211_X1 g_65_92 (.ZN (n_65_92), .A (n_66_93), .B (n_66_98), .C1 (n_64_98), .C2 (n_60_97) );
AOI211_X1 g_63_93 (.ZN (n_63_93), .A (n_64_94), .B (n_67_96), .C1 (n_65_100), .C2 (n_62_98) );
AOI211_X1 g_61_94 (.ZN (n_61_94), .A (n_65_92), .B (n_65_95), .C1 (n_66_98), .C2 (n_63_96) );
AOI211_X1 g_60_96 (.ZN (n_60_96), .A (n_63_93), .B (n_66_93), .C1 (n_67_96), .C2 (n_64_98) );
AOI211_X1 g_62_95 (.ZN (n_62_95), .A (n_61_94), .B (n_64_94), .C1 (n_65_95), .C2 (n_65_100) );
AOI211_X1 g_63_97 (.ZN (n_63_97), .A (n_60_96), .B (n_65_92), .C1 (n_66_93), .C2 (n_66_98) );
AOI211_X1 g_61_98 (.ZN (n_61_98), .A (n_62_95), .B (n_63_93), .C1 (n_64_94), .C2 (n_67_96) );
AOI211_X1 g_62_96 (.ZN (n_62_96), .A (n_63_97), .B (n_61_94), .C1 (n_65_92), .C2 (n_65_95) );
AOI211_X1 g_64_95 (.ZN (n_64_95), .A (n_61_98), .B (n_60_96), .C1 (n_63_93), .C2 (n_66_93) );
AOI211_X1 g_66_94 (.ZN (n_66_94), .A (n_62_96), .B (n_62_95), .C1 (n_61_94), .C2 (n_64_94) );
AOI211_X1 g_68_93 (.ZN (n_68_93), .A (n_64_95), .B (n_63_97), .C1 (n_60_96), .C2 (n_65_92) );
AOI211_X1 g_70_94 (.ZN (n_70_94), .A (n_66_94), .B (n_61_98), .C1 (n_62_95), .C2 (n_63_93) );
AOI211_X1 g_71_92 (.ZN (n_71_92), .A (n_68_93), .B (n_62_96), .C1 (n_63_97), .C2 (n_61_94) );
AOI211_X1 g_69_93 (.ZN (n_69_93), .A (n_70_94), .B (n_64_95), .C1 (n_61_98), .C2 (n_60_96) );
AOI211_X1 g_67_94 (.ZN (n_67_94), .A (n_71_92), .B (n_66_94), .C1 (n_62_96), .C2 (n_62_95) );
AOI211_X1 g_66_96 (.ZN (n_66_96), .A (n_69_93), .B (n_68_93), .C1 (n_64_95), .C2 (n_63_97) );
AOI211_X1 g_64_97 (.ZN (n_64_97), .A (n_67_94), .B (n_70_94), .C1 (n_66_94), .C2 (n_61_98) );
AOI211_X1 g_63_99 (.ZN (n_63_99), .A (n_66_96), .B (n_71_92), .C1 (n_68_93), .C2 (n_62_96) );
AOI211_X1 g_62_97 (.ZN (n_62_97), .A (n_64_97), .B (n_69_93), .C1 (n_70_94), .C2 (n_64_95) );
AOI211_X1 g_63_95 (.ZN (n_63_95), .A (n_63_99), .B (n_67_94), .C1 (n_71_92), .C2 (n_66_94) );
AOI211_X1 g_65_96 (.ZN (n_65_96), .A (n_62_97), .B (n_66_96), .C1 (n_69_93), .C2 (n_68_93) );
AOI211_X1 g_67_95 (.ZN (n_67_95), .A (n_63_95), .B (n_64_97), .C1 (n_67_94), .C2 (n_70_94) );
AOI211_X1 g_65_94 (.ZN (n_65_94), .A (n_65_96), .B (n_63_99), .C1 (n_66_96), .C2 (n_71_92) );
AOI211_X1 g_67_93 (.ZN (n_67_93), .A (n_67_95), .B (n_62_97), .C1 (n_64_97), .C2 (n_69_93) );
AOI211_X1 g_68_95 (.ZN (n_68_95), .A (n_65_94), .B (n_63_95), .C1 (n_63_99), .C2 (n_67_94) );
AOI211_X1 g_67_97 (.ZN (n_67_97), .A (n_67_93), .B (n_65_96), .C1 (n_62_97), .C2 (n_66_96) );
AOI211_X1 g_65_98 (.ZN (n_65_98), .A (n_68_95), .B (n_67_95), .C1 (n_63_95), .C2 (n_64_97) );
AOI211_X1 g_64_96 (.ZN (n_64_96), .A (n_67_97), .B (n_65_94), .C1 (n_65_96), .C2 (n_63_99) );
AOI211_X1 g_66_95 (.ZN (n_66_95), .A (n_65_98), .B (n_67_93), .C1 (n_67_95), .C2 (n_62_97) );
AOI211_X1 g_68_94 (.ZN (n_68_94), .A (n_64_96), .B (n_68_95), .C1 (n_65_94), .C2 (n_63_95) );
AOI211_X1 g_70_93 (.ZN (n_70_93), .A (n_66_95), .B (n_67_97), .C1 (n_67_93), .C2 (n_65_96) );
AOI211_X1 g_72_92 (.ZN (n_72_92), .A (n_68_94), .B (n_65_98), .C1 (n_68_95), .C2 (n_67_95) );
AOI211_X1 g_74_91 (.ZN (n_74_91), .A (n_70_93), .B (n_64_96), .C1 (n_67_97), .C2 (n_65_94) );
AOI211_X1 g_76_90 (.ZN (n_76_90), .A (n_72_92), .B (n_66_95), .C1 (n_65_98), .C2 (n_67_93) );
AOI211_X1 g_78_89 (.ZN (n_78_89), .A (n_74_91), .B (n_68_94), .C1 (n_64_96), .C2 (n_68_95) );
AOI211_X1 g_80_88 (.ZN (n_80_88), .A (n_76_90), .B (n_70_93), .C1 (n_66_95), .C2 (n_67_97) );
AOI211_X1 g_82_87 (.ZN (n_82_87), .A (n_78_89), .B (n_72_92), .C1 (n_68_94), .C2 (n_65_98) );
AOI211_X1 g_84_86 (.ZN (n_84_86), .A (n_80_88), .B (n_74_91), .C1 (n_70_93), .C2 (n_64_96) );
AOI211_X1 g_83_88 (.ZN (n_83_88), .A (n_82_87), .B (n_76_90), .C1 (n_72_92), .C2 (n_66_95) );
AOI211_X1 g_85_87 (.ZN (n_85_87), .A (n_84_86), .B (n_78_89), .C1 (n_74_91), .C2 (n_68_94) );
AOI211_X1 g_84_89 (.ZN (n_84_89), .A (n_83_88), .B (n_80_88), .C1 (n_76_90), .C2 (n_70_93) );
AOI211_X1 g_83_87 (.ZN (n_83_87), .A (n_85_87), .B (n_82_87), .C1 (n_78_89), .C2 (n_72_92) );
AOI211_X1 g_81_88 (.ZN (n_81_88), .A (n_84_89), .B (n_84_86), .C1 (n_80_88), .C2 (n_74_91) );
AOI211_X1 g_79_89 (.ZN (n_79_89), .A (n_83_87), .B (n_83_88), .C1 (n_82_87), .C2 (n_76_90) );
AOI211_X1 g_77_90 (.ZN (n_77_90), .A (n_81_88), .B (n_85_87), .C1 (n_84_86), .C2 (n_78_89) );
AOI211_X1 g_75_91 (.ZN (n_75_91), .A (n_79_89), .B (n_84_89), .C1 (n_83_88), .C2 (n_80_88) );
AOI211_X1 g_74_93 (.ZN (n_74_93), .A (n_77_90), .B (n_83_87), .C1 (n_85_87), .C2 (n_82_87) );
AOI211_X1 g_76_92 (.ZN (n_76_92), .A (n_75_91), .B (n_81_88), .C1 (n_84_89), .C2 (n_84_86) );
AOI211_X1 g_78_91 (.ZN (n_78_91), .A (n_74_93), .B (n_79_89), .C1 (n_83_87), .C2 (n_83_88) );
AOI211_X1 g_80_90 (.ZN (n_80_90), .A (n_76_92), .B (n_77_90), .C1 (n_81_88), .C2 (n_85_87) );
AOI211_X1 g_82_89 (.ZN (n_82_89), .A (n_78_91), .B (n_75_91), .C1 (n_79_89), .C2 (n_84_89) );
AOI211_X1 g_84_88 (.ZN (n_84_88), .A (n_80_90), .B (n_74_93), .C1 (n_77_90), .C2 (n_83_87) );
AOI211_X1 g_86_87 (.ZN (n_86_87), .A (n_82_89), .B (n_76_92), .C1 (n_75_91), .C2 (n_81_88) );
AOI211_X1 g_88_86 (.ZN (n_88_86), .A (n_84_88), .B (n_78_91), .C1 (n_74_93), .C2 (n_79_89) );
AOI211_X1 g_90_85 (.ZN (n_90_85), .A (n_86_87), .B (n_80_90), .C1 (n_76_92), .C2 (n_77_90) );
AOI211_X1 g_92_84 (.ZN (n_92_84), .A (n_88_86), .B (n_82_89), .C1 (n_78_91), .C2 (n_75_91) );
AOI211_X1 g_94_83 (.ZN (n_94_83), .A (n_90_85), .B (n_84_88), .C1 (n_80_90), .C2 (n_74_93) );
AOI211_X1 g_96_84 (.ZN (n_96_84), .A (n_92_84), .B (n_86_87), .C1 (n_82_89), .C2 (n_76_92) );
AOI211_X1 g_95_86 (.ZN (n_95_86), .A (n_94_83), .B (n_88_86), .C1 (n_84_88), .C2 (n_78_91) );
AOI211_X1 g_93_85 (.ZN (n_93_85), .A (n_96_84), .B (n_90_85), .C1 (n_86_87), .C2 (n_80_90) );
AOI211_X1 g_91_86 (.ZN (n_91_86), .A (n_95_86), .B (n_92_84), .C1 (n_88_86), .C2 (n_82_89) );
AOI211_X1 g_89_87 (.ZN (n_89_87), .A (n_93_85), .B (n_94_83), .C1 (n_90_85), .C2 (n_84_88) );
AOI211_X1 g_87_88 (.ZN (n_87_88), .A (n_91_86), .B (n_96_84), .C1 (n_92_84), .C2 (n_86_87) );
AOI211_X1 g_85_89 (.ZN (n_85_89), .A (n_89_87), .B (n_95_86), .C1 (n_94_83), .C2 (n_88_86) );
AOI211_X1 g_83_90 (.ZN (n_83_90), .A (n_87_88), .B (n_93_85), .C1 (n_96_84), .C2 (n_90_85) );
AOI211_X1 g_81_89 (.ZN (n_81_89), .A (n_85_89), .B (n_91_86), .C1 (n_95_86), .C2 (n_92_84) );
AOI211_X1 g_79_90 (.ZN (n_79_90), .A (n_83_90), .B (n_89_87), .C1 (n_93_85), .C2 (n_94_83) );
AOI211_X1 g_77_91 (.ZN (n_77_91), .A (n_81_89), .B (n_87_88), .C1 (n_91_86), .C2 (n_96_84) );
AOI211_X1 g_75_92 (.ZN (n_75_92), .A (n_79_90), .B (n_85_89), .C1 (n_89_87), .C2 (n_95_86) );
AOI211_X1 g_73_93 (.ZN (n_73_93), .A (n_77_91), .B (n_83_90), .C1 (n_87_88), .C2 (n_93_85) );
AOI211_X1 g_71_94 (.ZN (n_71_94), .A (n_75_92), .B (n_81_89), .C1 (n_85_89), .C2 (n_91_86) );
AOI211_X1 g_69_95 (.ZN (n_69_95), .A (n_73_93), .B (n_79_90), .C1 (n_83_90), .C2 (n_89_87) );
AOI211_X1 g_68_97 (.ZN (n_68_97), .A (n_71_94), .B (n_77_91), .C1 (n_81_89), .C2 (n_87_88) );
AOI211_X1 g_67_99 (.ZN (n_67_99), .A (n_69_95), .B (n_75_92), .C1 (n_79_90), .C2 (n_85_89) );
AOI211_X1 g_66_97 (.ZN (n_66_97), .A (n_68_97), .B (n_73_93), .C1 (n_77_91), .C2 (n_83_90) );
AOI211_X1 g_68_98 (.ZN (n_68_98), .A (n_67_99), .B (n_71_94), .C1 (n_75_92), .C2 (n_81_89) );
AOI211_X1 g_69_100 (.ZN (n_69_100), .A (n_66_97), .B (n_69_95), .C1 (n_73_93), .C2 (n_79_90) );
AOI211_X1 g_70_98 (.ZN (n_70_98), .A (n_68_98), .B (n_68_97), .C1 (n_71_94), .C2 (n_77_91) );
AOI211_X1 g_69_96 (.ZN (n_69_96), .A (n_69_100), .B (n_67_99), .C1 (n_69_95), .C2 (n_75_92) );
AOI211_X1 g_71_95 (.ZN (n_71_95), .A (n_70_98), .B (n_66_97), .C1 (n_68_97), .C2 (n_73_93) );
AOI211_X1 g_69_94 (.ZN (n_69_94), .A (n_69_96), .B (n_68_98), .C1 (n_67_99), .C2 (n_71_94) );
AOI211_X1 g_68_96 (.ZN (n_68_96), .A (n_71_95), .B (n_69_100), .C1 (n_66_97), .C2 (n_69_95) );
AOI211_X1 g_70_95 (.ZN (n_70_95), .A (n_69_94), .B (n_70_98), .C1 (n_68_98), .C2 (n_68_97) );
AOI211_X1 g_72_94 (.ZN (n_72_94), .A (n_68_96), .B (n_69_96), .C1 (n_69_100), .C2 (n_67_99) );
AOI211_X1 g_71_96 (.ZN (n_71_96), .A (n_70_95), .B (n_71_95), .C1 (n_70_98), .C2 (n_66_97) );
AOI211_X1 g_73_95 (.ZN (n_73_95), .A (n_72_94), .B (n_69_94), .C1 (n_69_96), .C2 (n_68_98) );
AOI211_X1 g_75_94 (.ZN (n_75_94), .A (n_71_96), .B (n_68_96), .C1 (n_71_95), .C2 (n_69_100) );
AOI211_X1 g_77_93 (.ZN (n_77_93), .A (n_73_95), .B (n_70_95), .C1 (n_69_94), .C2 (n_70_98) );
AOI211_X1 g_79_92 (.ZN (n_79_92), .A (n_75_94), .B (n_72_94), .C1 (n_68_96), .C2 (n_69_96) );
AOI211_X1 g_81_91 (.ZN (n_81_91), .A (n_77_93), .B (n_71_96), .C1 (n_70_95), .C2 (n_71_95) );
AOI211_X1 g_80_93 (.ZN (n_80_93), .A (n_79_92), .B (n_73_95), .C1 (n_72_94), .C2 (n_69_94) );
AOI211_X1 g_79_91 (.ZN (n_79_91), .A (n_81_91), .B (n_75_94), .C1 (n_71_96), .C2 (n_68_96) );
AOI211_X1 g_81_90 (.ZN (n_81_90), .A (n_80_93), .B (n_77_93), .C1 (n_73_95), .C2 (n_70_95) );
AOI211_X1 g_83_89 (.ZN (n_83_89), .A (n_79_91), .B (n_79_92), .C1 (n_75_94), .C2 (n_72_94) );
AOI211_X1 g_85_88 (.ZN (n_85_88), .A (n_81_90), .B (n_81_91), .C1 (n_77_93), .C2 (n_71_96) );
AOI211_X1 g_84_90 (.ZN (n_84_90), .A (n_83_89), .B (n_80_93), .C1 (n_79_92), .C2 (n_73_95) );
AOI211_X1 g_86_89 (.ZN (n_86_89), .A (n_85_88), .B (n_79_91), .C1 (n_81_91), .C2 (n_75_94) );
AOI211_X1 g_88_88 (.ZN (n_88_88), .A (n_84_90), .B (n_81_90), .C1 (n_80_93), .C2 (n_77_93) );
AOI211_X1 g_89_86 (.ZN (n_89_86), .A (n_86_89), .B (n_83_89), .C1 (n_79_91), .C2 (n_79_92) );
AOI211_X1 g_91_85 (.ZN (n_91_85), .A (n_88_88), .B (n_85_88), .C1 (n_81_90), .C2 (n_81_91) );
AOI211_X1 g_93_84 (.ZN (n_93_84), .A (n_89_86), .B (n_84_90), .C1 (n_83_89), .C2 (n_80_93) );
AOI211_X1 g_95_83 (.ZN (n_95_83), .A (n_91_85), .B (n_86_89), .C1 (n_85_88), .C2 (n_79_91) );
AOI211_X1 g_96_85 (.ZN (n_96_85), .A (n_93_84), .B (n_88_88), .C1 (n_84_90), .C2 (n_81_90) );
AOI211_X1 g_98_86 (.ZN (n_98_86), .A (n_95_83), .B (n_89_86), .C1 (n_86_89), .C2 (n_83_89) );
AOI211_X1 g_97_84 (.ZN (n_97_84), .A (n_96_85), .B (n_91_85), .C1 (n_88_88), .C2 (n_85_88) );
AOI211_X1 g_95_85 (.ZN (n_95_85), .A (n_98_86), .B (n_93_84), .C1 (n_89_86), .C2 (n_84_90) );
AOI211_X1 g_96_87 (.ZN (n_96_87), .A (n_97_84), .B (n_95_83), .C1 (n_91_85), .C2 (n_86_89) );
AOI211_X1 g_94_86 (.ZN (n_94_86), .A (n_95_85), .B (n_96_85), .C1 (n_93_84), .C2 (n_88_88) );
AOI211_X1 g_92_85 (.ZN (n_92_85), .A (n_96_87), .B (n_98_86), .C1 (n_95_83), .C2 (n_89_86) );
AOI211_X1 g_90_86 (.ZN (n_90_86), .A (n_94_86), .B (n_97_84), .C1 (n_96_85), .C2 (n_91_85) );
AOI211_X1 g_88_87 (.ZN (n_88_87), .A (n_92_85), .B (n_95_85), .C1 (n_98_86), .C2 (n_93_84) );
AOI211_X1 g_86_88 (.ZN (n_86_88), .A (n_90_86), .B (n_96_87), .C1 (n_97_84), .C2 (n_95_83) );
AOI211_X1 g_85_90 (.ZN (n_85_90), .A (n_88_87), .B (n_94_86), .C1 (n_95_85), .C2 (n_96_85) );
AOI211_X1 g_87_89 (.ZN (n_87_89), .A (n_86_88), .B (n_92_85), .C1 (n_96_87), .C2 (n_98_86) );
AOI211_X1 g_89_88 (.ZN (n_89_88), .A (n_85_90), .B (n_90_86), .C1 (n_94_86), .C2 (n_97_84) );
AOI211_X1 g_91_87 (.ZN (n_91_87), .A (n_87_89), .B (n_88_87), .C1 (n_92_85), .C2 (n_95_85) );
AOI211_X1 g_93_86 (.ZN (n_93_86), .A (n_89_88), .B (n_86_88), .C1 (n_90_86), .C2 (n_96_87) );
AOI211_X1 g_94_88 (.ZN (n_94_88), .A (n_91_87), .B (n_85_90), .C1 (n_88_87), .C2 (n_94_86) );
AOI211_X1 g_92_87 (.ZN (n_92_87), .A (n_93_86), .B (n_87_89), .C1 (n_86_88), .C2 (n_92_85) );
AOI211_X1 g_90_88 (.ZN (n_90_88), .A (n_94_88), .B (n_89_88), .C1 (n_85_90), .C2 (n_90_86) );
AOI211_X1 g_88_89 (.ZN (n_88_89), .A (n_92_87), .B (n_91_87), .C1 (n_87_89), .C2 (n_88_87) );
AOI211_X1 g_86_90 (.ZN (n_86_90), .A (n_90_88), .B (n_93_86), .C1 (n_89_88), .C2 (n_86_88) );
AOI211_X1 g_84_91 (.ZN (n_84_91), .A (n_88_89), .B (n_94_88), .C1 (n_91_87), .C2 (n_85_90) );
AOI211_X1 g_82_90 (.ZN (n_82_90), .A (n_86_90), .B (n_92_87), .C1 (n_93_86), .C2 (n_87_89) );
AOI211_X1 g_80_91 (.ZN (n_80_91), .A (n_84_91), .B (n_90_88), .C1 (n_94_88), .C2 (n_89_88) );
AOI211_X1 g_78_92 (.ZN (n_78_92), .A (n_82_90), .B (n_88_89), .C1 (n_92_87), .C2 (n_91_87) );
AOI211_X1 g_76_93 (.ZN (n_76_93), .A (n_80_91), .B (n_86_90), .C1 (n_90_88), .C2 (n_93_86) );
AOI211_X1 g_74_94 (.ZN (n_74_94), .A (n_78_92), .B (n_84_91), .C1 (n_88_89), .C2 (n_94_88) );
AOI211_X1 g_72_95 (.ZN (n_72_95), .A (n_76_93), .B (n_82_90), .C1 (n_86_90), .C2 (n_92_87) );
AOI211_X1 g_70_96 (.ZN (n_70_96), .A (n_74_94), .B (n_80_91), .C1 (n_84_91), .C2 (n_90_88) );
AOI211_X1 g_69_98 (.ZN (n_69_98), .A (n_72_95), .B (n_78_92), .C1 (n_82_90), .C2 (n_88_89) );
AOI211_X1 g_71_97 (.ZN (n_71_97), .A (n_70_96), .B (n_76_93), .C1 (n_80_91), .C2 (n_86_90) );
AOI211_X1 g_73_96 (.ZN (n_73_96), .A (n_69_98), .B (n_74_94), .C1 (n_78_92), .C2 (n_84_91) );
AOI211_X1 g_72_98 (.ZN (n_72_98), .A (n_71_97), .B (n_72_95), .C1 (n_76_93), .C2 (n_82_90) );
AOI211_X1 g_70_97 (.ZN (n_70_97), .A (n_73_96), .B (n_70_96), .C1 (n_74_94), .C2 (n_80_91) );
AOI211_X1 g_71_99 (.ZN (n_71_99), .A (n_72_98), .B (n_69_98), .C1 (n_72_95), .C2 (n_78_92) );
AOI211_X1 g_72_97 (.ZN (n_72_97), .A (n_70_97), .B (n_71_97), .C1 (n_70_96), .C2 (n_76_93) );
AOI211_X1 g_74_98 (.ZN (n_74_98), .A (n_71_99), .B (n_73_96), .C1 (n_69_98), .C2 (n_74_94) );
AOI211_X1 g_73_100 (.ZN (n_73_100), .A (n_72_97), .B (n_72_98), .C1 (n_71_97), .C2 (n_72_95) );
AOI211_X1 g_75_99 (.ZN (n_75_99), .A (n_74_98), .B (n_70_97), .C1 (n_73_96), .C2 (n_70_96) );
AOI211_X1 g_73_98 (.ZN (n_73_98), .A (n_73_100), .B (n_71_99), .C1 (n_72_98), .C2 (n_69_98) );
AOI211_X1 g_74_96 (.ZN (n_74_96), .A (n_75_99), .B (n_72_97), .C1 (n_70_97), .C2 (n_71_97) );
AOI211_X1 g_73_94 (.ZN (n_73_94), .A (n_73_98), .B (n_74_98), .C1 (n_71_99), .C2 (n_73_96) );
AOI211_X1 g_72_96 (.ZN (n_72_96), .A (n_74_96), .B (n_73_100), .C1 (n_72_97), .C2 (n_72_98) );
AOI211_X1 g_74_97 (.ZN (n_74_97), .A (n_73_94), .B (n_75_99), .C1 (n_74_98), .C2 (n_70_97) );
AOI211_X1 g_75_95 (.ZN (n_75_95), .A (n_72_96), .B (n_73_98), .C1 (n_73_100), .C2 (n_71_99) );
AOI211_X1 g_76_97 (.ZN (n_76_97), .A (n_74_97), .B (n_74_96), .C1 (n_75_99), .C2 (n_72_97) );
AOI211_X1 g_78_98 (.ZN (n_78_98), .A (n_75_95), .B (n_73_94), .C1 (n_73_98), .C2 (n_74_98) );
AOI211_X1 g_77_100 (.ZN (n_77_100), .A (n_76_97), .B (n_72_96), .C1 (n_74_96), .C2 (n_73_100) );
AOI211_X1 g_76_98 (.ZN (n_76_98), .A (n_78_98), .B (n_74_97), .C1 (n_73_94), .C2 (n_75_99) );
AOI211_X1 g_75_96 (.ZN (n_75_96), .A (n_77_100), .B (n_75_95), .C1 (n_72_96), .C2 (n_73_98) );
AOI211_X1 g_77_95 (.ZN (n_77_95), .A (n_76_98), .B (n_76_97), .C1 (n_74_97), .C2 (n_74_96) );
AOI211_X1 g_78_93 (.ZN (n_78_93), .A (n_75_96), .B (n_78_98), .C1 (n_75_95), .C2 (n_73_94) );
AOI211_X1 g_80_92 (.ZN (n_80_92), .A (n_77_95), .B (n_77_100), .C1 (n_76_97), .C2 (n_72_96) );
AOI211_X1 g_82_91 (.ZN (n_82_91), .A (n_78_93), .B (n_76_98), .C1 (n_78_98), .C2 (n_74_97) );
AOI211_X1 g_81_93 (.ZN (n_81_93), .A (n_80_92), .B (n_75_96), .C1 (n_77_100), .C2 (n_75_95) );
AOI211_X1 g_79_94 (.ZN (n_79_94), .A (n_82_91), .B (n_77_95), .C1 (n_76_98), .C2 (n_76_97) );
AOI211_X1 g_78_96 (.ZN (n_78_96), .A (n_81_93), .B (n_78_93), .C1 (n_75_96), .C2 (n_78_98) );
AOI211_X1 g_76_95 (.ZN (n_76_95), .A (n_79_94), .B (n_80_92), .C1 (n_77_95), .C2 (n_77_100) );
AOI211_X1 g_75_93 (.ZN (n_75_93), .A (n_78_96), .B (n_82_91), .C1 (n_78_93), .C2 (n_76_98) );
AOI211_X1 g_77_92 (.ZN (n_77_92), .A (n_76_95), .B (n_81_93), .C1 (n_80_92), .C2 (n_75_96) );
AOI211_X1 g_76_94 (.ZN (n_76_94), .A (n_75_93), .B (n_79_94), .C1 (n_82_91), .C2 (n_77_95) );
AOI211_X1 g_74_95 (.ZN (n_74_95), .A (n_77_92), .B (n_78_96), .C1 (n_81_93), .C2 (n_78_93) );
AOI211_X1 g_75_97 (.ZN (n_75_97), .A (n_76_94), .B (n_76_95), .C1 (n_79_94), .C2 (n_80_92) );
AOI211_X1 g_77_96 (.ZN (n_77_96), .A (n_74_95), .B (n_75_93), .C1 (n_78_96), .C2 (n_82_91) );
AOI211_X1 g_78_94 (.ZN (n_78_94), .A (n_75_97), .B (n_77_92), .C1 (n_76_95), .C2 (n_81_93) );
AOI211_X1 g_79_96 (.ZN (n_79_96), .A (n_77_96), .B (n_76_94), .C1 (n_75_93), .C2 (n_79_94) );
AOI211_X1 g_80_98 (.ZN (n_80_98), .A (n_78_94), .B (n_74_95), .C1 (n_77_92), .C2 (n_78_96) );
AOI211_X1 g_82_97 (.ZN (n_82_97), .A (n_79_96), .B (n_75_97), .C1 (n_76_94), .C2 (n_76_95) );
AOI211_X1 g_81_95 (.ZN (n_81_95), .A (n_80_98), .B (n_77_96), .C1 (n_74_95), .C2 (n_75_93) );
AOI211_X1 g_80_97 (.ZN (n_80_97), .A (n_82_97), .B (n_78_94), .C1 (n_75_97), .C2 (n_77_92) );
AOI211_X1 g_79_99 (.ZN (n_79_99), .A (n_81_95), .B (n_79_96), .C1 (n_77_96), .C2 (n_76_94) );
AOI211_X1 g_77_98 (.ZN (n_77_98), .A (n_80_97), .B (n_80_98), .C1 (n_78_94), .C2 (n_74_95) );
AOI211_X1 g_76_96 (.ZN (n_76_96), .A (n_79_99), .B (n_82_97), .C1 (n_79_96), .C2 (n_75_97) );
AOI211_X1 g_77_94 (.ZN (n_77_94), .A (n_77_98), .B (n_81_95), .C1 (n_80_98), .C2 (n_77_96) );
AOI211_X1 g_79_95 (.ZN (n_79_95), .A (n_76_96), .B (n_80_97), .C1 (n_82_97), .C2 (n_78_94) );
AOI211_X1 g_78_97 (.ZN (n_78_97), .A (n_77_94), .B (n_79_99), .C1 (n_81_95), .C2 (n_79_96) );
AOI211_X1 g_80_96 (.ZN (n_80_96), .A (n_79_95), .B (n_77_98), .C1 (n_80_97), .C2 (n_80_98) );
AOI211_X1 g_78_95 (.ZN (n_78_95), .A (n_78_97), .B (n_76_96), .C1 (n_79_99), .C2 (n_82_97) );
AOI211_X1 g_79_93 (.ZN (n_79_93), .A (n_80_96), .B (n_77_94), .C1 (n_77_98), .C2 (n_81_95) );
AOI211_X1 g_80_95 (.ZN (n_80_95), .A (n_78_95), .B (n_79_95), .C1 (n_76_96), .C2 (n_80_97) );
AOI211_X1 g_79_97 (.ZN (n_79_97), .A (n_79_93), .B (n_78_97), .C1 (n_77_94), .C2 (n_79_99) );
AOI211_X1 g_81_98 (.ZN (n_81_98), .A (n_80_95), .B (n_80_96), .C1 (n_79_95), .C2 (n_77_98) );
AOI211_X1 g_83_97 (.ZN (n_83_97), .A (n_79_97), .B (n_78_95), .C1 (n_78_97), .C2 (n_76_96) );
AOI211_X1 g_81_96 (.ZN (n_81_96), .A (n_81_98), .B (n_79_93), .C1 (n_80_96), .C2 (n_77_94) );
AOI211_X1 g_80_94 (.ZN (n_80_94), .A (n_83_97), .B (n_80_95), .C1 (n_78_95), .C2 (n_79_95) );
AOI211_X1 g_81_92 (.ZN (n_81_92), .A (n_81_96), .B (n_79_97), .C1 (n_79_93), .C2 (n_78_97) );
AOI211_X1 g_83_91 (.ZN (n_83_91), .A (n_80_94), .B (n_81_98), .C1 (n_80_95), .C2 (n_80_96) );
AOI211_X1 g_82_93 (.ZN (n_82_93), .A (n_81_92), .B (n_83_97), .C1 (n_79_97), .C2 (n_78_95) );
AOI211_X1 g_84_92 (.ZN (n_84_92), .A (n_83_91), .B (n_81_96), .C1 (n_81_98), .C2 (n_79_93) );
AOI211_X1 g_86_91 (.ZN (n_86_91), .A (n_82_93), .B (n_80_94), .C1 (n_83_97), .C2 (n_80_95) );
AOI211_X1 g_88_90 (.ZN (n_88_90), .A (n_84_92), .B (n_81_92), .C1 (n_81_96), .C2 (n_79_97) );
AOI211_X1 g_90_89 (.ZN (n_90_89), .A (n_86_91), .B (n_83_91), .C1 (n_80_94), .C2 (n_81_98) );
AOI211_X1 g_92_88 (.ZN (n_92_88), .A (n_88_90), .B (n_82_93), .C1 (n_81_92), .C2 (n_83_97) );
AOI211_X1 g_90_87 (.ZN (n_90_87), .A (n_90_89), .B (n_84_92), .C1 (n_83_91), .C2 (n_81_96) );
AOI211_X1 g_92_86 (.ZN (n_92_86), .A (n_92_88), .B (n_86_91), .C1 (n_82_93), .C2 (n_80_94) );
AOI211_X1 g_94_85 (.ZN (n_94_85), .A (n_90_87), .B (n_88_90), .C1 (n_84_92), .C2 (n_81_92) );
AOI211_X1 g_95_87 (.ZN (n_95_87), .A (n_92_86), .B (n_90_89), .C1 (n_86_91), .C2 (n_83_91) );
AOI211_X1 g_97_88 (.ZN (n_97_88), .A (n_94_85), .B (n_92_88), .C1 (n_88_90), .C2 (n_82_93) );
AOI211_X1 g_96_86 (.ZN (n_96_86), .A (n_95_87), .B (n_90_87), .C1 (n_90_89), .C2 (n_84_92) );
AOI211_X1 g_94_87 (.ZN (n_94_87), .A (n_97_88), .B (n_92_86), .C1 (n_92_88), .C2 (n_86_91) );
AOI211_X1 g_95_89 (.ZN (n_95_89), .A (n_96_86), .B (n_94_85), .C1 (n_90_87), .C2 (n_88_90) );
AOI211_X1 g_93_88 (.ZN (n_93_88), .A (n_94_87), .B (n_95_87), .C1 (n_92_86), .C2 (n_90_89) );
AOI211_X1 g_91_89 (.ZN (n_91_89), .A (n_95_89), .B (n_97_88), .C1 (n_94_85), .C2 (n_92_88) );
AOI211_X1 g_93_90 (.ZN (n_93_90), .A (n_93_88), .B (n_96_86), .C1 (n_95_87), .C2 (n_90_87) );
AOI211_X1 g_92_92 (.ZN (n_92_92), .A (n_91_89), .B (n_94_87), .C1 (n_97_88), .C2 (n_92_86) );
AOI211_X1 g_94_91 (.ZN (n_94_91), .A (n_93_90), .B (n_95_89), .C1 (n_96_86), .C2 (n_94_85) );
AOI211_X1 g_96_90 (.ZN (n_96_90), .A (n_92_92), .B (n_93_88), .C1 (n_94_87), .C2 (n_95_87) );
AOI211_X1 g_95_88 (.ZN (n_95_88), .A (n_94_91), .B (n_91_89), .C1 (n_95_89), .C2 (n_97_88) );
AOI211_X1 g_93_87 (.ZN (n_93_87), .A (n_96_90), .B (n_93_90), .C1 (n_93_88), .C2 (n_96_86) );
AOI211_X1 g_94_89 (.ZN (n_94_89), .A (n_95_88), .B (n_92_92), .C1 (n_91_89), .C2 (n_94_87) );
AOI211_X1 g_92_90 (.ZN (n_92_90), .A (n_93_87), .B (n_94_91), .C1 (n_93_90), .C2 (n_95_89) );
AOI211_X1 g_91_88 (.ZN (n_91_88), .A (n_94_89), .B (n_96_90), .C1 (n_92_92), .C2 (n_93_88) );
AOI211_X1 g_93_89 (.ZN (n_93_89), .A (n_92_90), .B (n_95_88), .C1 (n_94_91), .C2 (n_91_89) );
AOI211_X1 g_91_90 (.ZN (n_91_90), .A (n_91_88), .B (n_93_87), .C1 (n_96_90), .C2 (n_93_90) );
AOI211_X1 g_89_89 (.ZN (n_89_89), .A (n_93_89), .B (n_94_89), .C1 (n_95_88), .C2 (n_92_92) );
AOI211_X1 g_90_91 (.ZN (n_90_91), .A (n_91_90), .B (n_92_90), .C1 (n_93_87), .C2 (n_94_91) );
AOI211_X1 g_91_93 (.ZN (n_91_93), .A (n_89_89), .B (n_91_88), .C1 (n_94_89), .C2 (n_96_90) );
AOI211_X1 g_93_92 (.ZN (n_93_92), .A (n_90_91), .B (n_93_89), .C1 (n_92_90), .C2 (n_95_88) );
AOI211_X1 g_94_90 (.ZN (n_94_90), .A (n_91_93), .B (n_91_90), .C1 (n_91_88), .C2 (n_93_87) );
AOI211_X1 g_92_89 (.ZN (n_92_89), .A (n_93_92), .B (n_89_89), .C1 (n_93_89), .C2 (n_94_89) );
AOI211_X1 g_93_91 (.ZN (n_93_91), .A (n_94_90), .B (n_90_91), .C1 (n_91_90), .C2 (n_92_90) );
AOI211_X1 g_95_92 (.ZN (n_95_92), .A (n_92_89), .B (n_91_93), .C1 (n_89_89), .C2 (n_91_88) );
AOI211_X1 g_94_94 (.ZN (n_94_94), .A (n_93_91), .B (n_93_92), .C1 (n_90_91), .C2 (n_93_89) );
AOI211_X1 g_92_93 (.ZN (n_92_93), .A (n_95_92), .B (n_94_90), .C1 (n_91_93), .C2 (n_91_90) );
AOI211_X1 g_91_91 (.ZN (n_91_91), .A (n_94_94), .B (n_92_89), .C1 (n_93_92), .C2 (n_89_89) );
AOI211_X1 g_89_90 (.ZN (n_89_90), .A (n_92_93), .B (n_93_91), .C1 (n_94_90), .C2 (n_90_91) );
AOI211_X1 g_87_91 (.ZN (n_87_91), .A (n_91_91), .B (n_95_92), .C1 (n_92_89), .C2 (n_91_93) );
AOI211_X1 g_85_92 (.ZN (n_85_92), .A (n_89_90), .B (n_94_94), .C1 (n_93_91), .C2 (n_93_92) );
AOI211_X1 g_83_93 (.ZN (n_83_93), .A (n_87_91), .B (n_92_93), .C1 (n_95_92), .C2 (n_94_90) );
AOI211_X1 g_82_95 (.ZN (n_82_95), .A (n_85_92), .B (n_91_91), .C1 (n_94_94), .C2 (n_92_89) );
AOI211_X1 g_84_96 (.ZN (n_84_96), .A (n_83_93), .B (n_89_90), .C1 (n_92_93), .C2 (n_93_91) );
AOI211_X1 g_86_95 (.ZN (n_86_95), .A (n_82_95), .B (n_87_91), .C1 (n_91_91), .C2 (n_95_92) );
AOI211_X1 g_84_94 (.ZN (n_84_94), .A (n_84_96), .B (n_85_92), .C1 (n_89_90), .C2 (n_94_94) );
AOI211_X1 g_83_92 (.ZN (n_83_92), .A (n_86_95), .B (n_83_93), .C1 (n_87_91), .C2 (n_92_93) );
AOI211_X1 g_82_94 (.ZN (n_82_94), .A (n_84_94), .B (n_82_95), .C1 (n_85_92), .C2 (n_91_91) );
AOI211_X1 g_84_95 (.ZN (n_84_95), .A (n_83_92), .B (n_84_96), .C1 (n_83_93), .C2 (n_89_90) );
AOI211_X1 g_85_93 (.ZN (n_85_93), .A (n_82_94), .B (n_86_95), .C1 (n_82_95), .C2 (n_87_91) );
AOI211_X1 g_83_94 (.ZN (n_83_94), .A (n_84_95), .B (n_84_94), .C1 (n_84_96), .C2 (n_85_92) );
AOI211_X1 g_82_92 (.ZN (n_82_92), .A (n_85_93), .B (n_83_92), .C1 (n_86_95), .C2 (n_83_93) );
AOI211_X1 g_81_94 (.ZN (n_81_94), .A (n_83_94), .B (n_82_94), .C1 (n_84_94), .C2 (n_82_95) );
AOI211_X1 g_82_96 (.ZN (n_82_96), .A (n_82_92), .B (n_84_95), .C1 (n_83_92), .C2 (n_84_96) );
AOI211_X1 g_84_97 (.ZN (n_84_97), .A (n_81_94), .B (n_85_93), .C1 (n_82_94), .C2 (n_86_95) );
AOI211_X1 g_85_95 (.ZN (n_85_95), .A (n_82_96), .B (n_83_94), .C1 (n_84_95), .C2 (n_84_94) );
AOI211_X1 g_86_93 (.ZN (n_86_93), .A (n_84_97), .B (n_82_92), .C1 (n_85_93), .C2 (n_83_92) );
AOI211_X1 g_85_91 (.ZN (n_85_91), .A (n_85_95), .B (n_81_94), .C1 (n_83_94), .C2 (n_82_94) );
AOI211_X1 g_87_90 (.ZN (n_87_90), .A (n_86_93), .B (n_82_96), .C1 (n_82_92), .C2 (n_84_95) );
AOI211_X1 g_88_92 (.ZN (n_88_92), .A (n_85_91), .B (n_84_97), .C1 (n_81_94), .C2 (n_85_93) );
AOI211_X1 g_90_93 (.ZN (n_90_93), .A (n_87_90), .B (n_85_95), .C1 (n_82_96), .C2 (n_83_94) );
AOI211_X1 g_88_94 (.ZN (n_88_94), .A (n_88_92), .B (n_86_93), .C1 (n_84_97), .C2 (n_82_92) );
AOI211_X1 g_89_92 (.ZN (n_89_92), .A (n_90_93), .B (n_85_91), .C1 (n_85_95), .C2 (n_81_94) );
AOI211_X1 g_90_90 (.ZN (n_90_90), .A (n_88_94), .B (n_87_90), .C1 (n_86_93), .C2 (n_82_96) );
AOI211_X1 g_92_91 (.ZN (n_92_91), .A (n_89_92), .B (n_88_92), .C1 (n_85_91), .C2 (n_84_97) );
AOI211_X1 g_93_93 (.ZN (n_93_93), .A (n_90_90), .B (n_90_93), .C1 (n_87_90), .C2 (n_85_95) );
AOI211_X1 g_92_95 (.ZN (n_92_95), .A (n_92_91), .B (n_88_94), .C1 (n_88_92), .C2 (n_86_93) );
AOI211_X1 g_90_94 (.ZN (n_90_94), .A (n_93_93), .B (n_89_92), .C1 (n_90_93), .C2 (n_85_91) );
AOI211_X1 g_91_92 (.ZN (n_91_92), .A (n_92_95), .B (n_90_90), .C1 (n_88_94), .C2 (n_87_90) );
AOI211_X1 g_89_91 (.ZN (n_89_91), .A (n_90_94), .B (n_92_91), .C1 (n_89_92), .C2 (n_88_92) );
AOI211_X1 g_87_92 (.ZN (n_87_92), .A (n_91_92), .B (n_93_93), .C1 (n_90_90), .C2 (n_90_93) );
AOI211_X1 g_86_94 (.ZN (n_86_94), .A (n_89_91), .B (n_92_95), .C1 (n_92_91), .C2 (n_88_94) );
AOI211_X1 g_84_93 (.ZN (n_84_93), .A (n_87_92), .B (n_90_94), .C1 (n_93_93), .C2 (n_89_92) );
AOI211_X1 g_83_95 (.ZN (n_83_95), .A (n_86_94), .B (n_91_92), .C1 (n_92_95), .C2 (n_90_90) );
AOI211_X1 g_85_96 (.ZN (n_85_96), .A (n_84_93), .B (n_89_91), .C1 (n_90_94), .C2 (n_92_91) );
AOI211_X1 g_87_95 (.ZN (n_87_95), .A (n_83_95), .B (n_87_92), .C1 (n_91_92), .C2 (n_93_93) );
AOI211_X1 g_89_94 (.ZN (n_89_94), .A (n_85_96), .B (n_86_94), .C1 (n_89_91), .C2 (n_92_95) );
AOI211_X1 g_90_92 (.ZN (n_90_92), .A (n_87_95), .B (n_84_93), .C1 (n_87_92), .C2 (n_90_94) );
AOI211_X1 g_88_93 (.ZN (n_88_93), .A (n_89_94), .B (n_83_95), .C1 (n_86_94), .C2 (n_91_92) );
AOI211_X1 g_86_92 (.ZN (n_86_92), .A (n_90_92), .B (n_85_96), .C1 (n_84_93), .C2 (n_89_91) );
AOI211_X1 g_88_91 (.ZN (n_88_91), .A (n_88_93), .B (n_87_95), .C1 (n_83_95), .C2 (n_87_92) );
AOI211_X1 g_87_93 (.ZN (n_87_93), .A (n_86_92), .B (n_89_94), .C1 (n_85_96), .C2 (n_86_94) );
AOI211_X1 g_85_94 (.ZN (n_85_94), .A (n_88_91), .B (n_90_92), .C1 (n_87_95), .C2 (n_84_93) );
AOI211_X1 g_86_96 (.ZN (n_86_96), .A (n_87_93), .B (n_88_93), .C1 (n_89_94), .C2 (n_83_95) );
AOI211_X1 g_88_95 (.ZN (n_88_95), .A (n_85_94), .B (n_86_92), .C1 (n_90_92), .C2 (n_85_96) );
AOI211_X1 g_89_93 (.ZN (n_89_93), .A (n_86_96), .B (n_88_91), .C1 (n_88_93), .C2 (n_87_95) );
AOI211_X1 g_87_94 (.ZN (n_87_94), .A (n_88_95), .B (n_87_93), .C1 (n_86_92), .C2 (n_89_94) );
AOI211_X1 g_89_95 (.ZN (n_89_95), .A (n_89_93), .B (n_85_94), .C1 (n_88_91), .C2 (n_90_92) );
AOI211_X1 g_91_94 (.ZN (n_91_94), .A (n_87_94), .B (n_86_96), .C1 (n_87_93), .C2 (n_88_93) );
AOI211_X1 g_90_96 (.ZN (n_90_96), .A (n_89_95), .B (n_88_95), .C1 (n_85_94), .C2 (n_86_92) );
AOI211_X1 g_88_97 (.ZN (n_88_97), .A (n_91_94), .B (n_89_93), .C1 (n_86_96), .C2 (n_88_91) );
endmodule
