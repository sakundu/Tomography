VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram45_2048x42
  FOREIGN fakeram45_2048x42 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 193.420 BY 383.600 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.765 0.070 2.835 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.285 0.070 5.355 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.805 0.070 7.875 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.325 0.070 10.395 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.845 0.070 12.915 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.365 0.070 15.435 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.885 0.070 17.955 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.405 0.070 20.475 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.925 0.070 22.995 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.445 0.070 25.515 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.965 0.070 28.035 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.485 0.070 30.555 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.005 0.070 33.075 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.525 0.070 35.595 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.045 0.070 38.115 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.565 0.070 40.635 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.085 0.070 43.155 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.605 0.070 45.675 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.125 0.070 48.195 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.645 0.070 50.715 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.165 0.070 53.235 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.685 0.070 55.755 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 58.205 0.070 58.275 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.725 0.070 60.795 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 63.245 0.070 63.315 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 65.765 0.070 65.835 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.285 0.070 68.355 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.805 0.070 70.875 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.325 0.070 73.395 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.845 0.070 75.915 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.365 0.070 78.435 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.885 0.070 80.955 ;
    END
  END w_mask_in[31]
  PIN w_mask_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.405 0.070 83.475 ;
    END
  END w_mask_in[32]
  PIN w_mask_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.925 0.070 85.995 ;
    END
  END w_mask_in[33]
  PIN w_mask_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 88.445 0.070 88.515 ;
    END
  END w_mask_in[34]
  PIN w_mask_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 90.965 0.070 91.035 ;
    END
  END w_mask_in[35]
  PIN w_mask_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 93.485 0.070 93.555 ;
    END
  END w_mask_in[36]
  PIN w_mask_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 96.005 0.070 96.075 ;
    END
  END w_mask_in[37]
  PIN w_mask_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 98.525 0.070 98.595 ;
    END
  END w_mask_in[38]
  PIN w_mask_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 101.045 0.070 101.115 ;
    END
  END w_mask_in[39]
  PIN w_mask_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 103.565 0.070 103.635 ;
    END
  END w_mask_in[40]
  PIN w_mask_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 106.085 0.070 106.155 ;
    END
  END w_mask_in[41]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 112.245 0.070 112.315 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 114.765 0.070 114.835 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 117.285 0.070 117.355 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 119.805 0.070 119.875 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 122.325 0.070 122.395 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 124.845 0.070 124.915 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 127.365 0.070 127.435 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 129.885 0.070 129.955 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 132.405 0.070 132.475 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 134.925 0.070 134.995 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 137.445 0.070 137.515 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 139.965 0.070 140.035 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 142.485 0.070 142.555 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 145.005 0.070 145.075 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 147.525 0.070 147.595 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 150.045 0.070 150.115 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 152.565 0.070 152.635 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 155.085 0.070 155.155 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 157.605 0.070 157.675 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 160.125 0.070 160.195 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 162.645 0.070 162.715 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 165.165 0.070 165.235 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 167.685 0.070 167.755 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 170.205 0.070 170.275 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 172.725 0.070 172.795 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 175.245 0.070 175.315 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 177.765 0.070 177.835 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 180.285 0.070 180.355 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 182.805 0.070 182.875 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 185.325 0.070 185.395 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 187.845 0.070 187.915 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 190.365 0.070 190.435 ;
    END
  END rd_out[31]
  PIN rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 192.885 0.070 192.955 ;
    END
  END rd_out[32]
  PIN rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 195.405 0.070 195.475 ;
    END
  END rd_out[33]
  PIN rd_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 197.925 0.070 197.995 ;
    END
  END rd_out[34]
  PIN rd_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 200.445 0.070 200.515 ;
    END
  END rd_out[35]
  PIN rd_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 202.965 0.070 203.035 ;
    END
  END rd_out[36]
  PIN rd_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 205.485 0.070 205.555 ;
    END
  END rd_out[37]
  PIN rd_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 208.005 0.070 208.075 ;
    END
  END rd_out[38]
  PIN rd_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 210.525 0.070 210.595 ;
    END
  END rd_out[39]
  PIN rd_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 213.045 0.070 213.115 ;
    END
  END rd_out[40]
  PIN rd_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 215.565 0.070 215.635 ;
    END
  END rd_out[41]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 221.725 0.070 221.795 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 224.245 0.070 224.315 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 226.765 0.070 226.835 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 229.285 0.070 229.355 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 231.805 0.070 231.875 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 234.325 0.070 234.395 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 236.845 0.070 236.915 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 239.365 0.070 239.435 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 241.885 0.070 241.955 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 244.405 0.070 244.475 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 246.925 0.070 246.995 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 249.445 0.070 249.515 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 251.965 0.070 252.035 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 254.485 0.070 254.555 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 257.005 0.070 257.075 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 259.525 0.070 259.595 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 262.045 0.070 262.115 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 264.565 0.070 264.635 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 267.085 0.070 267.155 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 269.605 0.070 269.675 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 272.125 0.070 272.195 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 274.645 0.070 274.715 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 277.165 0.070 277.235 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 279.685 0.070 279.755 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 282.205 0.070 282.275 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 284.725 0.070 284.795 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 287.245 0.070 287.315 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 289.765 0.070 289.835 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 292.285 0.070 292.355 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 294.805 0.070 294.875 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 297.325 0.070 297.395 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 299.845 0.070 299.915 ;
    END
  END wd_in[31]
  PIN wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 302.365 0.070 302.435 ;
    END
  END wd_in[32]
  PIN wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 304.885 0.070 304.955 ;
    END
  END wd_in[33]
  PIN wd_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 307.405 0.070 307.475 ;
    END
  END wd_in[34]
  PIN wd_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 309.925 0.070 309.995 ;
    END
  END wd_in[35]
  PIN wd_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 312.445 0.070 312.515 ;
    END
  END wd_in[36]
  PIN wd_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 314.965 0.070 315.035 ;
    END
  END wd_in[37]
  PIN wd_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 317.485 0.070 317.555 ;
    END
  END wd_in[38]
  PIN wd_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 320.005 0.070 320.075 ;
    END
  END wd_in[39]
  PIN wd_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 322.525 0.070 322.595 ;
    END
  END wd_in[40]
  PIN wd_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 325.045 0.070 325.115 ;
    END
  END wd_in[41]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 331.205 0.070 331.275 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 333.725 0.070 333.795 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 336.245 0.070 336.315 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 338.765 0.070 338.835 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 341.285 0.070 341.355 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 343.805 0.070 343.875 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 346.325 0.070 346.395 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 348.845 0.070 348.915 ;
    END
  END addr_in[7]
  PIN addr_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 351.365 0.070 351.435 ;
    END
  END addr_in[8]
  PIN addr_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 353.885 0.070 353.955 ;
    END
  END addr_in[9]
  PIN addr_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 356.405 0.070 356.475 ;
    END
  END addr_in[10]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 362.565 0.070 362.635 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 365.085 0.070 365.155 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 367.605 0.070 367.675 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 2.660 2.800 2.940 380.800 ;
      RECT 7.140 2.800 7.420 380.800 ;
      RECT 11.620 2.800 11.900 380.800 ;
      RECT 16.100 2.800 16.380 380.800 ;
      RECT 20.580 2.800 20.860 380.800 ;
      RECT 25.060 2.800 25.340 380.800 ;
      RECT 29.540 2.800 29.820 380.800 ;
      RECT 34.020 2.800 34.300 380.800 ;
      RECT 38.500 2.800 38.780 380.800 ;
      RECT 42.980 2.800 43.260 380.800 ;
      RECT 47.460 2.800 47.740 380.800 ;
      RECT 51.940 2.800 52.220 380.800 ;
      RECT 56.420 2.800 56.700 380.800 ;
      RECT 60.900 2.800 61.180 380.800 ;
      RECT 65.380 2.800 65.660 380.800 ;
      RECT 69.860 2.800 70.140 380.800 ;
      RECT 74.340 2.800 74.620 380.800 ;
      RECT 78.820 2.800 79.100 380.800 ;
      RECT 83.300 2.800 83.580 380.800 ;
      RECT 87.780 2.800 88.060 380.800 ;
      RECT 92.260 2.800 92.540 380.800 ;
      RECT 96.740 2.800 97.020 380.800 ;
      RECT 101.220 2.800 101.500 380.800 ;
      RECT 105.700 2.800 105.980 380.800 ;
      RECT 110.180 2.800 110.460 380.800 ;
      RECT 114.660 2.800 114.940 380.800 ;
      RECT 119.140 2.800 119.420 380.800 ;
      RECT 123.620 2.800 123.900 380.800 ;
      RECT 128.100 2.800 128.380 380.800 ;
      RECT 132.580 2.800 132.860 380.800 ;
      RECT 137.060 2.800 137.340 380.800 ;
      RECT 141.540 2.800 141.820 380.800 ;
      RECT 146.020 2.800 146.300 380.800 ;
      RECT 150.500 2.800 150.780 380.800 ;
      RECT 154.980 2.800 155.260 380.800 ;
      RECT 159.460 2.800 159.740 380.800 ;
      RECT 163.940 2.800 164.220 380.800 ;
      RECT 168.420 2.800 168.700 380.800 ;
      RECT 172.900 2.800 173.180 380.800 ;
      RECT 177.380 2.800 177.660 380.800 ;
      RECT 181.860 2.800 182.140 380.800 ;
      RECT 186.340 2.800 186.620 380.800 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 4.900 2.800 5.180 380.800 ;
      RECT 9.380 2.800 9.660 380.800 ;
      RECT 13.860 2.800 14.140 380.800 ;
      RECT 18.340 2.800 18.620 380.800 ;
      RECT 22.820 2.800 23.100 380.800 ;
      RECT 27.300 2.800 27.580 380.800 ;
      RECT 31.780 2.800 32.060 380.800 ;
      RECT 36.260 2.800 36.540 380.800 ;
      RECT 40.740 2.800 41.020 380.800 ;
      RECT 45.220 2.800 45.500 380.800 ;
      RECT 49.700 2.800 49.980 380.800 ;
      RECT 54.180 2.800 54.460 380.800 ;
      RECT 58.660 2.800 58.940 380.800 ;
      RECT 63.140 2.800 63.420 380.800 ;
      RECT 67.620 2.800 67.900 380.800 ;
      RECT 72.100 2.800 72.380 380.800 ;
      RECT 76.580 2.800 76.860 380.800 ;
      RECT 81.060 2.800 81.340 380.800 ;
      RECT 85.540 2.800 85.820 380.800 ;
      RECT 90.020 2.800 90.300 380.800 ;
      RECT 94.500 2.800 94.780 380.800 ;
      RECT 98.980 2.800 99.260 380.800 ;
      RECT 103.460 2.800 103.740 380.800 ;
      RECT 107.940 2.800 108.220 380.800 ;
      RECT 112.420 2.800 112.700 380.800 ;
      RECT 116.900 2.800 117.180 380.800 ;
      RECT 121.380 2.800 121.660 380.800 ;
      RECT 125.860 2.800 126.140 380.800 ;
      RECT 130.340 2.800 130.620 380.800 ;
      RECT 134.820 2.800 135.100 380.800 ;
      RECT 139.300 2.800 139.580 380.800 ;
      RECT 143.780 2.800 144.060 380.800 ;
      RECT 148.260 2.800 148.540 380.800 ;
      RECT 152.740 2.800 153.020 380.800 ;
      RECT 157.220 2.800 157.500 380.800 ;
      RECT 161.700 2.800 161.980 380.800 ;
      RECT 166.180 2.800 166.460 380.800 ;
      RECT 170.660 2.800 170.940 380.800 ;
      RECT 175.140 2.800 175.420 380.800 ;
      RECT 179.620 2.800 179.900 380.800 ;
      RECT 184.100 2.800 184.380 380.800 ;
      RECT 188.580 2.800 188.860 380.800 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 193.420 383.600 ;
    LAYER metal2 ;
    RECT 0 0 193.420 383.600 ;
    LAYER metal3 ;
    RECT 0.070 0 193.420 383.600 ;
    RECT 0 0.000 0.070 2.765 ;
    RECT 0 2.835 0.070 5.285 ;
    RECT 0 5.355 0.070 7.805 ;
    RECT 0 7.875 0.070 10.325 ;
    RECT 0 10.395 0.070 12.845 ;
    RECT 0 12.915 0.070 15.365 ;
    RECT 0 15.435 0.070 17.885 ;
    RECT 0 17.955 0.070 20.405 ;
    RECT 0 20.475 0.070 22.925 ;
    RECT 0 22.995 0.070 25.445 ;
    RECT 0 25.515 0.070 27.965 ;
    RECT 0 28.035 0.070 30.485 ;
    RECT 0 30.555 0.070 33.005 ;
    RECT 0 33.075 0.070 35.525 ;
    RECT 0 35.595 0.070 38.045 ;
    RECT 0 38.115 0.070 40.565 ;
    RECT 0 40.635 0.070 43.085 ;
    RECT 0 43.155 0.070 45.605 ;
    RECT 0 45.675 0.070 48.125 ;
    RECT 0 48.195 0.070 50.645 ;
    RECT 0 50.715 0.070 53.165 ;
    RECT 0 53.235 0.070 55.685 ;
    RECT 0 55.755 0.070 58.205 ;
    RECT 0 58.275 0.070 60.725 ;
    RECT 0 60.795 0.070 63.245 ;
    RECT 0 63.315 0.070 65.765 ;
    RECT 0 65.835 0.070 68.285 ;
    RECT 0 68.355 0.070 70.805 ;
    RECT 0 70.875 0.070 73.325 ;
    RECT 0 73.395 0.070 75.845 ;
    RECT 0 75.915 0.070 78.365 ;
    RECT 0 78.435 0.070 80.885 ;
    RECT 0 80.955 0.070 83.405 ;
    RECT 0 83.475 0.070 85.925 ;
    RECT 0 85.995 0.070 88.445 ;
    RECT 0 88.515 0.070 90.965 ;
    RECT 0 91.035 0.070 93.485 ;
    RECT 0 93.555 0.070 96.005 ;
    RECT 0 96.075 0.070 98.525 ;
    RECT 0 98.595 0.070 101.045 ;
    RECT 0 101.115 0.070 103.565 ;
    RECT 0 103.635 0.070 106.085 ;
    RECT 0 106.155 0.070 112.245 ;
    RECT 0 112.315 0.070 114.765 ;
    RECT 0 114.835 0.070 117.285 ;
    RECT 0 117.355 0.070 119.805 ;
    RECT 0 119.875 0.070 122.325 ;
    RECT 0 122.395 0.070 124.845 ;
    RECT 0 124.915 0.070 127.365 ;
    RECT 0 127.435 0.070 129.885 ;
    RECT 0 129.955 0.070 132.405 ;
    RECT 0 132.475 0.070 134.925 ;
    RECT 0 134.995 0.070 137.445 ;
    RECT 0 137.515 0.070 139.965 ;
    RECT 0 140.035 0.070 142.485 ;
    RECT 0 142.555 0.070 145.005 ;
    RECT 0 145.075 0.070 147.525 ;
    RECT 0 147.595 0.070 150.045 ;
    RECT 0 150.115 0.070 152.565 ;
    RECT 0 152.635 0.070 155.085 ;
    RECT 0 155.155 0.070 157.605 ;
    RECT 0 157.675 0.070 160.125 ;
    RECT 0 160.195 0.070 162.645 ;
    RECT 0 162.715 0.070 165.165 ;
    RECT 0 165.235 0.070 167.685 ;
    RECT 0 167.755 0.070 170.205 ;
    RECT 0 170.275 0.070 172.725 ;
    RECT 0 172.795 0.070 175.245 ;
    RECT 0 175.315 0.070 177.765 ;
    RECT 0 177.835 0.070 180.285 ;
    RECT 0 180.355 0.070 182.805 ;
    RECT 0 182.875 0.070 185.325 ;
    RECT 0 185.395 0.070 187.845 ;
    RECT 0 187.915 0.070 190.365 ;
    RECT 0 190.435 0.070 192.885 ;
    RECT 0 192.955 0.070 195.405 ;
    RECT 0 195.475 0.070 197.925 ;
    RECT 0 197.995 0.070 200.445 ;
    RECT 0 200.515 0.070 202.965 ;
    RECT 0 203.035 0.070 205.485 ;
    RECT 0 205.555 0.070 208.005 ;
    RECT 0 208.075 0.070 210.525 ;
    RECT 0 210.595 0.070 213.045 ;
    RECT 0 213.115 0.070 215.565 ;
    RECT 0 215.635 0.070 221.725 ;
    RECT 0 221.795 0.070 224.245 ;
    RECT 0 224.315 0.070 226.765 ;
    RECT 0 226.835 0.070 229.285 ;
    RECT 0 229.355 0.070 231.805 ;
    RECT 0 231.875 0.070 234.325 ;
    RECT 0 234.395 0.070 236.845 ;
    RECT 0 236.915 0.070 239.365 ;
    RECT 0 239.435 0.070 241.885 ;
    RECT 0 241.955 0.070 244.405 ;
    RECT 0 244.475 0.070 246.925 ;
    RECT 0 246.995 0.070 249.445 ;
    RECT 0 249.515 0.070 251.965 ;
    RECT 0 252.035 0.070 254.485 ;
    RECT 0 254.555 0.070 257.005 ;
    RECT 0 257.075 0.070 259.525 ;
    RECT 0 259.595 0.070 262.045 ;
    RECT 0 262.115 0.070 264.565 ;
    RECT 0 264.635 0.070 267.085 ;
    RECT 0 267.155 0.070 269.605 ;
    RECT 0 269.675 0.070 272.125 ;
    RECT 0 272.195 0.070 274.645 ;
    RECT 0 274.715 0.070 277.165 ;
    RECT 0 277.235 0.070 279.685 ;
    RECT 0 279.755 0.070 282.205 ;
    RECT 0 282.275 0.070 284.725 ;
    RECT 0 284.795 0.070 287.245 ;
    RECT 0 287.315 0.070 289.765 ;
    RECT 0 289.835 0.070 292.285 ;
    RECT 0 292.355 0.070 294.805 ;
    RECT 0 294.875 0.070 297.325 ;
    RECT 0 297.395 0.070 299.845 ;
    RECT 0 299.915 0.070 302.365 ;
    RECT 0 302.435 0.070 304.885 ;
    RECT 0 304.955 0.070 307.405 ;
    RECT 0 307.475 0.070 309.925 ;
    RECT 0 309.995 0.070 312.445 ;
    RECT 0 312.515 0.070 314.965 ;
    RECT 0 315.035 0.070 317.485 ;
    RECT 0 317.555 0.070 320.005 ;
    RECT 0 320.075 0.070 322.525 ;
    RECT 0 322.595 0.070 325.045 ;
    RECT 0 325.115 0.070 331.205 ;
    RECT 0 331.275 0.070 333.725 ;
    RECT 0 333.795 0.070 336.245 ;
    RECT 0 336.315 0.070 338.765 ;
    RECT 0 338.835 0.070 341.285 ;
    RECT 0 341.355 0.070 343.805 ;
    RECT 0 343.875 0.070 346.325 ;
    RECT 0 346.395 0.070 348.845 ;
    RECT 0 348.915 0.070 351.365 ;
    RECT 0 351.435 0.070 353.885 ;
    RECT 0 353.955 0.070 356.405 ;
    RECT 0 356.475 0.070 362.565 ;
    RECT 0 362.635 0.070 365.085 ;
    RECT 0 365.155 0.070 367.605 ;
    RECT 0 367.675 0.070 383.600 ;
    LAYER metal4 ;
    RECT 0 0 193.420 2.800 ;
    RECT 0 380.800 193.420 383.600 ;
    RECT 0.000 2.800 2.660 380.800 ;
    RECT 2.940 2.800 4.900 380.800 ;
    RECT 5.180 2.800 7.140 380.800 ;
    RECT 7.420 2.800 9.380 380.800 ;
    RECT 9.660 2.800 11.620 380.800 ;
    RECT 11.900 2.800 13.860 380.800 ;
    RECT 14.140 2.800 16.100 380.800 ;
    RECT 16.380 2.800 18.340 380.800 ;
    RECT 18.620 2.800 20.580 380.800 ;
    RECT 20.860 2.800 22.820 380.800 ;
    RECT 23.100 2.800 25.060 380.800 ;
    RECT 25.340 2.800 27.300 380.800 ;
    RECT 27.580 2.800 29.540 380.800 ;
    RECT 29.820 2.800 31.780 380.800 ;
    RECT 32.060 2.800 34.020 380.800 ;
    RECT 34.300 2.800 36.260 380.800 ;
    RECT 36.540 2.800 38.500 380.800 ;
    RECT 38.780 2.800 40.740 380.800 ;
    RECT 41.020 2.800 42.980 380.800 ;
    RECT 43.260 2.800 45.220 380.800 ;
    RECT 45.500 2.800 47.460 380.800 ;
    RECT 47.740 2.800 49.700 380.800 ;
    RECT 49.980 2.800 51.940 380.800 ;
    RECT 52.220 2.800 54.180 380.800 ;
    RECT 54.460 2.800 56.420 380.800 ;
    RECT 56.700 2.800 58.660 380.800 ;
    RECT 58.940 2.800 60.900 380.800 ;
    RECT 61.180 2.800 63.140 380.800 ;
    RECT 63.420 2.800 65.380 380.800 ;
    RECT 65.660 2.800 67.620 380.800 ;
    RECT 67.900 2.800 69.860 380.800 ;
    RECT 70.140 2.800 72.100 380.800 ;
    RECT 72.380 2.800 74.340 380.800 ;
    RECT 74.620 2.800 76.580 380.800 ;
    RECT 76.860 2.800 78.820 380.800 ;
    RECT 79.100 2.800 81.060 380.800 ;
    RECT 81.340 2.800 83.300 380.800 ;
    RECT 83.580 2.800 85.540 380.800 ;
    RECT 85.820 2.800 87.780 380.800 ;
    RECT 88.060 2.800 90.020 380.800 ;
    RECT 90.300 2.800 92.260 380.800 ;
    RECT 92.540 2.800 94.500 380.800 ;
    RECT 94.780 2.800 96.740 380.800 ;
    RECT 97.020 2.800 98.980 380.800 ;
    RECT 99.260 2.800 101.220 380.800 ;
    RECT 101.500 2.800 103.460 380.800 ;
    RECT 103.740 2.800 105.700 380.800 ;
    RECT 105.980 2.800 107.940 380.800 ;
    RECT 108.220 2.800 110.180 380.800 ;
    RECT 110.460 2.800 112.420 380.800 ;
    RECT 112.700 2.800 114.660 380.800 ;
    RECT 114.940 2.800 116.900 380.800 ;
    RECT 117.180 2.800 119.140 380.800 ;
    RECT 119.420 2.800 121.380 380.800 ;
    RECT 121.660 2.800 123.620 380.800 ;
    RECT 123.900 2.800 125.860 380.800 ;
    RECT 126.140 2.800 128.100 380.800 ;
    RECT 128.380 2.800 130.340 380.800 ;
    RECT 130.620 2.800 132.580 380.800 ;
    RECT 132.860 2.800 134.820 380.800 ;
    RECT 135.100 2.800 137.060 380.800 ;
    RECT 137.340 2.800 139.300 380.800 ;
    RECT 139.580 2.800 141.540 380.800 ;
    RECT 141.820 2.800 143.780 380.800 ;
    RECT 144.060 2.800 146.020 380.800 ;
    RECT 146.300 2.800 148.260 380.800 ;
    RECT 148.540 2.800 150.500 380.800 ;
    RECT 150.780 2.800 152.740 380.800 ;
    RECT 153.020 2.800 154.980 380.800 ;
    RECT 155.260 2.800 157.220 380.800 ;
    RECT 157.500 2.800 159.460 380.800 ;
    RECT 159.740 2.800 161.700 380.800 ;
    RECT 161.980 2.800 163.940 380.800 ;
    RECT 164.220 2.800 166.180 380.800 ;
    RECT 166.460 2.800 168.420 380.800 ;
    RECT 168.700 2.800 170.660 380.800 ;
    RECT 170.940 2.800 172.900 380.800 ;
    RECT 173.180 2.800 175.140 380.800 ;
    RECT 175.420 2.800 177.380 380.800 ;
    RECT 177.660 2.800 179.620 380.800 ;
    RECT 179.900 2.800 181.860 380.800 ;
    RECT 182.140 2.800 184.100 380.800 ;
    RECT 184.380 2.800 186.340 380.800 ;
    RECT 186.620 2.800 188.580 380.800 ;
    RECT 188.860 2.800 193.420 380.800 ;
    LAYER OVERLAP ;
    RECT 0 0 193.420 383.600 ;
  END
END fakeram45_2048x42

END LIBRARY
